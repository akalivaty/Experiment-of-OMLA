

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n684), .A2(n798), .ZN(n725) );
  NAND2_X1 U552 ( .A1(G8), .A2(n725), .ZN(n767) );
  AND2_X1 U553 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U554 ( .A1(G651), .A2(n644), .ZN(n656) );
  NOR2_X1 U555 ( .A1(n743), .A2(n687), .ZN(n688) );
  NOR2_X1 U556 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U557 ( .A1(n725), .A2(G2084), .ZN(n686) );
  AND2_X1 U558 ( .A1(n761), .A2(n752), .ZN(n753) );
  AND2_X1 U559 ( .A1(n813), .A2(n823), .ZN(n814) );
  INV_X1 U560 ( .A(KEYINPUT17), .ZN(n524) );
  AND2_X1 U561 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U562 ( .A1(n997), .A2(G138), .ZN(n534) );
  XOR2_X1 U563 ( .A(G2104), .B(KEYINPUT64), .Z(n519) );
  NOR2_X1 U564 ( .A1(n519), .A2(G2105), .ZN(n620) );
  NAND2_X1 U565 ( .A1(G101), .A2(n620), .ZN(n518) );
  XOR2_X1 U566 ( .A(n518), .B(KEYINPUT23), .Z(n523) );
  AND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n993) );
  NAND2_X1 U568 ( .A1(G113), .A2(n993), .ZN(n521) );
  AND2_X2 U569 ( .A1(G2105), .A2(n519), .ZN(n994) );
  NAND2_X1 U570 ( .A1(G125), .A2(n994), .ZN(n520) );
  AND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XNOR2_X2 U574 ( .A(n525), .B(n524), .ZN(n997) );
  AND2_X1 U575 ( .A1(n997), .A2(G137), .ZN(n527) );
  INV_X1 U576 ( .A(KEYINPUT65), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n527), .B(n526), .ZN(n528) );
  NOR2_X2 U578 ( .A1(n529), .A2(n528), .ZN(G160) );
  AND2_X1 U579 ( .A1(G114), .A2(n993), .ZN(n533) );
  NAND2_X1 U580 ( .A1(G102), .A2(n620), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G126), .A2(n994), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n534), .B(KEYINPUT80), .ZN(n535) );
  AND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(G164) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U587 ( .A1(G85), .A2(n649), .ZN(n538) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  INV_X1 U589 ( .A(G651), .ZN(n539) );
  NOR2_X1 U590 ( .A1(n644), .A2(n539), .ZN(n652) );
  NAND2_X1 U591 ( .A1(G72), .A2(n652), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U593 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n540), .Z(n648) );
  NAND2_X1 U595 ( .A1(G60), .A2(n648), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G47), .A2(n656), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G290) );
  XNOR2_X1 U599 ( .A(G1348), .B(G2427), .ZN(n554) );
  XOR2_X1 U600 ( .A(G2451), .B(KEYINPUT103), .Z(n546) );
  XNOR2_X1 U601 ( .A(G1341), .B(G2443), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n546), .B(n545), .ZN(n550) );
  XOR2_X1 U603 ( .A(G2438), .B(G2435), .Z(n548) );
  XNOR2_X1 U604 ( .A(G2430), .B(G2454), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U606 ( .A(n550), .B(n549), .Z(n552) );
  XNOR2_X1 U607 ( .A(G2446), .B(KEYINPUT104), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n554), .B(n553), .ZN(n555) );
  AND2_X1 U610 ( .A1(n555), .A2(G14), .ZN(G401) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(G88), .A2(n649), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G75), .A2(n652), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G62), .A2(n648), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G50), .A2(n656), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U620 ( .A1(n561), .A2(n560), .ZN(G166) );
  NAND2_X1 U621 ( .A1(G63), .A2(n648), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G51), .A2(n656), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT6), .B(n564), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n649), .A2(G89), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G76), .A2(n652), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U629 ( .A(n568), .B(KEYINPUT5), .Z(n569) );
  NOR2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT7), .B(n571), .Z(n572) );
  XNOR2_X1 U632 ( .A(KEYINPUT70), .B(n572), .ZN(G168) );
  XOR2_X1 U633 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U634 ( .A1(G94), .A2(G452), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n573), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n834) );
  NAND2_X1 U639 ( .A1(n834), .A2(G567), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n648), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n576), .Z(n582) );
  NAND2_X1 U643 ( .A1(n649), .A2(G81), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G68), .A2(n652), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n656), .A2(G43), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n967) );
  INV_X1 U651 ( .A(G860), .ZN(n612) );
  OR2_X1 U652 ( .A1(n967), .A2(n612), .ZN(G153) );
  NAND2_X1 U653 ( .A1(n649), .A2(G90), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n585), .B(KEYINPUT66), .ZN(n587) );
  NAND2_X1 U655 ( .A1(G77), .A2(n652), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U657 ( .A(KEYINPUT9), .B(n588), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G64), .A2(n648), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G52), .A2(n656), .ZN(n589) );
  AND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G301) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n656), .A2(G54), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G66), .A2(n648), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G79), .A2(n652), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G92), .A2(n649), .ZN(n595) );
  XNOR2_X1 U668 ( .A(KEYINPUT69), .B(n595), .ZN(n596) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X2 U671 ( .A(KEYINPUT15), .B(n600), .Z(n970) );
  INV_X1 U672 ( .A(G868), .ZN(n666) );
  NAND2_X1 U673 ( .A1(n970), .A2(n666), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G65), .A2(n648), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G53), .A2(n656), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G91), .A2(n649), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G78), .A2(n652), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n948) );
  XOR2_X1 U682 ( .A(n948), .B(KEYINPUT68), .Z(G299) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(G868), .ZN(n609) );
  NOR2_X1 U684 ( .A1(G286), .A2(n609), .ZN(n611) );
  NOR2_X1 U685 ( .A1(G299), .A2(G868), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n612), .A2(G559), .ZN(n613) );
  INV_X1 U688 ( .A(n970), .ZN(n701) );
  NAND2_X1 U689 ( .A1(n613), .A2(n701), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT72), .ZN(n615) );
  XNOR2_X1 U691 ( .A(KEYINPUT16), .B(n615), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G559), .A2(n666), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n701), .A2(n616), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT73), .ZN(n619) );
  NOR2_X1 U695 ( .A1(n967), .A2(G868), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(G282) );
  BUF_X1 U697 ( .A(n620), .Z(n998) );
  NAND2_X1 U698 ( .A1(G99), .A2(n998), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G111), .A2(n993), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT74), .B(n623), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G123), .A2(n994), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT18), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n997), .A2(G135), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n1018) );
  XNOR2_X1 U707 ( .A(n1018), .B(G2096), .ZN(n630) );
  INV_X1 U708 ( .A(G2100), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G559), .A2(n701), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n967), .B(n631), .ZN(n664) );
  NOR2_X1 U712 ( .A1(n664), .A2(G860), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G93), .A2(n649), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G80), .A2(n652), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G67), .A2(n648), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G55), .A2(n656), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U719 ( .A(KEYINPUT75), .B(n636), .Z(n637) );
  NOR2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n667) );
  XNOR2_X1 U721 ( .A(n639), .B(n667), .ZN(G145) );
  NAND2_X1 U722 ( .A1(n656), .A2(G49), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(KEYINPUT76), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U726 ( .A1(n648), .A2(n643), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G87), .A2(n644), .ZN(n645) );
  XOR2_X1 U728 ( .A(KEYINPUT77), .B(n645), .Z(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U730 ( .A1(G61), .A2(n648), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G86), .A2(n649), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n652), .A2(G73), .ZN(n653) );
  XOR2_X1 U734 ( .A(KEYINPUT2), .B(n653), .Z(n654) );
  NOR2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n656), .A2(G48), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(G305) );
  XNOR2_X1 U738 ( .A(KEYINPUT19), .B(G299), .ZN(n660) );
  XNOR2_X1 U739 ( .A(G305), .B(G166), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U741 ( .A(n661), .B(G290), .Z(n662) );
  XNOR2_X1 U742 ( .A(G288), .B(n662), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n667), .B(n663), .ZN(n968) );
  XOR2_X1 U744 ( .A(n664), .B(n968), .Z(n665) );
  NAND2_X1 U745 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U748 ( .A(KEYINPUT78), .B(n670), .Z(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U757 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G96), .A2(n677), .ZN(n965) );
  NAND2_X1 U759 ( .A1(n965), .A2(G2106), .ZN(n681) );
  NAND2_X1 U760 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U761 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U762 ( .A1(G108), .A2(n679), .ZN(n966) );
  NAND2_X1 U763 ( .A1(n966), .A2(G567), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n1028) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n682) );
  NOR2_X1 U766 ( .A1(n1028), .A2(n682), .ZN(n683) );
  XOR2_X1 U767 ( .A(KEYINPUT79), .B(n683), .Z(n838) );
  NAND2_X1 U768 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G301), .ZN(G171) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n797) );
  INV_X1 U772 ( .A(n797), .ZN(n684) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n798) );
  NOR2_X1 U774 ( .A1(n767), .A2(G1966), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT88), .ZN(n743) );
  XNOR2_X1 U776 ( .A(n686), .B(KEYINPUT87), .ZN(n739) );
  NAND2_X1 U777 ( .A1(G8), .A2(n739), .ZN(n687) );
  XOR2_X1 U778 ( .A(KEYINPUT30), .B(n688), .Z(n689) );
  NOR2_X1 U779 ( .A1(G168), .A2(n689), .ZN(n693) );
  XNOR2_X1 U780 ( .A(G1961), .B(KEYINPUT89), .ZN(n871) );
  NAND2_X1 U781 ( .A1(n725), .A2(n871), .ZN(n691) );
  INV_X1 U782 ( .A(n725), .ZN(n706) );
  XNOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .ZN(n854) );
  NAND2_X1 U784 ( .A1(n706), .A2(n854), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n696) );
  NOR2_X1 U786 ( .A1(G171), .A2(n696), .ZN(n692) );
  XOR2_X1 U787 ( .A(n694), .B(KEYINPUT31), .Z(n695) );
  XNOR2_X1 U788 ( .A(n695), .B(KEYINPUT94), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n696), .A2(G171), .ZN(n724) );
  NAND2_X1 U790 ( .A1(n706), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U791 ( .A(n697), .B(KEYINPUT27), .ZN(n699) );
  XOR2_X1 U792 ( .A(G1956), .B(KEYINPUT90), .Z(n883) );
  NOR2_X1 U793 ( .A1(n706), .A2(n883), .ZN(n698) );
  NOR2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n716) );
  NOR2_X1 U795 ( .A1(n716), .A2(n948), .ZN(n700) );
  XOR2_X1 U796 ( .A(KEYINPUT28), .B(n700), .Z(n721) );
  NAND2_X1 U797 ( .A1(G1341), .A2(n725), .ZN(n711) );
  AND2_X1 U798 ( .A1(n701), .A2(n711), .ZN(n704) );
  XNOR2_X1 U799 ( .A(G1996), .B(KEYINPUT91), .ZN(n853) );
  NOR2_X1 U800 ( .A1(n725), .A2(n853), .ZN(n702) );
  XNOR2_X1 U801 ( .A(n702), .B(KEYINPUT26), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n703), .A2(n967), .ZN(n712) );
  AND2_X1 U803 ( .A1(n704), .A2(n712), .ZN(n705) );
  XOR2_X1 U804 ( .A(n705), .B(KEYINPUT92), .Z(n710) );
  NOR2_X1 U805 ( .A1(n706), .A2(G1348), .ZN(n708) );
  NOR2_X1 U806 ( .A1(G2067), .A2(n725), .ZN(n707) );
  NOR2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U810 ( .A1(n970), .A2(n713), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n948), .A2(n716), .ZN(n717) );
  XOR2_X1 U813 ( .A(KEYINPUT93), .B(n717), .Z(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U816 ( .A(KEYINPUT29), .B(n722), .Z(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n741) );
  INV_X1 U818 ( .A(G8), .ZN(n730) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n767), .ZN(n727) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n728), .A2(G303), .ZN(n729) );
  OR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n732) );
  AND2_X1 U824 ( .A1(n741), .A2(n732), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n742), .A2(n731), .ZN(n736) );
  INV_X1 U826 ( .A(n732), .ZN(n734) );
  AND2_X1 U827 ( .A1(G286), .A2(G8), .ZN(n733) );
  OR2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n738) );
  XOR2_X1 U830 ( .A(KEYINPUT32), .B(KEYINPUT95), .Z(n737) );
  XNOR2_X1 U831 ( .A(n738), .B(n737), .ZN(n748) );
  INV_X1 U832 ( .A(n739), .ZN(n740) );
  NAND2_X1 U833 ( .A1(G8), .A2(n740), .ZN(n746) );
  AND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n761) );
  NOR2_X1 U838 ( .A1(G288), .A2(G1976), .ZN(n749) );
  XOR2_X1 U839 ( .A(n749), .B(KEYINPUT96), .Z(n951) );
  INV_X1 U840 ( .A(n951), .ZN(n751) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n767), .A2(n753), .ZN(n754) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NAND2_X1 U845 ( .A1(n754), .A2(n952), .ZN(n765) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n755) );
  XOR2_X1 U848 ( .A(n755), .B(KEYINPUT24), .Z(n756) );
  NOR2_X1 U849 ( .A1(n767), .A2(n756), .ZN(n757) );
  XNOR2_X1 U850 ( .A(n757), .B(KEYINPUT86), .ZN(n774) );
  INV_X1 U851 ( .A(n774), .ZN(n758) );
  AND2_X1 U852 ( .A1(n769), .A2(n758), .ZN(n763) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U854 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n767), .A2(n762), .ZN(n766) );
  AND2_X1 U857 ( .A1(n763), .A2(n766), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n778) );
  INV_X1 U859 ( .A(n766), .ZN(n776) );
  XNOR2_X1 U860 ( .A(G1981), .B(G305), .ZN(n941) );
  INV_X1 U861 ( .A(n941), .ZN(n772) );
  OR2_X1 U862 ( .A1(n767), .A2(n951), .ZN(n768) );
  NOR2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U864 ( .A(n770), .B(KEYINPUT97), .ZN(n771) );
  AND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  OR2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n779), .B(KEYINPUT98), .ZN(n815) );
  NAND2_X1 U869 ( .A1(G141), .A2(n997), .ZN(n780) );
  XNOR2_X1 U870 ( .A(n780), .B(KEYINPUT84), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G117), .A2(n993), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G129), .A2(n994), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n998), .A2(G105), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n1009) );
  NAND2_X1 U878 ( .A1(G1996), .A2(n1009), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G131), .A2(n997), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G95), .A2(n998), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U882 ( .A(KEYINPUT83), .B(n790), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G107), .A2(n993), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G119), .A2(n994), .ZN(n791) );
  AND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n1004) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n1004), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n908) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U890 ( .A(KEYINPUT81), .B(n799), .Z(n827) );
  NAND2_X1 U891 ( .A1(n908), .A2(n827), .ZN(n800) );
  XNOR2_X1 U892 ( .A(n800), .B(KEYINPUT85), .ZN(n820) );
  XOR2_X1 U893 ( .A(G1986), .B(G290), .Z(n939) );
  INV_X1 U894 ( .A(n827), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n939), .A2(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n820), .A2(n802), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G140), .A2(n997), .ZN(n804) );
  NAND2_X1 U898 ( .A1(G104), .A2(n998), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U900 ( .A(KEYINPUT34), .B(n805), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G116), .A2(n993), .ZN(n807) );
  NAND2_X1 U902 ( .A1(G128), .A2(n994), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U904 ( .A(KEYINPUT82), .B(n808), .Z(n809) );
  XNOR2_X1 U905 ( .A(KEYINPUT35), .B(n809), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U907 ( .A(KEYINPUT36), .B(n812), .ZN(n1014) );
  XNOR2_X1 U908 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NOR2_X1 U909 ( .A1(n1014), .A2(n825), .ZN(n909) );
  NAND2_X1 U910 ( .A1(n827), .A2(n909), .ZN(n823) );
  XNOR2_X1 U911 ( .A(n816), .B(KEYINPUT99), .ZN(n830) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n1009), .ZN(n906) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n1004), .ZN(n902) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n902), .A2(n817), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n818), .B(KEYINPUT100), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n906), .A2(n821), .ZN(n822) );
  XNOR2_X1 U919 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n1014), .A2(n825), .ZN(n903) );
  NAND2_X1 U922 ( .A1(n826), .A2(n903), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n833) );
  XOR2_X1 U925 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n831), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n836) );
  INV_X1 U930 ( .A(G661), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n837), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G1), .A2(G3), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U935 ( .A(n840), .B(KEYINPUT106), .ZN(G188) );
  NAND2_X1 U937 ( .A1(G124), .A2(n994), .ZN(n841) );
  XOR2_X1 U938 ( .A(KEYINPUT109), .B(n841), .Z(n842) );
  XNOR2_X1 U939 ( .A(n842), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U940 ( .A1(G136), .A2(n997), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U942 ( .A(KEYINPUT110), .B(n845), .ZN(n849) );
  NAND2_X1 U943 ( .A1(G100), .A2(n998), .ZN(n847) );
  NAND2_X1 U944 ( .A1(G112), .A2(n993), .ZN(n846) );
  NAND2_X1 U945 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U946 ( .A1(n849), .A2(n848), .ZN(G162) );
  INV_X1 U947 ( .A(KEYINPUT55), .ZN(n931) );
  XNOR2_X1 U948 ( .A(G2090), .B(G35), .ZN(n863) );
  XOR2_X1 U949 ( .A(G1991), .B(G25), .Z(n850) );
  NAND2_X1 U950 ( .A1(n850), .A2(G28), .ZN(n860) );
  XNOR2_X1 U951 ( .A(G2067), .B(G26), .ZN(n852) );
  XNOR2_X1 U952 ( .A(G33), .B(G2072), .ZN(n851) );
  NOR2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n858) );
  XOR2_X1 U954 ( .A(n853), .B(G32), .Z(n856) );
  XOR2_X1 U955 ( .A(n854), .B(G27), .Z(n855) );
  NOR2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U959 ( .A(KEYINPUT53), .B(n861), .ZN(n862) );
  NOR2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n866) );
  XOR2_X1 U961 ( .A(G2084), .B(G34), .Z(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT54), .B(n864), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n931), .B(n867), .ZN(n869) );
  INV_X1 U965 ( .A(G29), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G11), .A2(n870), .ZN(n901) );
  XOR2_X1 U968 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n897) );
  XNOR2_X1 U969 ( .A(KEYINPUT121), .B(G5), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n879) );
  XNOR2_X1 U971 ( .A(G1976), .B(G23), .ZN(n874) );
  XNOR2_X1 U972 ( .A(G1971), .B(G22), .ZN(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n876) );
  XOR2_X1 U974 ( .A(G1986), .B(G24), .Z(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U976 ( .A(KEYINPUT58), .B(n877), .ZN(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n895) );
  XNOR2_X1 U978 ( .A(G1966), .B(G21), .ZN(n893) );
  XNOR2_X1 U979 ( .A(G1981), .B(G6), .ZN(n881) );
  XNOR2_X1 U980 ( .A(G19), .B(G1341), .ZN(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT122), .B(n882), .Z(n885) );
  XOR2_X1 U983 ( .A(n883), .B(G20), .Z(n884) );
  NOR2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n889) );
  XOR2_X1 U985 ( .A(G4), .B(KEYINPUT123), .Z(n887) );
  XNOR2_X1 U986 ( .A(G1348), .B(KEYINPUT59), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n890), .B(KEYINPUT60), .ZN(n891) );
  XNOR2_X1 U990 ( .A(KEYINPUT124), .B(n891), .ZN(n892) );
  NOR2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U994 ( .A1(n898), .A2(G16), .ZN(n899) );
  XNOR2_X1 U995 ( .A(KEYINPUT126), .B(n899), .ZN(n900) );
  NOR2_X1 U996 ( .A1(n901), .A2(n900), .ZN(n935) );
  NOR2_X1 U997 ( .A1(n902), .A2(n1018), .ZN(n904) );
  NAND2_X1 U998 ( .A1(n904), .A2(n903), .ZN(n929) );
  XOR2_X1 U999 ( .A(G2090), .B(G162), .Z(n905) );
  NOR2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1001 ( .A(KEYINPUT51), .B(n907), .Z(n927) );
  XNOR2_X1 U1002 ( .A(G160), .B(G2084), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n925) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n997), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n998), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(n920) );
  NAND2_X1 U1008 ( .A1(n993), .A2(G115), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n914), .B(KEYINPUT112), .ZN(n916) );
  NAND2_X1 U1010 ( .A1(G127), .A2(n994), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT47), .B(n917), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT113), .B(n918), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n1017) );
  XOR2_X1 U1015 ( .A(G2072), .B(n1017), .Z(n922) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n921) );
  NOR2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1018 ( .A(KEYINPUT50), .B(n923), .Z(n924) );
  NOR2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(KEYINPUT52), .B(n930), .ZN(n932) );
  NAND2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1024 ( .A1(n933), .A2(G29), .ZN(n934) );
  NAND2_X1 U1025 ( .A1(n935), .A2(n934), .ZN(n963) );
  XNOR2_X1 U1026 ( .A(G301), .B(G1961), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(n967), .B(G1341), .ZN(n936) );
  NOR2_X1 U1028 ( .A1(n937), .A2(n936), .ZN(n947) );
  XOR2_X1 U1029 ( .A(G1348), .B(n970), .Z(n938) );
  NAND2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1031 ( .A(G1966), .B(G168), .Z(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT57), .B(n942), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(KEYINPUT118), .B(n943), .ZN(n944) );
  NOR2_X1 U1035 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1036 ( .A1(n947), .A2(n946), .ZN(n958) );
  XNOR2_X1 U1037 ( .A(n948), .B(G1956), .ZN(n950) );
  XNOR2_X1 U1038 ( .A(G166), .B(G1971), .ZN(n949) );
  NAND2_X1 U1039 ( .A1(n950), .A2(n949), .ZN(n955) );
  NAND2_X1 U1040 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1041 ( .A(KEYINPUT119), .B(n953), .Z(n954) );
  NOR2_X1 U1042 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1043 ( .A(KEYINPUT120), .B(n956), .Z(n957) );
  NOR2_X1 U1044 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .ZN(n959) );
  XNOR2_X1 U1046 ( .A(KEYINPUT117), .B(n959), .ZN(n960) );
  NOR2_X1 U1047 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1048 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1049 ( .A(n964), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1050 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1051 ( .A(G120), .ZN(G236) );
  INV_X1 U1052 ( .A(G96), .ZN(G221) );
  INV_X1 U1053 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1054 ( .A1(n966), .A2(n965), .ZN(G325) );
  INV_X1 U1055 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1056 ( .A(n968), .B(n967), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(n969), .B(G286), .ZN(n972) );
  XNOR2_X1 U1058 ( .A(n970), .B(G171), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(n972), .B(n971), .ZN(n973) );
  NOR2_X1 U1060 ( .A1(G37), .A2(n973), .ZN(G397) );
  XOR2_X1 U1061 ( .A(G2678), .B(G2100), .Z(n975) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G2084), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1064 ( .A(n976), .B(KEYINPUT107), .Z(n978) );
  XNOR2_X1 U1065 ( .A(G2090), .B(KEYINPUT42), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(n978), .B(n977), .ZN(n982) );
  XOR2_X1 U1067 ( .A(G2096), .B(KEYINPUT43), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G2078), .B(G2072), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n980), .B(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(n982), .B(n981), .Z(G227) );
  XNOR2_X1 U1071 ( .A(G1986), .B(G1976), .ZN(n992) );
  XOR2_X1 U1072 ( .A(G1966), .B(G1971), .Z(n984) );
  XNOR2_X1 U1073 ( .A(G1996), .B(G1981), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n984), .B(n983), .ZN(n988) );
  XOR2_X1 U1075 ( .A(KEYINPUT108), .B(G2474), .Z(n986) );
  XNOR2_X1 U1076 ( .A(G1991), .B(G1961), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1078 ( .A(n988), .B(n987), .Z(n990) );
  XNOR2_X1 U1079 ( .A(G1956), .B(KEYINPUT41), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n992), .B(n991), .ZN(G229) );
  NAND2_X1 U1082 ( .A1(G118), .A2(n993), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(G130), .A2(n994), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1003) );
  NAND2_X1 U1085 ( .A1(G142), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(G106), .A2(n998), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1088 ( .A(n1001), .B(KEYINPUT45), .Z(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1005), .B(n1004), .ZN(n1013) );
  XOR2_X1 U1091 ( .A(KEYINPUT114), .B(KEYINPUT111), .Z(n1007) );
  XNOR2_X1 U1092 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1007), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(n1009), .B(n1008), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(G160), .B(G164), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1013), .B(n1012), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(n1014), .B(G162), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(n1020) );
  XNOR2_X1 U1100 ( .A(n1018), .B(n1017), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1102 ( .A1(G37), .A2(n1021), .ZN(G395) );
  NOR2_X1 U1103 ( .A1(G401), .A2(n1028), .ZN(n1025) );
  NOR2_X1 U1104 ( .A1(G227), .A2(G229), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(KEYINPUT49), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1106 ( .A1(G397), .A2(n1023), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1108 ( .A1(n1026), .A2(G395), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(n1027), .B(KEYINPUT115), .ZN(G225) );
  XOR2_X1 U1110 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1111 ( .A(n1028), .ZN(G319) );
  INV_X1 U1112 ( .A(G108), .ZN(G238) );
endmodule

