//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT21), .B(G898), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(G234), .A2(G237), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G902), .A3(G953), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n191), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G214), .B1(G237), .B2(G902), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT83), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT5), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G116), .ZN(new_n202));
  XNOR2_X1  g016(.A(G116), .B(G119), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(G113), .B(new_n202), .C1(new_n204), .C2(new_n200), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT84), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT2), .B(G113), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n203), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n206), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT78), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT78), .A2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT78), .B(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G107), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n216), .A2(KEYINPUT3), .A3(G107), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n221), .A2(new_n222), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n220), .B2(KEYINPUT3), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(KEYINPUT79), .A3(new_n222), .A4(new_n224), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n216), .A2(G107), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n222), .B1(new_n220), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n214), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  AOI211_X1 g050(.A(KEYINPUT80), .B(new_n234), .C1(new_n229), .C2(new_n231), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n213), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n222), .B1(new_n230), .B2(new_n224), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n229), .B2(new_n231), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n242), .B2(new_n239), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n209), .B1(new_n244), .B2(new_n203), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n204), .A2(KEYINPUT67), .A3(new_n208), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G110), .B(G122), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n238), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n205), .A2(new_n210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT86), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n234), .B1(new_n229), .B2(new_n231), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n249), .B(KEYINPUT85), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT8), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(new_n256), .C1(new_n253), .C2(new_n212), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .A4(G128), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT65), .B1(new_n258), .B2(G143), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n260), .A3(G146), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n264), .A2(new_n266), .B1(G143), .B2(new_n258), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n259), .B2(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  INV_X1    g085(.A(G125), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n259), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT0), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n268), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n275), .A3(new_n268), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n259), .A2(new_n261), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n274), .A2(new_n280), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n271), .B1(new_n272), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n187), .A2(G224), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n283), .B(new_n285), .Z(new_n286));
  NAND3_X1  g100(.A1(new_n250), .A2(new_n257), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n238), .A2(new_n248), .ZN(new_n292));
  INV_X1    g106(.A(new_n249), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT6), .A3(new_n250), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n283), .B(new_n284), .Z(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n288), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n291), .A2(new_n299), .A3(new_n302), .A4(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n199), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(G128), .B(G143), .Z(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G134), .ZN(new_n308));
  XNOR2_X1  g122(.A(G128), .B(G143), .ZN(new_n309));
  INV_X1    g123(.A(G134), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT14), .A3(G122), .ZN(new_n314));
  XOR2_X1   g128(.A(G116), .B(G122), .Z(new_n315));
  OAI211_X1 g129(.A(G107), .B(new_n314), .C1(new_n315), .C2(KEYINPUT14), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n315), .A2(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT95), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT13), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n260), .A3(G128), .ZN(new_n322));
  OAI211_X1 g136(.A(G134), .B(new_n322), .C1(new_n307), .C2(new_n321), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT93), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n315), .A2(G107), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n311), .B(KEYINPUT94), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT73), .B(G217), .Z(new_n330));
  XOR2_X1   g144(.A(KEYINPUT9), .B(G234), .Z(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n187), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n329), .B(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n288), .ZN(new_n334));
  INV_X1    g148(.A(G478), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(KEYINPUT15), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G475), .A2(G902), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT91), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n272), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(G125), .A2(G140), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n272), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n258), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n343), .ZN(new_n347));
  NOR2_X1   g161(.A1(G125), .A2(G140), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT16), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n345), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n346), .A2(KEYINPUT75), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n350), .A3(new_n353), .A4(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT89), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n357));
  NOR2_X1   g171(.A1(G237), .A2(G953), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G214), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n260), .ZN(new_n360));
  INV_X1    g174(.A(G131), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(G143), .A3(G214), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n360), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n357), .B2(new_n364), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n352), .A2(new_n367), .A3(new_n354), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(KEYINPUT18), .ZN(new_n370));
  NAND2_X1  g184(.A1(KEYINPUT18), .A2(G131), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n360), .A2(new_n362), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n342), .A2(new_n343), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n258), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(G113), .B(G122), .Z(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT88), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(G104), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n369), .A2(KEYINPUT90), .A3(new_n375), .A4(new_n378), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n373), .B(KEYINPUT19), .Z(new_n384));
  OAI221_X1 g198(.A(new_n351), .B1(new_n364), .B2(new_n363), .C1(new_n384), .C2(G146), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(new_n375), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n378), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n339), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  AOI211_X1 g203(.A(KEYINPUT91), .B(new_n387), .C1(new_n381), .C2(new_n382), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT20), .B(new_n338), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n387), .B1(new_n381), .B2(new_n382), .ZN(new_n393));
  INV_X1    g207(.A(new_n338), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n378), .B1(new_n369), .B2(new_n375), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n381), .B2(new_n382), .ZN(new_n397));
  OAI21_X1  g211(.A(G475), .B1(new_n397), .B2(G902), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT92), .A4(new_n398), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n306), .A2(new_n337), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G221), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n331), .B2(new_n288), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n187), .A2(G227), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n263), .B1(new_n281), .B2(new_n269), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n232), .A2(new_n235), .A3(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n243), .A2(new_n282), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n310), .B2(G137), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n310), .A2(G137), .ZN(new_n416));
  INV_X1    g230(.A(G137), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT11), .A3(G134), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT66), .A3(G131), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT66), .A2(G131), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n415), .A2(new_n418), .A3(new_n421), .A4(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(KEYINPUT10), .B(new_n270), .C1(new_n236), .C2(new_n237), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n413), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n413), .B2(new_n425), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n409), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT82), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(new_n409), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n426), .A2(new_n409), .ZN(new_n432));
  INV_X1    g246(.A(new_n412), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n253), .A2(new_n270), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT12), .B(new_n423), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n412), .B1(new_n253), .B2(new_n270), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n423), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT12), .A4(new_n423), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n429), .A2(new_n431), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n288), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n413), .A2(new_n424), .A3(new_n425), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n408), .B(KEYINPUT77), .ZN(new_n450));
  INV_X1    g264(.A(new_n427), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n449), .A2(new_n450), .B1(new_n432), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G469), .B1(new_n452), .B2(G902), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n405), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT23), .B1(new_n268), .B2(G119), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT74), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n201), .B2(G128), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT76), .B(G110), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G119), .B(G128), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT24), .B(G110), .Z(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n373), .A2(new_n258), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n351), .ZN(new_n465));
  INV_X1    g279(.A(G110), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n461), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n354), .A3(new_n352), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT22), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n417), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OR3_X1    g291(.A1(new_n477), .A2(KEYINPUT25), .A3(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n330), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(G234), .B2(new_n288), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT25), .B1(new_n477), .B2(G902), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n477), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT68), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT68), .B1(new_n245), .B2(new_n246), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n282), .A2(new_n423), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n419), .A2(G131), .ZN(new_n491));
  INV_X1    g305(.A(new_n416), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n310), .A2(G137), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n270), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(KEYINPUT30), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n501), .B2(new_n247), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT26), .B(G101), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n358), .A2(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT29), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g324(.A(new_n489), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n490), .A2(new_n495), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n490), .A2(new_n495), .B1(new_n245), .B2(new_n246), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT28), .B1(new_n497), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n508), .A2(new_n509), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n511), .B(new_n496), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n515), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n515), .B2(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(new_n507), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(new_n509), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n288), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G472), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n507), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n490), .A2(new_n499), .A3(new_n495), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n499), .B1(new_n490), .B2(new_n495), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n247), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n489), .A2(new_n496), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(KEYINPUT70), .A3(new_n533), .A4(new_n507), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n507), .B1(new_n516), .B2(new_n518), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT72), .B1(G472), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(KEYINPUT72), .A2(G472), .A3(G902), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n538), .B1(new_n529), .B2(new_n536), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT32), .B1(new_n548), .B2(new_n545), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n486), .B1(new_n528), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n454), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n403), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n222), .ZN(G3));
  NAND2_X1  g368(.A1(new_n447), .A2(new_n453), .ZN(new_n555));
  INV_X1    g369(.A(new_n405), .ZN(new_n556));
  INV_X1    g370(.A(new_n486), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n548), .A2(new_n545), .ZN(new_n558));
  INV_X1    g372(.A(G472), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n548), .A2(G902), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(KEYINPUT96), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n540), .A2(new_n288), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n558), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n333), .B(KEYINPUT33), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n568), .A2(new_n335), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n333), .A2(new_n335), .A3(new_n288), .ZN(new_n570));
  NAND2_X1  g384(.A1(G478), .A2(G902), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n401), .B2(new_n402), .ZN(new_n573));
  INV_X1    g387(.A(new_n197), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n574), .B(new_n195), .C1(new_n304), .C2(new_n305), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n567), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G104), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n576), .B(new_n578), .ZN(G6));
  AND2_X1   g393(.A1(new_n391), .A2(new_n398), .ZN(new_n580));
  INV_X1    g394(.A(new_n337), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n389), .A2(new_n390), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n392), .B1(new_n582), .B2(new_n394), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n567), .A2(new_n575), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G107), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n585), .B(new_n587), .ZN(G9));
  NOR2_X1   g402(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n470), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n484), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n593), .A2(new_n482), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n454), .A2(new_n565), .A3(new_n595), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n596), .A2(new_n403), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT37), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n466), .ZN(G12));
  NAND2_X1  g413(.A1(new_n528), .A2(new_n550), .ZN(new_n600));
  AND4_X1   g414(.A1(new_n556), .A2(new_n555), .A3(new_n600), .A4(new_n595), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n574), .B1(new_n304), .B2(new_n305), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G900), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n189), .B1(new_n194), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n580), .A2(new_n581), .A3(new_n583), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G128), .ZN(G30));
  NAND2_X1  g424(.A1(new_n401), .A2(new_n402), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(new_n581), .A3(new_n197), .A4(new_n594), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT101), .Z(new_n613));
  XOR2_X1   g427(.A(new_n605), .B(KEYINPUT39), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n454), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n615), .A2(KEYINPUT40), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n304), .A2(new_n305), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n521), .A2(new_n524), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n288), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n502), .A2(new_n524), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n541), .B1(new_n540), .B2(new_n546), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n548), .A2(KEYINPUT32), .A3(new_n545), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT100), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n550), .A2(new_n628), .A3(new_n623), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n615), .A2(KEYINPUT40), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n613), .A2(new_n616), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G143), .ZN(G45));
  AND3_X1   g449(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n611), .A2(new_n602), .A3(new_n636), .A4(new_n606), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT102), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n573), .A2(new_n639), .A3(new_n602), .A4(new_n606), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n601), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G146), .ZN(G48));
  INV_X1    g457(.A(new_n447), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n446), .B1(new_n445), .B2(new_n288), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n644), .A2(new_n645), .A3(new_n405), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(new_n573), .A3(new_n575), .A4(new_n551), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT41), .B(G113), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G15));
  NAND4_X1  g463(.A1(new_n646), .A2(new_n551), .A3(new_n575), .A4(new_n584), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT104), .B(G116), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G18));
  AND4_X1   g466(.A1(new_n337), .A2(new_n401), .A3(new_n402), .A4(new_n196), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n574), .B(new_n594), .C1(new_n304), .C2(new_n305), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n646), .A3(new_n654), .A4(new_n600), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G119), .ZN(G21));
  NAND2_X1  g470(.A1(new_n611), .A2(new_n581), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n445), .A2(new_n288), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(G469), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n556), .A3(new_n447), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n486), .A2(KEYINPUT106), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n537), .B1(new_n523), .B2(new_n507), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n545), .B(KEYINPUT105), .Z(new_n665));
  AOI22_X1  g479(.A1(new_n562), .A2(G472), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n486), .A2(KEYINPUT106), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n611), .A2(KEYINPUT107), .A3(new_n581), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n659), .A2(new_n669), .A3(new_n575), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  NAND2_X1  g486(.A1(new_n602), .A2(new_n595), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n662), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n611), .A2(new_n636), .A3(new_n606), .A4(new_n666), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G125), .ZN(G27));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT110), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n678), .A2(KEYINPUT110), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n304), .A2(new_n305), .A3(new_n197), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT109), .ZN(new_n682));
  NAND2_X1  g496(.A1(G469), .A2(G902), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT108), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n452), .B2(G469), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n405), .B1(new_n447), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n304), .A2(new_n688), .A3(new_n305), .A4(new_n197), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n682), .A2(new_n551), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n573), .A2(new_n606), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n679), .B(new_n680), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n682), .A2(new_n689), .A3(new_n687), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n611), .A2(new_n636), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n605), .ZN(new_n695));
  INV_X1    g509(.A(new_n600), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n663), .A2(new_n667), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n696), .A2(new_n697), .A3(new_n678), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n693), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n692), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G131), .ZN(G33));
  NOR2_X1   g515(.A1(new_n690), .A2(new_n607), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT111), .B(G134), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G36));
  NAND2_X1  g518(.A1(new_n449), .A2(new_n450), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n432), .A2(new_n451), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n452), .A2(KEYINPUT45), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(G469), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT46), .B1(new_n711), .B2(new_n684), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n644), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n684), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n556), .A3(new_n614), .ZN(new_n716));
  NOR2_X1   g530(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n636), .A2(new_n401), .A3(new_n402), .ZN(new_n718));
  NAND2_X1  g532(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n717), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n565), .A2(new_n594), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n716), .B1(new_n726), .B2(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n682), .A2(new_n689), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g543(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n723), .C2(new_n724), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n731), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n727), .B(new_n729), .C1(new_n730), .C2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G137), .ZN(G39));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  INV_X1    g550(.A(new_n714), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(new_n644), .A3(new_n712), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n738), .B2(new_n405), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n715), .A2(KEYINPUT47), .A3(new_n556), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n691), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n696), .A3(new_n486), .A4(new_n729), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  AOI22_X1  g557(.A1(new_n674), .A2(new_n675), .B1(new_n601), .B2(new_n608), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n593), .A2(new_n482), .A3(new_n606), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n630), .A2(new_n747), .A3(new_n687), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n602), .A3(new_n659), .A4(new_n670), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n749), .A3(new_n641), .A4(KEYINPUT52), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n749), .A3(new_n641), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n655), .A2(new_n647), .A3(new_n650), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n401), .A2(new_n581), .A3(new_n402), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n566), .B1(new_n694), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n553), .B1(new_n760), .B2(new_n306), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n761), .A3(new_n597), .A4(new_n671), .ZN(new_n762));
  INV_X1    g576(.A(new_n702), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n700), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n675), .A2(new_n687), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n580), .A2(new_n583), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT114), .A3(new_n337), .A4(new_n606), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n580), .A2(new_n337), .A3(new_n583), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n605), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(new_n454), .A3(new_n770), .A4(new_n600), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n594), .B(new_n728), .C1(new_n765), .C2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n762), .A2(new_n764), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT53), .B1(new_n757), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n756), .A2(new_n750), .ZN(new_n775));
  INV_X1    g589(.A(new_n553), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n694), .A2(new_n759), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n567), .A3(new_n306), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n776), .A2(new_n671), .A3(new_n597), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n702), .B1(new_n692), .B2(new_n699), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n771), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n595), .A3(new_n729), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n779), .A2(new_n780), .A3(new_n758), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n775), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT54), .B1(new_n774), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n722), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n189), .B(new_n669), .C1(new_n788), .C2(new_n720), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(new_n603), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n756), .B1(new_n751), .B2(new_n750), .ZN(new_n791));
  INV_X1    g605(.A(new_n753), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n773), .B(KEYINPUT53), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n785), .B1(new_n775), .B2(new_n783), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n787), .A2(new_n790), .A3(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n728), .A2(new_n630), .A3(new_n662), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n189), .A3(new_n557), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n573), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n189), .B(new_n729), .C1(new_n788), .C2(new_n720), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n696), .A2(new_n697), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n646), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT48), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(KEYINPUT48), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n188), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n801), .A2(new_n594), .A3(new_n662), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n666), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n619), .A2(new_n574), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n789), .A2(KEYINPUT50), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n810), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n723), .A2(new_n812), .A3(new_n189), .A4(new_n669), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT50), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n799), .A2(new_n401), .A3(new_n402), .A4(new_n572), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n809), .A2(new_n811), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n644), .A2(new_n645), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n405), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n739), .A2(new_n740), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n668), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n802), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT118), .B(KEYINPUT51), .C1(new_n816), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n808), .A2(new_n666), .B1(new_n813), .B2(KEYINPUT50), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n821), .A3(new_n811), .A4(new_n815), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n826), .B2(KEYINPUT118), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n800), .B(new_n807), .C1(new_n824), .C2(new_n827), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n797), .A2(new_n828), .B1(G952), .B2(G953), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n817), .B(KEYINPUT49), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n198), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n718), .A2(new_n405), .A3(new_n697), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n631), .A3(new_n619), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(G75));
  NAND2_X1  g648(.A1(new_n295), .A2(new_n297), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(new_n298), .Z(new_n836));
  XOR2_X1   g650(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n837));
  XNOR2_X1  g651(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(KEYINPUT120), .B2(KEYINPUT56), .ZN(new_n839));
  INV_X1    g653(.A(G210), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n840), .B(new_n288), .C1(new_n793), .C2(new_n794), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(KEYINPUT56), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n843));
  INV_X1    g657(.A(new_n839), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n793), .A2(new_n794), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(G902), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n843), .B(new_n844), .C1(new_n846), .C2(new_n840), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n187), .A2(G952), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n842), .A2(new_n847), .A3(new_n849), .ZN(G51));
  NAND2_X1  g664(.A1(new_n684), .A2(KEYINPUT57), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n684), .A2(KEYINPUT57), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n793), .A2(new_n795), .A3(new_n794), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n795), .B1(new_n793), .B2(new_n794), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n445), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n846), .A2(new_n711), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n848), .B1(new_n856), .B2(new_n857), .ZN(G54));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n845), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n582), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n848), .B1(new_n860), .B2(new_n582), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n863), .B(new_n288), .C1(new_n793), .C2(new_n794), .ZN(new_n864));
  INV_X1    g678(.A(new_n582), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(KEYINPUT121), .A3(G475), .A4(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n861), .A2(new_n862), .A3(new_n866), .ZN(G60));
  XOR2_X1   g681(.A(new_n571), .B(KEYINPUT59), .Z(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n568), .B(new_n869), .C1(new_n853), .C2(new_n854), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n787), .B2(new_n796), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n870), .B(new_n849), .C1(new_n871), .C2(new_n568), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(G63));
  NAND2_X1  g687(.A1(G217), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT60), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n845), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n848), .B1(new_n877), .B2(new_n477), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT122), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT123), .Z(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n793), .B2(new_n794), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n590), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(KEYINPUT122), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n878), .A2(new_n881), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n881), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n849), .B(new_n884), .C1(new_n882), .C2(new_n483), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n882), .A2(new_n590), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(G66));
  AOI21_X1  g704(.A(new_n187), .B1(new_n190), .B2(G224), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n762), .B2(new_n187), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n835), .B1(G898), .B2(new_n187), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n892), .B(new_n893), .Z(G69));
  AOI21_X1  g708(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n501), .B(new_n384), .Z(new_n896));
  NAND2_X1  g710(.A1(G900), .A2(G953), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n744), .A2(new_n641), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n716), .A2(new_n696), .A3(new_n697), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n659), .A2(new_n602), .A3(new_n670), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n764), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n734), .A2(new_n742), .A3(new_n898), .A4(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n896), .B(new_n897), .C1(new_n902), .C2(G953), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n634), .A2(new_n898), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n634), .A2(KEYINPUT62), .A3(new_n898), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n777), .A2(new_n551), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n910), .A2(new_n615), .A3(new_n728), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT124), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n734), .A3(new_n742), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n896), .B1(new_n913), .B2(new_n187), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n895), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n895), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n913), .A2(new_n187), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n903), .C1(new_n917), .C2(new_n896), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(G72));
  XNOR2_X1  g733(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n559), .A2(new_n288), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n920), .B(new_n921), .Z(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n913), .B2(new_n762), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n848), .B1(new_n923), .B2(new_n622), .ZN(new_n924));
  INV_X1    g738(.A(new_n922), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n502), .A2(new_n507), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n508), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT126), .Z(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n774), .B2(new_n786), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n922), .B1(new_n902), .B2(new_n762), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n524), .A3(new_n502), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n924), .A2(new_n929), .A3(new_n931), .ZN(G57));
endmodule


