//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n465), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT69), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n475), .A2(new_n463), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(G136), .B2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n463), .A2(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(new_n484), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n489));
  INV_X1    g064(.A(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n463), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n485), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n488), .A2(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .A3(new_n485), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(new_n511), .B1(G75), .B2(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(KEYINPUT72), .A3(G62), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n509), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n514), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(new_n518), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(new_n531), .B1(new_n507), .B2(new_n508), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n518), .A2(G52), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n506), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n520), .A2(new_n509), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G81), .B1(G43), .B2(new_n518), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n545), .A2(KEYINPUT75), .A3(G91), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n521), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n518), .A2(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n518), .A2(new_n559), .A3(G53), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n553), .A2(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n509), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n507), .A2(KEYINPUT76), .A3(new_n508), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(G78), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n561), .A2(new_n568), .ZN(G299));
  XNOR2_X1  g144(.A(G168), .B(KEYINPUT77), .ZN(G286));
  OR2_X1    g145(.A1(new_n514), .A2(new_n523), .ZN(G303));
  NAND2_X1  g146(.A1(new_n545), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n507), .B2(new_n508), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n579), .B2(new_n506), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(G48), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n520), .A2(new_n509), .A3(G86), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n584), .B(G651), .C1(new_n577), .C2(new_n578), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n583), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n506), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n518), .A2(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n521), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n520), .A2(new_n509), .A3(G92), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n527), .B2(KEYINPUT79), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(KEYINPUT79), .B2(new_n527), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n564), .B2(new_n565), .ZN(new_n602));
  AND2_X1   g177(.A1(G79), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT80), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G321));
  NOR2_X1   g183(.A1(G299), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G286), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  AOI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n481), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n476), .A2(G123), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n621), .A2(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n622), .B2(new_n621), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n619), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT82), .B(G2096), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n490), .A2(G2105), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n493), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n642), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2100), .Z(new_n661));
  NOR2_X1   g236(.A1(G2072), .A2(G2078), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n442), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2096), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G29), .A2(G35), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G162), .B2(G29), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(G2090), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT97), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n606), .A2(G16), .ZN(new_n691));
  NOR2_X1   g266(.A1(G4), .A2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT90), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G1348), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G27), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT95), .Z(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G164), .B2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(G2078), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT26), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n706), .A2(new_n707), .B1(G105), .B2(new_n629), .ZN(new_n708));
  INV_X1    g283(.A(new_n476), .ZN(new_n709));
  INV_X1    g284(.A(G129), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n475), .A2(new_n463), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n713));
  INV_X1    g288(.A(G141), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n698), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n698), .B2(G32), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n703), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n723), .B2(KEYINPUT24), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(KEYINPUT24), .B2(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(G160), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n698), .ZN(new_n727));
  INV_X1    g302(.A(G2084), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n547), .A2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G16), .B2(G19), .ZN(new_n731));
  INV_X1    g306(.A(G1341), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n731), .A2(new_n732), .B1(new_n698), .B2(new_n626), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n729), .B(new_n733), .C1(new_n732), .C2(new_n731), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G5), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G171), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT31), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G11), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G11), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n698), .B1(new_n743), .B2(G28), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n741), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n727), .B2(new_n728), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n734), .A2(new_n739), .A3(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n722), .B(new_n748), .C1(G2090), .C2(new_n688), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n720), .A2(new_n721), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n735), .A2(G20), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1956), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n698), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  OAI21_X1  g331(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n757));
  INV_X1    g332(.A(G116), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G2105), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n476), .B2(G128), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n481), .A2(G140), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n735), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n735), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT94), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1966), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n750), .A2(new_n754), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n698), .A2(G33), .B1(KEYINPUT92), .B2(G2072), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n463), .ZN(new_n772));
  INV_X1    g347(.A(G139), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n712), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT25), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT91), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n778));
  INV_X1    g353(.A(new_n776), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n778), .B(new_n779), .C1(new_n712), .C2(new_n773), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n772), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n770), .B1(new_n781), .B2(new_n698), .ZN(new_n782));
  NOR2_X1   g357(.A1(KEYINPUT92), .A2(G2072), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n782), .B(new_n783), .Z(new_n784));
  NOR2_X1   g359(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n697), .A2(new_n749), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n735), .A2(G22), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT87), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G303), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  OR2_X1    g365(.A1(G6), .A2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G305), .B2(new_n735), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n789), .A2(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n790), .B2(new_n789), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n735), .A2(G23), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n735), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n792), .B2(new_n793), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n795), .A2(new_n801), .A3(KEYINPUT34), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT34), .B1(new_n795), .B2(new_n801), .ZN(new_n803));
  OR2_X1    g378(.A1(G25), .A2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n481), .A2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n476), .A2(G119), .ZN(new_n806));
  OR2_X1    g381(.A1(G95), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n804), .B1(new_n809), .B2(new_n698), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n735), .A2(G24), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n592), .B2(new_n735), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1986), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n802), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT89), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT88), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n821), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n786), .B1(new_n822), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n822), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n825), .A2(new_n697), .A3(new_n749), .A4(new_n785), .ZN(G150));
  NAND2_X1  g401(.A1(new_n606), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n545), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n506), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n547), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n828), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n831), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(KEYINPUT101), .B(G37), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n781), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n762), .A2(new_n499), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n760), .A2(new_n485), .A3(new_n502), .A4(new_n761), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n781), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n849), .A3(new_n718), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n718), .B1(new_n847), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n481), .A2(G142), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT99), .Z(new_n854));
  INV_X1    g429(.A(new_n631), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n809), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(G130), .ZN(new_n860));
  OR3_X1    g435(.A1(new_n709), .A2(KEYINPUT100), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT100), .B1(new_n709), .B2(new_n860), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n809), .A2(new_n855), .ZN(new_n864));
  AND4_X1   g439(.A1(new_n854), .A2(new_n856), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n863), .A2(new_n854), .B1(new_n856), .B2(new_n864), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n851), .A2(new_n852), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n847), .A2(new_n849), .ZN(new_n869));
  INV_X1    g444(.A(new_n718), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n850), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n626), .B(new_n726), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(G162), .Z(new_n875));
  AOI21_X1  g450(.A(new_n843), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(KEYINPUT102), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n868), .A2(new_n871), .A3(new_n878), .A4(new_n850), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n877), .A2(new_n879), .A3(new_n867), .A4(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n876), .A2(new_n881), .A3(KEYINPUT103), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT103), .B1(new_n876), .B2(new_n881), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n876), .A2(new_n881), .A3(KEYINPUT103), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT40), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n885), .A2(new_n890), .ZN(G395));
  XNOR2_X1  g466(.A(G166), .B(KEYINPUT104), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G305), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n797), .B(new_n592), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G305), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n892), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n899), .A3(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n605), .ZN(new_n908));
  INV_X1    g483(.A(G299), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n605), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n615), .B(new_n833), .ZN(new_n917));
  MUX2_X1   g492(.A(new_n916), .B(new_n912), .S(new_n917), .Z(new_n918));
  AND2_X1   g493(.A1(new_n907), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n907), .A2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G868), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n831), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n923), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  INV_X1    g501(.A(G168), .ZN(new_n927));
  NAND2_X1  g502(.A1(G301), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G301), .B2(G286), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(new_n833), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n913), .B2(new_n915), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n929), .B(new_n832), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n911), .A3(new_n910), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n895), .A2(new_n899), .A3(KEYINPUT105), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT105), .B1(new_n895), .B2(new_n899), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n931), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n932), .B1(new_n939), .B2(new_n915), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n936), .B(new_n842), .C1(new_n941), .C2(new_n904), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n926), .B1(new_n942), .B2(KEYINPUT43), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n931), .A2(new_n933), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n902), .A3(new_n903), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n936), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(KEYINPUT108), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT108), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(new_n944), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n904), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n946), .B1(new_n955), .B2(new_n945), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n951), .A2(new_n957), .ZN(G397));
  INV_X1    g533(.A(G2067), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n762), .B(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT111), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n718), .ZN(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G125), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n491), .B2(new_n492), .ZN(new_n966));
  INV_X1    g541(.A(new_n467), .ZN(new_n967));
  OAI21_X1  g542(.A(G2105), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n470), .B1(new_n969), .B2(G137), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n970), .A3(G40), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT109), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND3_X1  g548(.A1(G160), .A2(new_n973), .A3(G40), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  AND2_X1   g551(.A1(G126), .A2(G2105), .ZN(new_n977));
  INV_X1    g552(.A(G138), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G2105), .ZN(new_n979));
  INV_X1    g554(.A(new_n484), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n498), .B1(new_n981), .B2(new_n474), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n969), .B2(G138), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n975), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n962), .A2(new_n964), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n963), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT110), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(new_n870), .ZN(new_n991));
  INV_X1    g566(.A(new_n811), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n809), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n809), .A2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1986), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n592), .B(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n987), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(G166), .B2(new_n1001), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n502), .A2(KEYINPUT71), .A3(new_n485), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT71), .B1(new_n502), .B2(new_n485), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n976), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1010));
  NAND3_X1  g585(.A1(new_n499), .A2(new_n976), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT113), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n502), .B2(new_n485), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n1010), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G2090), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n973), .B1(G160), .B2(G40), .ZN(new_n1018));
  AND4_X1   g593(.A1(new_n973), .A2(new_n968), .A3(new_n970), .A4(G40), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1009), .A2(new_n1016), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1008), .A2(new_n985), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n972), .A2(new_n974), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1021), .A2(new_n1022), .B1(new_n1026), .B2(new_n790), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n975), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(KEYINPUT114), .A3(new_n1017), .A4(new_n1009), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1001), .B(new_n1005), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G305), .A2(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n580), .A2(new_n583), .A3(new_n1032), .A4(new_n585), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n972), .A2(new_n974), .A3(new_n1013), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n797), .A2(G1976), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1039), .A3(G8), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1037), .A2(new_n1038), .B1(KEYINPUT52), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1035), .A2(new_n1039), .A3(new_n1043), .A4(G8), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n504), .B2(new_n976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n972), .A2(new_n974), .A3(new_n1024), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n790), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n504), .A2(new_n1050), .A3(new_n976), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1013), .A2(new_n1010), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1017), .A3(new_n1020), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1001), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1041), .B(new_n1045), .C1(new_n1046), .C2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1000), .B1(new_n1030), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(G8), .A3(new_n1046), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1054), .A2(new_n1046), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1058), .A2(new_n1059), .A3(KEYINPUT126), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1026), .B2(G2078), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1009), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n738), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n986), .A2(new_n1067), .A3(new_n972), .A4(new_n974), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n986), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT116), .B1(new_n1071), .B2(new_n975), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n702), .A2(KEYINPUT53), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1064), .B(new_n1066), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1056), .A2(new_n1062), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1067), .B1(new_n1020), .B2(new_n986), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT117), .B(G2084), .Z(new_n1082));
  NAND3_X1  g657(.A1(new_n1028), .A2(new_n1009), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(G168), .A3(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(KEYINPUT125), .A2(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(KEYINPUT51), .A3(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1966), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1082), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1065), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(G8), .B(new_n927), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT124), .A3(G8), .A4(new_n927), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1090), .A2(KEYINPUT62), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT62), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1077), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT127), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1077), .B(new_n1104), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1035), .A2(G2067), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1065), .B2(new_n695), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(KEYINPUT122), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1110), .B(new_n1107), .C1(new_n1065), .C2(new_n695), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n558), .A2(new_n560), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT120), .B1(new_n558), .B2(new_n560), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT121), .B1(new_n1119), .B2(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G299), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n909), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1051), .A2(new_n1020), .A3(new_n1052), .ZN(new_n1128));
  INV_X1    g703(.A(G1956), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1124), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1112), .A2(new_n908), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1124), .A2(KEYINPUT123), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1122), .A2(new_n1123), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n908), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1109), .A2(new_n1111), .A3(KEYINPUT60), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1131), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1124), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1124), .B1(new_n1130), .B2(new_n1127), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT60), .B(new_n605), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1026), .A2(G1996), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT58), .B(G1341), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n547), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n547), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1138), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1159));
  XNOR2_X1  g734(.A(G301), .B(KEYINPUT54), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1071), .A2(new_n971), .A3(new_n1074), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1024), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1075), .A2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1158), .A2(new_n1159), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1097), .A2(G8), .A3(new_n610), .ZN(new_n1168));
  OR3_X1    g743(.A1(new_n1030), .A2(new_n1055), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1057), .A2(G8), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1005), .A2(KEYINPUT119), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1168), .A2(new_n1177), .A3(new_n1171), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1030), .A2(new_n1055), .A3(new_n1168), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT118), .B1(new_n1180), .B2(KEYINPUT63), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1172), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1183), .A2(new_n1042), .A3(new_n797), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1036), .B1(new_n1184), .B2(new_n1033), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n1030), .B2(new_n1059), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1167), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n999), .B1(new_n1106), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n987), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n990), .B(KEYINPUT46), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT47), .Z(new_n1192));
  NAND3_X1  g767(.A1(new_n988), .A2(new_n991), .A3(new_n994), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n760), .A2(new_n959), .A3(new_n761), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n975), .B(new_n986), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n987), .A2(new_n997), .A3(new_n592), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT48), .Z(new_n1197));
  NOR2_X1   g772(.A1(new_n996), .A2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1192), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1188), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g775(.A1(new_n953), .A2(new_n956), .ZN(new_n1202));
  OAI21_X1  g776(.A(G319), .B1(new_n650), .B2(new_n651), .ZN(new_n1203));
  NOR3_X1   g777(.A1(G229), .A2(G227), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1204), .B1(new_n882), .B2(new_n883), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1202), .A2(new_n1205), .ZN(G308));
  OAI221_X1 g780(.A(new_n1204), .B1(new_n882), .B2(new_n883), .C1(new_n953), .C2(new_n956), .ZN(G225));
endmodule


