//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AOI211_X1 g043(.A(new_n467), .B(new_n468), .C1(new_n463), .C2(new_n464), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G137), .A4(new_n468), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n461), .A2(new_n462), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT70), .Z(new_n486));
  NOR2_X1   g061(.A1(new_n483), .A2(new_n468), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n482), .B(new_n486), .C1(G124), .C2(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G138), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n474), .A2(KEYINPUT4), .A3(G138), .A4(new_n468), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n474), .A2(G126), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(G50), .A3(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n508), .A2(new_n500), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n503), .A2(new_n511), .A3(new_n513), .ZN(G166));
  AND2_X1   g089(.A1(G63), .A2(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n518), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n508), .A2(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(new_n500), .A3(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n498), .A2(KEYINPUT73), .A3(new_n499), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(new_n526), .A3(G543), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n520), .B(new_n521), .C1(new_n527), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND4_X1  g105(.A1(new_n522), .A2(new_n526), .A3(G52), .A4(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n508), .A2(new_n500), .A3(G90), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n510), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n506), .B2(new_n507), .ZN(new_n537));
  AND2_X1   g112(.A1(G68), .A2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G81), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n508), .A2(new_n500), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n539), .B(new_n541), .C1(new_n542), .C2(new_n527), .ZN(new_n543));
  INV_X1    g118(.A(G860), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT9), .B1(new_n527), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n505), .B1(new_n500), .B2(new_n523), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n552), .A2(new_n553), .A3(G53), .A4(new_n522), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n506), .A2(new_n507), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n512), .B2(G91), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n555), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(G299));
  NAND3_X1  g138(.A1(new_n503), .A2(new_n511), .A3(new_n513), .ZN(G303));
  OAI21_X1  g139(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n508), .A2(new_n500), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n522), .A2(new_n526), .A3(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(KEYINPUT76), .A3(G49), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n527), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n568), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(G288));
  NAND2_X1  g150(.A1(new_n512), .A2(G86), .ZN(new_n576));
  AND2_X1   g151(.A1(G48), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT78), .B1(new_n500), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n500), .A2(KEYINPUT78), .A3(new_n577), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n510), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n583), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n580), .A2(new_n578), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n576), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n522), .A2(new_n526), .A3(G47), .A4(G543), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n508), .A2(new_n500), .A3(G85), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n592), .A2(new_n591), .A3(new_n593), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n557), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n506), .B2(new_n507), .ZN(new_n602));
  INV_X1    g177(.A(new_n599), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT80), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(G651), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT82), .B1(new_n597), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n592), .A2(new_n593), .A3(new_n591), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n605), .B(KEYINPUT82), .C1(new_n607), .C2(new_n594), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n506), .B2(new_n507), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n614), .A2(KEYINPUT83), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT83), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n617), .A2(G651), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n567), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n569), .A2(G54), .ZN(new_n625));
  AND3_X1   g200(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n612), .B1(new_n626), .B2(G868), .ZN(G284));
  XOR2_X1   g202(.A(G284), .B(KEYINPUT84), .Z(G321));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(G299), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(G168), .ZN(G297));
  XOR2_X1   g206(.A(G297), .B(KEYINPUT85), .Z(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n543), .A2(new_n629), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n635), .B1(new_n637), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g214(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n643), .A2(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n484), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n487), .A2(G123), .ZN(new_n647));
  OR2_X1    g222(.A1(G99), .A2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n648), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(G2100), .B2(new_n643), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT89), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2451), .B(G2454), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT90), .Z(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(G2100), .Z(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(G2096), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n689), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n691), .B(new_n694), .C1(new_n686), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G35), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G162), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT29), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G2090), .ZN(new_n707));
  MUX2_X1   g282(.A(G19), .B(new_n543), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1341), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n703), .A2(G33), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n474), .A2(G127), .ZN(new_n711));
  AND2_X1   g286(.A1(G115), .A2(G2104), .ZN(new_n712));
  OAI21_X1  g287(.A(G2105), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT25), .ZN(new_n714));
  NAND2_X1  g289(.A1(G103), .A2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G2105), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n484), .A2(G139), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n710), .B1(new_n719), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2072), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n650), .A2(new_n703), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n725), .A2(new_n703), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n703), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n703), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2078), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n707), .A2(new_n709), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G20), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT23), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G299), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1956), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n703), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(KEYINPUT26), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n484), .A2(G141), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT99), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n739), .B1(new_n749), .B2(new_n703), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT100), .Z(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT101), .B1(G16), .B2(G21), .ZN(new_n755));
  NAND2_X1  g330(.A1(G168), .A2(G16), .ZN(new_n756));
  MUX2_X1   g331(.A(KEYINPUT101), .B(new_n755), .S(new_n756), .Z(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n703), .A2(G26), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT28), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n484), .A2(G140), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(G116), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G2105), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n487), .B2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NOR2_X1   g346(.A1(G171), .A2(new_n734), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G5), .B2(new_n734), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G1961), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n754), .A2(new_n759), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n703), .B1(KEYINPUT24), .B2(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(KEYINPUT24), .B2(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n478), .B2(G29), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n777), .A2(new_n780), .B1(new_n774), .B2(G1961), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n781), .B1(new_n758), .B2(new_n757), .C1(new_n752), .C2(new_n753), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n777), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT98), .ZN(new_n785));
  NOR2_X1   g360(.A1(G4), .A2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT96), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n636), .B2(new_n734), .ZN(new_n788));
  INV_X1    g363(.A(G1348), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n733), .A2(new_n738), .A3(new_n783), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n574), .A2(new_n734), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n734), .B2(G23), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT33), .B(G1976), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n734), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n734), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(G1971), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n734), .A2(G6), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n589), .B2(new_n734), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT32), .B(G1981), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n803), .A2(new_n805), .B1(new_n794), .B2(new_n795), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n803), .A2(new_n805), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n801), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n811));
  NOR2_X1   g386(.A1(G25), .A2(G29), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n484), .A2(G131), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n487), .A2(G119), .ZN(new_n814));
  INV_X1    g389(.A(G95), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n815), .A2(new_n468), .A3(KEYINPUT92), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT92), .B1(new_n815), .B2(new_n468), .ZN(new_n817));
  OAI221_X1 g392(.A(G2104), .B1(G107), .B2(new_n468), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n813), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n812), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT93), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n610), .A2(G16), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G16), .B2(G24), .ZN(new_n825));
  INV_X1    g400(.A(G1986), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n810), .A2(new_n811), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n811), .B1(new_n810), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n792), .B1(new_n835), .B2(new_n837), .ZN(G311));
  INV_X1    g413(.A(G311), .ZN(G150));
  NAND2_X1  g414(.A1(new_n626), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT103), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n522), .A2(new_n526), .A3(G55), .A4(G543), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT102), .B(G93), .Z(new_n844));
  NAND3_X1  g419(.A1(new_n844), .A2(new_n508), .A3(new_n500), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n845), .C1(new_n846), .C2(new_n510), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n543), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n543), .A2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n842), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  NOR2_X1   g433(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n769), .B(G164), .ZN(new_n860));
  INV_X1    g435(.A(new_n749), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n487), .A2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n468), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n484), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n641), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n819), .ZN(new_n872));
  XNOR2_X1  g447(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n865), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n478), .B(new_n650), .ZN(new_n878));
  XOR2_X1   g453(.A(G162), .B(new_n878), .Z(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n875), .A2(new_n879), .A3(new_n876), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g460(.A1(new_n847), .A2(new_n629), .ZN(new_n886));
  AND3_X1   g461(.A1(G166), .A2(new_n584), .A3(new_n588), .ZN(new_n887));
  AOI21_X1  g462(.A(G166), .B1(new_n584), .B2(new_n588), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n605), .B1(new_n607), .B2(new_n594), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT82), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n892), .A2(new_n574), .A3(new_n608), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n574), .B1(new_n892), .B2(new_n608), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT107), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n570), .A2(new_n573), .ZN(new_n896));
  INV_X1    g471(.A(new_n568), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n606), .B2(new_n609), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n574), .A3(new_n608), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n889), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n887), .A2(new_n888), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(KEYINPUT107), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n851), .B(new_n637), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n636), .B1(new_n561), .B2(new_n562), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n555), .A2(new_n560), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT75), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n560), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n626), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n910), .A2(new_n915), .A3(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n918), .B1(new_n909), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n908), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n886), .B1(new_n924), .B2(new_n629), .ZN(G295));
  OAI21_X1  g500(.A(new_n886), .B1(new_n924), .B2(new_n629), .ZN(G331));
  XOR2_X1   g501(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n927));
  AND3_X1   g502(.A1(new_n910), .A2(new_n915), .A3(KEYINPUT41), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(new_n910), .B2(new_n915), .ZN(new_n929));
  NOR2_X1   g504(.A1(G301), .A2(G286), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G301), .A2(G286), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n849), .A2(new_n931), .A3(new_n850), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n850), .ZN(new_n934));
  AND2_X1   g509(.A1(G301), .A2(G286), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n934), .A2(new_n848), .B1(new_n935), .B2(new_n930), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n932), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n851), .B2(new_n939), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n928), .A2(new_n929), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n936), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n910), .B2(new_n915), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n907), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n938), .ZN(new_n947));
  INV_X1    g522(.A(new_n940), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n943), .B1(new_n922), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n951), .C1(new_n903), .C2(new_n906), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n949), .B2(new_n917), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n922), .A2(new_n942), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT112), .A4(new_n916), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n907), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n907), .B2(new_n945), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n954), .B1(new_n953), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(KEYINPUT111), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  AOI211_X1 g540(.A(new_n965), .B(new_n954), .C1(new_n953), .C2(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n927), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n953), .A2(new_n960), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n953), .A2(new_n954), .A3(new_n962), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(KEYINPUT44), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n970), .A2(KEYINPUT114), .A3(KEYINPUT44), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n927), .C1(new_n964), .C2(new_n966), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n968), .A2(new_n976), .A3(new_n978), .ZN(G397));
  OAI211_X1 g554(.A(new_n477), .B(G40), .C1(new_n466), .C2(new_n469), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n496), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n769), .A2(G2067), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n769), .A2(G2067), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(new_n749), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT46), .B1(new_n984), .B2(G1996), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n984), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n992));
  XNOR2_X1  g567(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n984), .A2(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n749), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT115), .Z(new_n996));
  INV_X1    g571(.A(new_n984), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n987), .B1(new_n998), .B2(new_n749), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n819), .A2(new_n821), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n984), .B1(new_n1002), .B2(new_n985), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n819), .A2(new_n821), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n997), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n997), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT48), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n993), .B(new_n1003), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT126), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1981), .B1(new_n581), .B2(new_n583), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n585), .A2(new_n586), .A3(new_n1013), .A4(new_n576), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1012), .A2(new_n1014), .A3(KEYINPUT49), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT49), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n496), .A2(new_n982), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n980), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G288), .A2(G1976), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT120), .B1(new_n1022), .B2(new_n1014), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1018), .B(KEYINPUT119), .Z(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(KEYINPUT120), .A3(new_n1014), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n574), .A2(KEYINPUT118), .A3(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT118), .B1(new_n574), .B2(G1976), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1018), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1019), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1031), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT52), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G303), .A2(G8), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT55), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n980), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1017), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT116), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n983), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1971), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n496), .A2(new_n1049), .A3(new_n982), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n496), .A2(KEYINPUT117), .A3(new_n1049), .A4(new_n982), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1049), .B1(new_n496), .B2(new_n982), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n980), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2090), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1038), .B(G8), .C1(new_n1048), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1025), .A2(new_n1026), .B1(new_n1035), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1056), .A2(new_n1050), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G2090), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1064), .A2(new_n1065), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1037), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1059), .A2(new_n1068), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1039), .A2(new_n980), .A3(new_n983), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(G1966), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1054), .A2(new_n777), .A3(new_n1056), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n981), .A2(new_n1042), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(KEYINPUT121), .A3(new_n758), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G8), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G286), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1062), .B1(new_n1069), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1048), .B2(new_n1058), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1062), .B1(new_n1082), .B2(new_n1037), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1035), .A2(new_n1083), .A3(new_n1059), .A4(new_n1079), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1061), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1063), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n911), .B(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1040), .A2(new_n1043), .A3(new_n1045), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1057), .A2(new_n789), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n980), .A2(G2067), .A3(new_n1017), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n636), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n626), .B(new_n1096), .C1(new_n1057), .C2(new_n789), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1099), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1091), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1103), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n636), .A2(KEYINPUT60), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1095), .A2(new_n1097), .A3(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1040), .A2(new_n1043), .A3(new_n998), .A4(new_n1045), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n980), .B2(new_n1017), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n543), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(KEYINPUT59), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(KEYINPUT59), .B2(new_n1117), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1101), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  INV_X1    g697(.A(G2078), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1040), .A2(new_n1043), .A3(new_n1123), .A4(new_n1045), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT123), .B(G1961), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1057), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n465), .B2(G2105), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1042), .A2(new_n1130), .A3(new_n477), .A4(new_n1074), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1126), .A2(G301), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1122), .B1(new_n1132), .B2(KEYINPUT124), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(KEYINPUT124), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1124), .A2(new_n1125), .B1(new_n1057), .B2(new_n1127), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n1123), .ZN(new_n1137));
  AOI21_X1  g712(.A(G301), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1133), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(G286), .A2(G8), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1077), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1078), .A2(new_n1141), .A3(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(G8), .B(new_n1147), .C1(new_n1077), .C2(G286), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1144), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1136), .A2(G301), .A3(new_n1137), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(KEYINPUT54), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1140), .A2(new_n1151), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1150), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1142), .B(new_n1147), .C1(new_n1077), .C2(G8), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1143), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1139), .B1(new_n1160), .B2(KEYINPUT62), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1151), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1121), .A2(new_n1157), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1069), .B(KEYINPUT125), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1087), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n610), .A2(new_n826), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n997), .B1(new_n1007), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1006), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1011), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1132), .A2(KEYINPUT124), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1173), .B(new_n1122), .C1(new_n1138), .C2(new_n1134), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n1160), .A3(new_n1155), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1138), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1176));
  AOI211_X1 g751(.A(KEYINPUT62), .B(new_n1144), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1175), .A2(new_n1120), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1086), .B1(new_n1178), .B2(new_n1165), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1179), .A2(KEYINPUT126), .A3(new_n1170), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1010), .B1(new_n1172), .B2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g756(.A(G227), .ZN(new_n1183));
  NAND2_X1  g757(.A1(G319), .A2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g758(.A1(G229), .A2(new_n670), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n884), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n964), .A2(new_n966), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1186), .A2(new_n1187), .ZN(G308));
  OR2_X1    g762(.A1(new_n1186), .A2(new_n1187), .ZN(G225));
endmodule


