

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U555 ( .A1(G101), .A2(n561), .ZN(n537) );
  AND2_X1 U556 ( .A1(n724), .A2(n723), .ZN(n524) );
  NAND2_X1 U557 ( .A1(G286), .A2(G8), .ZN(n525) );
  NOR2_X1 U558 ( .A1(n759), .A2(n769), .ZN(n526) );
  NOR2_X1 U559 ( .A1(n811), .A2(n528), .ZN(n527) );
  AND2_X1 U560 ( .A1(n984), .A2(n822), .ZN(n528) );
  INV_X1 U561 ( .A(G168), .ZN(n723) );
  NAND2_X1 U562 ( .A1(G8), .A2(n730), .ZN(n769) );
  NOR2_X1 U563 ( .A1(G651), .A2(n614), .ZN(n650) );
  XNOR2_X1 U564 ( .A(n542), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  XOR2_X2 U566 ( .A(KEYINPUT68), .B(n529), .Z(n863) );
  NAND2_X1 U567 ( .A1(n863), .A2(G113), .ZN(n541) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X1 U569 ( .A(KEYINPUT17), .B(n530), .Z(n681) );
  NAND2_X1 U570 ( .A1(n681), .A2(G137), .ZN(n534) );
  INV_X1 U571 ( .A(G2105), .ZN(n531) );
  NOR2_X1 U572 ( .A1(n531), .A2(G2104), .ZN(n532) );
  XNOR2_X2 U573 ( .A(n532), .B(KEYINPUT66), .ZN(n862) );
  NAND2_X1 U574 ( .A1(G125), .A2(n862), .ZN(n533) );
  NAND2_X1 U575 ( .A1(n534), .A2(n533), .ZN(n539) );
  NAND2_X1 U576 ( .A1(n531), .A2(G2104), .ZN(n535) );
  XNOR2_X1 U577 ( .A(n535), .B(KEYINPUT67), .ZN(n561) );
  INV_X1 U578 ( .A(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U579 ( .A(n537), .B(n536), .ZN(n538) );
  NOR2_X1 U580 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U581 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n543) );
  XNOR2_X1 U583 ( .A(n543), .B(KEYINPUT64), .ZN(n655) );
  NAND2_X1 U584 ( .A1(G89), .A2(n655), .ZN(n544) );
  XNOR2_X1 U585 ( .A(n544), .B(KEYINPUT4), .ZN(n547) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n545) );
  XNOR2_X1 U587 ( .A(KEYINPUT70), .B(n545), .ZN(n614) );
  XNOR2_X1 U588 ( .A(G651), .B(KEYINPUT71), .ZN(n549) );
  NOR2_X1 U589 ( .A1(n614), .A2(n549), .ZN(n654) );
  NAND2_X1 U590 ( .A1(G76), .A2(n654), .ZN(n546) );
  NAND2_X1 U591 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U592 ( .A(KEYINPUT5), .B(n548), .ZN(n557) );
  NAND2_X1 U593 ( .A1(n650), .A2(G51), .ZN(n553) );
  NOR2_X1 U594 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n550), .Z(n551) );
  XNOR2_X1 U596 ( .A(KEYINPUT72), .B(n551), .ZN(n651) );
  NAND2_X1 U597 ( .A1(G63), .A2(n651), .ZN(n552) );
  NAND2_X1 U598 ( .A1(n553), .A2(n552), .ZN(n555) );
  XOR2_X1 U599 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n554) );
  XNOR2_X1 U600 ( .A(n555), .B(n554), .ZN(n556) );
  NAND2_X1 U601 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(n558), .ZN(G168) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U604 ( .A1(n862), .A2(G123), .ZN(n559) );
  XNOR2_X1 U605 ( .A(n559), .B(KEYINPUT76), .ZN(n560) );
  XNOR2_X1 U606 ( .A(n560), .B(KEYINPUT18), .ZN(n563) );
  BUF_X1 U607 ( .A(n561), .Z(n858) );
  NAND2_X1 U608 ( .A1(G99), .A2(n858), .ZN(n562) );
  NAND2_X1 U609 ( .A1(n563), .A2(n562), .ZN(n567) );
  BUF_X1 U610 ( .A(n681), .Z(n859) );
  NAND2_X1 U611 ( .A1(G135), .A2(n859), .ZN(n565) );
  NAND2_X1 U612 ( .A1(G111), .A2(n863), .ZN(n564) );
  NAND2_X1 U613 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U614 ( .A1(n567), .A2(n566), .ZN(n926) );
  XNOR2_X1 U615 ( .A(n926), .B(G2096), .ZN(n568) );
  XNOR2_X1 U616 ( .A(n568), .B(KEYINPUT77), .ZN(n569) );
  OR2_X1 U617 ( .A1(G2100), .A2(n569), .ZN(G156) );
  NAND2_X1 U618 ( .A1(n650), .A2(G53), .ZN(n571) );
  NAND2_X1 U619 ( .A1(G65), .A2(n651), .ZN(n570) );
  NAND2_X1 U620 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U621 ( .A1(n654), .A2(G78), .ZN(n573) );
  NAND2_X1 U622 ( .A1(G91), .A2(n655), .ZN(n572) );
  NAND2_X1 U623 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U624 ( .A1(n575), .A2(n574), .ZN(n695) );
  INV_X1 U625 ( .A(n695), .ZN(G299) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G120), .ZN(G236) );
  INV_X1 U628 ( .A(G132), .ZN(G219) );
  INV_X1 U629 ( .A(G82), .ZN(G220) );
  NAND2_X1 U630 ( .A1(n650), .A2(G52), .ZN(n577) );
  NAND2_X1 U631 ( .A1(G64), .A2(n651), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U633 ( .A1(n654), .A2(G77), .ZN(n579) );
  NAND2_X1 U634 ( .A1(G90), .A2(n655), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n580), .Z(n581) );
  NOR2_X1 U637 ( .A1(n582), .A2(n581), .ZN(G171) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n583) );
  XOR2_X1 U641 ( .A(n583), .B(KEYINPUT10), .Z(n925) );
  NAND2_X1 U642 ( .A1(n925), .A2(G567), .ZN(n584) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U644 ( .A1(n651), .A2(G56), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n585), .Z(n592) );
  NAND2_X1 U646 ( .A1(n655), .A2(G81), .ZN(n586) );
  XOR2_X1 U647 ( .A(KEYINPUT73), .B(n586), .Z(n587) );
  XNOR2_X1 U648 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U649 ( .A1(G68), .A2(n654), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U652 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U653 ( .A1(n650), .A2(G43), .ZN(n593) );
  NAND2_X1 U654 ( .A1(n594), .A2(n593), .ZN(n978) );
  INV_X1 U655 ( .A(G860), .ZN(n606) );
  OR2_X1 U656 ( .A1(n978), .A2(n606), .ZN(G153) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U658 ( .A1(G92), .A2(n655), .ZN(n596) );
  NAND2_X1 U659 ( .A1(G66), .A2(n651), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U661 ( .A1(G79), .A2(n654), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G54), .A2(n650), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U664 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U665 ( .A(KEYINPUT15), .B(n601), .ZN(n607) );
  INV_X1 U666 ( .A(G868), .ZN(n664) );
  NAND2_X1 U667 ( .A1(n607), .A2(n664), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U670 ( .A1(G286), .A2(n664), .ZN(n604) );
  NOR2_X1 U671 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n606), .A2(G559), .ZN(n608) );
  INV_X1 U673 ( .A(n607), .ZN(n973) );
  NAND2_X1 U674 ( .A1(n608), .A2(n973), .ZN(n609) );
  XNOR2_X1 U675 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n978), .ZN(n612) );
  NAND2_X1 U677 ( .A1(G868), .A2(n973), .ZN(n610) );
  NOR2_X1 U678 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U680 ( .A(KEYINPUT75), .B(n613), .Z(G282) );
  NAND2_X1 U681 ( .A1(n614), .A2(G87), .ZN(n615) );
  XNOR2_X1 U682 ( .A(n615), .B(KEYINPUT80), .ZN(n620) );
  NAND2_X1 U683 ( .A1(G49), .A2(n650), .ZN(n617) );
  NAND2_X1 U684 ( .A1(G74), .A2(G651), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U686 ( .A1(n651), .A2(n618), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(G288) );
  NAND2_X1 U688 ( .A1(n650), .A2(G47), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G60), .A2(n651), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U691 ( .A1(G85), .A2(n655), .ZN(n623) );
  XNOR2_X1 U692 ( .A(KEYINPUT69), .B(n623), .ZN(n624) );
  NOR2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n654), .A2(G72), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U696 ( .A1(G88), .A2(n655), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G62), .A2(n651), .ZN(n628) );
  NAND2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U699 ( .A1(G50), .A2(n650), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT82), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n654), .A2(G75), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U703 ( .A1(n634), .A2(n633), .ZN(G166) );
  INV_X1 U704 ( .A(G166), .ZN(G303) );
  NAND2_X1 U705 ( .A1(G73), .A2(n654), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n635), .Z(n640) );
  NAND2_X1 U707 ( .A1(G86), .A2(n655), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G61), .A2(n651), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U710 ( .A(KEYINPUT81), .B(n638), .Z(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n650), .A2(G48), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G559), .A2(n973), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(n978), .ZN(n833) );
  XNOR2_X1 U716 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n645) );
  XNOR2_X1 U717 ( .A(G290), .B(KEYINPUT83), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U719 ( .A(G288), .B(n646), .ZN(n648) );
  XOR2_X1 U720 ( .A(G303), .B(n695), .Z(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(G305), .ZN(n662) );
  NAND2_X1 U723 ( .A1(n650), .A2(G55), .ZN(n653) );
  NAND2_X1 U724 ( .A1(G67), .A2(n651), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n660) );
  NAND2_X1 U726 ( .A1(n654), .A2(G80), .ZN(n657) );
  NAND2_X1 U727 ( .A1(G93), .A2(n655), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT78), .B(n658), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT79), .ZN(n835) );
  XNOR2_X1 U732 ( .A(n662), .B(n835), .ZN(n892) );
  XNOR2_X1 U733 ( .A(n833), .B(n892), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n663), .A2(G868), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n664), .A2(n835), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U745 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U746 ( .A1(G96), .A2(n673), .ZN(n831) );
  NAND2_X1 U747 ( .A1(n831), .A2(G2106), .ZN(n679) );
  NOR2_X1 U748 ( .A1(G236), .A2(G237), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G69), .A2(n674), .ZN(n675) );
  XNOR2_X1 U750 ( .A(KEYINPUT85), .B(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G108), .ZN(n677) );
  XNOR2_X1 U752 ( .A(KEYINPUT86), .B(n677), .ZN(n832) );
  NAND2_X1 U753 ( .A1(n832), .A2(G567), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n679), .A2(n678), .ZN(n924) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U756 ( .A1(n924), .A2(n680), .ZN(n830) );
  NAND2_X1 U757 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(n681), .A2(G138), .ZN(n683) );
  NAND2_X1 U759 ( .A1(G126), .A2(n862), .ZN(n682) );
  NAND2_X1 U760 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U761 ( .A1(G102), .A2(n858), .ZN(n685) );
  NAND2_X1 U762 ( .A1(G114), .A2(n863), .ZN(n684) );
  NAND2_X1 U763 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U764 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U765 ( .A(KEYINPUT87), .B(n688), .Z(G164) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n776) );
  NAND2_X1 U767 ( .A1(G40), .A2(G160), .ZN(n689) );
  XOR2_X1 U768 ( .A(n689), .B(KEYINPUT88), .Z(n775) );
  NAND2_X2 U769 ( .A1(n776), .A2(n775), .ZN(n730) );
  INV_X1 U770 ( .A(n730), .ZN(n714) );
  NAND2_X1 U771 ( .A1(n714), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U772 ( .A(n690), .B(KEYINPUT27), .ZN(n692) );
  INV_X1 U773 ( .A(G1956), .ZN(n897) );
  NOR2_X1 U774 ( .A1(n897), .A2(n714), .ZN(n691) );
  NOR2_X1 U775 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U776 ( .A1(n696), .A2(n695), .ZN(n694) );
  XOR2_X1 U777 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n693) );
  XNOR2_X1 U778 ( .A(n694), .B(n693), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n710) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n730), .ZN(n698) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n714), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U783 ( .A(KEYINPUT97), .B(n699), .ZN(n706) );
  OR2_X1 U784 ( .A1(n973), .A2(n706), .ZN(n705) );
  AND2_X1 U785 ( .A1(n714), .A2(G1996), .ZN(n700) );
  XOR2_X1 U786 ( .A(n700), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U787 ( .A1(n730), .A2(G1341), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U789 ( .A1(n978), .A2(n703), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U791 ( .A1(n706), .A2(n973), .ZN(n707) );
  AND2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U793 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U794 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U795 ( .A(n713), .B(KEYINPUT29), .ZN(n718) );
  NAND2_X1 U796 ( .A1(G1961), .A2(n730), .ZN(n716) );
  XOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .Z(n957) );
  NAND2_X1 U798 ( .A1(n714), .A2(n957), .ZN(n715) );
  NAND2_X1 U799 ( .A1(n716), .A2(n715), .ZN(n725) );
  NOR2_X1 U800 ( .A1(G301), .A2(n725), .ZN(n717) );
  NOR2_X1 U801 ( .A1(n718), .A2(n717), .ZN(n729) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n769), .ZN(n742) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n730), .ZN(n743) );
  NOR2_X1 U804 ( .A1(n742), .A2(n743), .ZN(n719) );
  XNOR2_X1 U805 ( .A(n719), .B(KEYINPUT98), .ZN(n720) );
  NAND2_X1 U806 ( .A1(n720), .A2(G8), .ZN(n721) );
  XNOR2_X1 U807 ( .A(n721), .B(KEYINPUT30), .ZN(n722) );
  XNOR2_X1 U808 ( .A(n722), .B(KEYINPUT99), .ZN(n724) );
  AND2_X1 U809 ( .A1(G301), .A2(n725), .ZN(n726) );
  NOR2_X1 U810 ( .A1(n524), .A2(n726), .ZN(n727) );
  XNOR2_X1 U811 ( .A(n727), .B(KEYINPUT31), .ZN(n728) );
  NOR2_X1 U812 ( .A1(n729), .A2(n728), .ZN(n741) );
  OR2_X1 U813 ( .A1(n741), .A2(n525), .ZN(n739) );
  INV_X1 U814 ( .A(G8), .ZN(n737) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n769), .ZN(n732) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U817 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U818 ( .A(KEYINPUT101), .B(n733), .Z(n734) );
  NAND2_X1 U819 ( .A1(n734), .A2(G303), .ZN(n735) );
  XNOR2_X1 U820 ( .A(n735), .B(KEYINPUT102), .ZN(n736) );
  OR2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n738) );
  AND2_X1 U822 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U823 ( .A(n740), .B(KEYINPUT32), .ZN(n748) );
  NOR2_X1 U824 ( .A1(n742), .A2(n741), .ZN(n745) );
  NAND2_X1 U825 ( .A1(G8), .A2(n743), .ZN(n744) );
  NAND2_X1 U826 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U827 ( .A(n746), .B(KEYINPUT100), .ZN(n747) );
  NAND2_X1 U828 ( .A1(n748), .A2(n747), .ZN(n758) );
  NOR2_X1 U829 ( .A1(G2090), .A2(G303), .ZN(n749) );
  NAND2_X1 U830 ( .A1(G8), .A2(n749), .ZN(n750) );
  NAND2_X1 U831 ( .A1(n758), .A2(n750), .ZN(n751) );
  XNOR2_X1 U832 ( .A(n751), .B(KEYINPUT104), .ZN(n752) );
  AND2_X1 U833 ( .A1(n752), .A2(n769), .ZN(n773) );
  XOR2_X1 U834 ( .A(G1981), .B(G305), .Z(n990) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n760) );
  INV_X1 U836 ( .A(n760), .ZN(n977) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n753) );
  XNOR2_X1 U838 ( .A(n753), .B(KEYINPUT103), .ZN(n754) );
  AND2_X1 U839 ( .A1(n977), .A2(n754), .ZN(n756) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n755) );
  AND2_X1 U841 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n758), .A2(n757), .ZN(n765) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n976) );
  INV_X1 U844 ( .A(n976), .ZN(n759) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n526), .ZN(n763) );
  NAND2_X1 U846 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U847 ( .A1(n761), .A2(n769), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n764) );
  AND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U850 ( .A1(n990), .A2(n766), .ZN(n771) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U852 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  OR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U855 ( .A1(n773), .A2(n772), .ZN(n774) );
  INV_X1 U856 ( .A(n774), .ZN(n812) );
  INV_X1 U857 ( .A(n775), .ZN(n777) );
  NOR2_X1 U858 ( .A1(n777), .A2(n776), .ZN(n822) );
  XNOR2_X1 U859 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n782) );
  NAND2_X1 U860 ( .A1(G128), .A2(n862), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G116), .A2(n863), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U863 ( .A(n780), .B(KEYINPUT35), .ZN(n781) );
  XNOR2_X1 U864 ( .A(n782), .B(n781), .ZN(n788) );
  NAND2_X1 U865 ( .A1(n858), .A2(G104), .ZN(n783) );
  XOR2_X1 U866 ( .A(KEYINPUT89), .B(n783), .Z(n785) );
  NAND2_X1 U867 ( .A1(n859), .A2(G140), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U869 ( .A(KEYINPUT34), .B(n786), .ZN(n787) );
  NOR2_X1 U870 ( .A1(n788), .A2(n787), .ZN(n790) );
  XNOR2_X1 U871 ( .A(KEYINPUT92), .B(KEYINPUT36), .ZN(n789) );
  XNOR2_X1 U872 ( .A(n790), .B(n789), .ZN(n876) );
  XNOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NOR2_X1 U874 ( .A1(n876), .A2(n820), .ZN(n946) );
  NAND2_X1 U875 ( .A1(n822), .A2(n946), .ZN(n818) );
  NAND2_X1 U876 ( .A1(n859), .A2(G131), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G119), .A2(n862), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G95), .A2(n858), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G107), .A2(n863), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n854) );
  AND2_X1 U883 ( .A1(n854), .A2(G1991), .ZN(n808) );
  NAND2_X1 U884 ( .A1(G105), .A2(n858), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n797), .B(KEYINPUT38), .ZN(n806) );
  NAND2_X1 U886 ( .A1(n863), .A2(G117), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT94), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G141), .A2(n859), .ZN(n799) );
  XOR2_X1 U889 ( .A(KEYINPUT95), .B(n799), .Z(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G129), .A2(n862), .ZN(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT93), .B(n802), .ZN(n803) );
  NOR2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n870) );
  AND2_X1 U895 ( .A1(n870), .A2(G1996), .ZN(n807) );
  NOR2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n936) );
  INV_X1 U897 ( .A(n822), .ZN(n809) );
  NOR2_X1 U898 ( .A1(n936), .A2(n809), .ZN(n815) );
  INV_X1 U899 ( .A(n815), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n818), .A2(n810), .ZN(n811) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U902 ( .A1(n812), .A2(n527), .ZN(n825) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n870), .ZN(n931) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n854), .ZN(n927) );
  NOR2_X1 U906 ( .A1(n813), .A2(n927), .ZN(n814) );
  NOR2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U908 ( .A1(n931), .A2(n816), .ZN(n817) );
  XNOR2_X1 U909 ( .A(KEYINPUT39), .B(n817), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n876), .A2(n820), .ZN(n943) );
  NAND2_X1 U912 ( .A1(n821), .A2(n943), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U915 ( .A(KEYINPUT40), .B(n826), .ZN(G329) );
  NAND2_X1 U916 ( .A1(n925), .A2(G2106), .ZN(n827) );
  XNOR2_X1 U917 ( .A(n827), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  NOR2_X1 U927 ( .A1(G860), .A2(n833), .ZN(n834) );
  XOR2_X1 U928 ( .A(n835), .B(n834), .Z(G145) );
  NAND2_X1 U929 ( .A1(n862), .A2(G124), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT44), .ZN(n837) );
  XNOR2_X1 U931 ( .A(KEYINPUT110), .B(n837), .ZN(n840) );
  NAND2_X1 U932 ( .A1(G100), .A2(n858), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT111), .B(n838), .Z(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n844) );
  NAND2_X1 U935 ( .A1(G136), .A2(n859), .ZN(n842) );
  NAND2_X1 U936 ( .A1(G112), .A2(n863), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G162) );
  NAND2_X1 U939 ( .A1(G130), .A2(n862), .ZN(n846) );
  NAND2_X1 U940 ( .A1(G118), .A2(n863), .ZN(n845) );
  NAND2_X1 U941 ( .A1(n846), .A2(n845), .ZN(n851) );
  NAND2_X1 U942 ( .A1(G106), .A2(n858), .ZN(n848) );
  NAND2_X1 U943 ( .A1(G142), .A2(n859), .ZN(n847) );
  NAND2_X1 U944 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U945 ( .A(n849), .B(KEYINPUT45), .Z(n850) );
  NOR2_X1 U946 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U947 ( .A(KEYINPUT113), .B(n852), .Z(n853) );
  XOR2_X1 U948 ( .A(n853), .B(KEYINPUT48), .Z(n856) );
  XOR2_X1 U949 ( .A(n854), .B(KEYINPUT46), .Z(n855) );
  XNOR2_X1 U950 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U951 ( .A(n857), .B(G162), .Z(n872) );
  NAND2_X1 U952 ( .A1(G103), .A2(n858), .ZN(n861) );
  NAND2_X1 U953 ( .A1(G139), .A2(n859), .ZN(n860) );
  NAND2_X1 U954 ( .A1(n861), .A2(n860), .ZN(n868) );
  NAND2_X1 U955 ( .A1(G127), .A2(n862), .ZN(n865) );
  NAND2_X1 U956 ( .A1(G115), .A2(n863), .ZN(n864) );
  NAND2_X1 U957 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U958 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U959 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U960 ( .A(KEYINPUT112), .B(n869), .Z(n937) );
  XOR2_X1 U961 ( .A(n870), .B(n937), .Z(n871) );
  XNOR2_X1 U962 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U963 ( .A(n873), .B(n926), .Z(n875) );
  XNOR2_X1 U964 ( .A(G160), .B(G164), .ZN(n874) );
  XNOR2_X1 U965 ( .A(n875), .B(n874), .ZN(n877) );
  XNOR2_X1 U966 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U967 ( .A1(G37), .A2(n878), .ZN(n879) );
  XNOR2_X1 U968 ( .A(KEYINPUT114), .B(n879), .ZN(G395) );
  XNOR2_X1 U969 ( .A(G1348), .B(G2454), .ZN(n880) );
  XNOR2_X1 U970 ( .A(n880), .B(G2430), .ZN(n881) );
  XNOR2_X1 U971 ( .A(n881), .B(G1341), .ZN(n887) );
  XOR2_X1 U972 ( .A(G2443), .B(G2427), .Z(n883) );
  XNOR2_X1 U973 ( .A(G2438), .B(G2446), .ZN(n882) );
  XNOR2_X1 U974 ( .A(n883), .B(n882), .ZN(n885) );
  XOR2_X1 U975 ( .A(G2451), .B(G2435), .Z(n884) );
  XNOR2_X1 U976 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U977 ( .A(n887), .B(n886), .ZN(n888) );
  NAND2_X1 U978 ( .A1(n888), .A2(G14), .ZN(n889) );
  XNOR2_X1 U979 ( .A(KEYINPUT105), .B(n889), .ZN(G401) );
  XNOR2_X1 U980 ( .A(n978), .B(KEYINPUT115), .ZN(n891) );
  XOR2_X1 U981 ( .A(G301), .B(n973), .Z(n890) );
  XNOR2_X1 U982 ( .A(n891), .B(n890), .ZN(n894) );
  XNOR2_X1 U983 ( .A(G286), .B(n892), .ZN(n893) );
  XNOR2_X1 U984 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U985 ( .A1(G37), .A2(n895), .ZN(n896) );
  XNOR2_X1 U986 ( .A(KEYINPUT116), .B(n896), .ZN(G397) );
  XOR2_X1 U987 ( .A(G1976), .B(G1981), .Z(n899) );
  XOR2_X1 U988 ( .A(G1991), .B(n897), .Z(n898) );
  XNOR2_X1 U989 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U990 ( .A(G1971), .B(G1966), .Z(n901) );
  XNOR2_X1 U991 ( .A(G1986), .B(G1961), .ZN(n900) );
  XNOR2_X1 U992 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U993 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U994 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n904) );
  XNOR2_X1 U995 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U996 ( .A(G2474), .B(n906), .ZN(n907) );
  XOR2_X1 U997 ( .A(n907), .B(G1996), .Z(G229) );
  XOR2_X1 U998 ( .A(KEYINPUT108), .B(G2678), .Z(n909) );
  XNOR2_X1 U999 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1001 ( .A(KEYINPUT42), .B(G2072), .Z(n911) );
  XNOR2_X1 U1002 ( .A(G2067), .B(G2090), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1004 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1005 ( .A(G2096), .B(G2100), .ZN(n914) );
  XNOR2_X1 U1006 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1007 ( .A(G2078), .B(G2084), .Z(n916) );
  XNOR2_X1 U1008 ( .A(n917), .B(n916), .ZN(G227) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n924), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(KEYINPUT117), .B(n918), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G395), .A2(n919), .ZN(n923) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n921), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n924), .ZN(G319) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  INV_X1 U1019 ( .A(n925), .ZN(G223) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n929) );
  NOR2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1022 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(n932), .B(KEYINPUT51), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n939) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n937), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1032 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1033 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1034 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1035 ( .A(KEYINPUT52), .B(n947), .Z(n948) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n948), .ZN(n949) );
  XOR2_X1 U1037 ( .A(KEYINPUT118), .B(n949), .Z(n950) );
  NAND2_X1 U1038 ( .A1(n950), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1039 ( .A(G2072), .B(G33), .Z(n951) );
  NAND2_X1 U1040 ( .A1(n951), .A2(G28), .ZN(n954) );
  XOR2_X1 U1041 ( .A(G25), .B(G1991), .Z(n952) );
  XNOR2_X1 U1042 ( .A(KEYINPUT119), .B(n952), .ZN(n953) );
  NOR2_X1 U1043 ( .A1(n954), .A2(n953), .ZN(n961) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n956) );
  XOR2_X1 U1045 ( .A(G1996), .B(G32), .Z(n955) );
  NAND2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1047 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1048 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1049 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1050 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1051 ( .A(G2084), .B(KEYINPUT54), .Z(n963) );
  XNOR2_X1 U1052 ( .A(G34), .B(n963), .ZN(n964) );
  NAND2_X1 U1053 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1055 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n968), .ZN(n970) );
  INV_X1 U1057 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1058 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1059 ( .A1(n971), .A2(G11), .ZN(n1027) );
  XOR2_X1 U1060 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n972) );
  XOR2_X1 U1061 ( .A(G16), .B(n972), .Z(n997) );
  XOR2_X1 U1062 ( .A(G171), .B(G1961), .Z(n975) );
  XOR2_X1 U1063 ( .A(n973), .B(G1348), .Z(n974) );
  NOR2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n986) );
  XOR2_X1 U1065 ( .A(G299), .B(G1956), .Z(n982) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1071 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1072 ( .A(G1971), .B(G166), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NOR2_X1 U1074 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1075 ( .A(G168), .B(G1966), .ZN(n991) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(n992), .B(KEYINPUT57), .ZN(n993) );
  NAND2_X1 U1078 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(n995), .B(KEYINPUT122), .ZN(n996) );
  NAND2_X1 U1080 ( .A1(n997), .A2(n996), .ZN(n1025) );
  INV_X1 U1081 ( .A(G16), .ZN(n1023) );
  XOR2_X1 U1082 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n1021) );
  XNOR2_X1 U1083 ( .A(G1961), .B(G5), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G21), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1019) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n1006) );
  XNOR2_X1 U1087 ( .A(G1986), .B(G24), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1090 ( .A(G1971), .B(KEYINPUT124), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(G22), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(n1006), .B(n1005), .ZN(n1017) );
  XOR2_X1 U1094 ( .A(G20), .B(G1956), .Z(n1010) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT59), .B(G1348), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT123), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT60), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1110 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(n1030), .B(KEYINPUT62), .ZN(n1031) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1031), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

