//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT0), .A3(G128), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G134), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G137), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n200), .A2(new_n202), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n198), .A4(new_n199), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n198), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n191), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n188), .A2(new_n212), .A3(G128), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n212), .A2(new_n217), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n199), .B1(G134), .B2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n193), .A2(new_n195), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT66), .B(new_n224), .C1(new_n225), .C2(G137), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n208), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n223), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n205), .A2(new_n207), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n211), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n236), .B2(KEYINPUT30), .ZN(new_n237));
  XNOR2_X1  g051(.A(G116), .B(G119), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n240), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(KEYINPUT70), .A3(new_n240), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n208), .A2(new_n210), .ZN(new_n248));
  INV_X1    g062(.A(new_n191), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n221), .A2(new_n222), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n234), .B2(KEYINPUT67), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n208), .A2(KEYINPUT67), .A3(new_n230), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n211), .B1(new_n251), .B2(new_n234), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT30), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n237), .A2(new_n247), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n250), .B(new_n246), .C1(new_n223), .C2(new_n231), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n261), .A2(KEYINPUT71), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT71), .B1(new_n261), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n260), .A2(KEYINPUT72), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n260), .A2(new_n270), .A3(KEYINPUT72), .A4(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n267), .B(KEYINPUT73), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n254), .A2(new_n278), .A3(new_n247), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n236), .A2(new_n246), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n261), .A2(KEYINPUT74), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT28), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n261), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT28), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n277), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n286), .B1(new_n273), .B2(new_n274), .ZN(new_n292));
  INV_X1    g106(.A(new_n290), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT32), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G472), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n260), .A2(new_n261), .ZN(new_n297));
  INV_X1    g111(.A(new_n267), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n282), .A2(new_n285), .A3(new_n277), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n258), .B(new_n246), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n284), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n298), .A2(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n296), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n187), .B1(new_n295), .B2(new_n308), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT75), .B(new_n307), .C1(new_n291), .C2(new_n294), .ZN(new_n310));
  INV_X1    g124(.A(G217), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(G234), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n219), .A2(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(KEYINPUT77), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(KEYINPUT77), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT23), .A3(new_n315), .ZN(new_n320));
  INV_X1    g134(.A(G110), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT24), .B(G110), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n315), .A2(new_n317), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT76), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT78), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n326), .A2(new_n327), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n330), .B(new_n331), .C1(new_n332), .C2(new_n323), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT16), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n343), .A2(KEYINPUT79), .A3(G146), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n343), .B2(G146), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n340), .A2(G146), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(new_n333), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n332), .A2(new_n323), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n318), .A2(new_n320), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G110), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n340), .A2(G146), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n339), .A2(new_n214), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n348), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n347), .A2(new_n353), .A3(KEYINPUT80), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT25), .B1(new_n364), .B2(new_n312), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  AOI211_X1 g180(.A(new_n366), .B(G902), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n313), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT81), .B(new_n313), .C1(new_n365), .C2(new_n367), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n313), .A2(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n309), .A2(new_n310), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n208), .A2(new_n210), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G107), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n377), .A2(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n251), .A2(KEYINPUT10), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n213), .A2(new_n220), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n216), .A2(KEYINPUT1), .A3(G146), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(G101), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n249), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n376), .A2(new_n390), .A3(new_n395), .A4(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G140), .ZN(new_n403));
  INV_X1    g217(.A(G227), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G953), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n402), .A2(KEYINPUT84), .A3(new_n407), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n390), .A2(new_n395), .A3(new_n401), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n248), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n221), .A2(new_n222), .A3(new_n388), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n393), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT12), .A3(new_n248), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n416), .A2(KEYINPUT83), .A3(new_n248), .A4(KEYINPUT12), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n248), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n407), .B1(new_n424), .B2(new_n402), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT85), .B1(new_n414), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n424), .A2(new_n402), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n427), .B(new_n428), .C1(new_n429), .C2(new_n407), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n430), .A3(new_n312), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G469), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n434), .A3(G469), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n408), .B1(new_n424), .B2(KEYINPUT87), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n419), .A2(new_n423), .A3(new_n437), .A4(new_n420), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n413), .A2(new_n402), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n406), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n312), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n433), .A2(new_n435), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT9), .B(G234), .ZN(new_n446));
  OAI21_X1  g260(.A(G221), .B1(new_n446), .B2(G902), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT82), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n398), .A2(new_n400), .A3(new_n245), .A4(new_n244), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n314), .A3(G116), .ZN(new_n452));
  OAI211_X1 g266(.A(G113), .B(new_n452), .C1(new_n239), .C2(new_n451), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n389), .A2(new_n241), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n241), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n388), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n454), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(KEYINPUT88), .A3(new_n388), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n455), .B(KEYINPUT8), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n251), .A2(new_n341), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n249), .A2(G125), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n263), .A2(G224), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT7), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n466), .B2(new_n467), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n456), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n472), .A2(new_n312), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n450), .A2(new_n454), .ZN(new_n474));
  INV_X1    g288(.A(new_n455), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n466), .B(new_n468), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT90), .Z(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n473), .A2(new_n483), .A3(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G475), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(G143), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT91), .ZN(new_n493));
  AND2_X1   g307(.A1(KEYINPUT18), .A2(G131), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n344), .A2(new_n345), .B1(G146), .B2(new_n343), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n377), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n351), .A2(new_n352), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n492), .A2(new_n199), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT17), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n492), .B(new_n199), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(new_n502), .C1(KEYINPUT17), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n497), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n334), .B(KEYINPUT19), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n352), .B1(new_n214), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n503), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n499), .B1(new_n497), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n490), .B(new_n312), .C1(new_n506), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT20), .ZN(new_n512));
  INV_X1    g326(.A(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n505), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT20), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n490), .A4(new_n312), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n499), .B1(new_n497), .B2(new_n504), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n312), .B1(new_n506), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n512), .A2(new_n516), .B1(G475), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n263), .A2(G952), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT94), .Z(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT21), .B(G898), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n527), .B(KEYINPUT95), .Z(new_n528));
  XNOR2_X1  g342(.A(G116), .B(G122), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G122), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(G116), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n380), .B1(new_n533), .B2(KEYINPUT14), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n531), .A2(new_n534), .B1(new_n380), .B2(new_n529), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT92), .B1(new_n219), .B2(G143), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n216), .A3(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT64), .B(G134), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n219), .A2(G143), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT93), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n535), .B(new_n546), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n529), .A2(new_n380), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n529), .A2(new_n380), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n539), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT13), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n553), .A2(new_n541), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n555), .B2(new_n192), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n446), .A2(new_n311), .A3(G953), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n548), .A2(new_n556), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n312), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n519), .A2(new_n528), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n489), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n445), .A2(new_n449), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT96), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n375), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  NAND2_X1  g389(.A1(new_n288), .A2(new_n312), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT97), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n288), .A2(new_n290), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n580), .A3(G472), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n445), .A2(new_n449), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n582), .A2(new_n374), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n562), .A2(new_n564), .A3(new_n312), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n548), .A2(new_n556), .A3(new_n558), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n558), .B1(new_n548), .B2(new_n556), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT33), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n560), .A2(new_n589), .A3(new_n561), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n585), .B1(new_n591), .B2(new_n564), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT98), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n585), .C1(new_n591), .C2(new_n564), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n512), .A2(new_n516), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n518), .A2(G475), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n488), .ZN(new_n601));
  INV_X1    g415(.A(new_n483), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n482), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n603), .B2(new_n486), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n528), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n584), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT99), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT34), .B(G104), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  NOR2_X1   g425(.A1(new_n599), .A2(new_n569), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n528), .B(KEYINPUT100), .Z(new_n613));
  AND3_X1   g427(.A1(new_n612), .A2(new_n604), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n584), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n354), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n372), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n370), .A2(new_n371), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n370), .A2(KEYINPUT102), .A3(new_n371), .A4(new_n621), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT103), .B1(new_n582), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n581), .A2(new_n579), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n630));
  INV_X1    g444(.A(new_n626), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n578), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n627), .A2(new_n573), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G12));
  AOI21_X1  g450(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n293), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n308), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT75), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n295), .A2(new_n187), .A3(new_n308), .ZN(new_n641));
  INV_X1    g455(.A(new_n583), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n523), .B1(G900), .B2(new_n526), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n599), .A2(new_n569), .A3(new_n644), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n604), .A2(new_n624), .A3(new_n625), .A4(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n640), .A2(new_n641), .A3(new_n642), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  XNOR2_X1  g462(.A(new_n643), .B(KEYINPUT39), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n445), .A2(new_n449), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n260), .A2(new_n270), .B1(new_n276), .B2(new_n303), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n653), .B2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n295), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n487), .B(KEYINPUT38), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n599), .A2(new_n568), .A3(new_n488), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n622), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n652), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G143), .ZN(G45));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n600), .B2(new_n644), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n519), .B1(new_n593), .B2(new_n595), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT105), .A3(new_n643), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n624), .A2(new_n604), .A3(new_n625), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n436), .A2(new_n438), .B1(new_n406), .B2(new_n440), .ZN(new_n672));
  OAI21_X1  g486(.A(G469), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n444), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n674), .B2(new_n448), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n444), .A2(new_n673), .A3(KEYINPUT106), .A4(new_n449), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n375), .A2(new_n607), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT107), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(G15));
  NOR2_X1   g495(.A1(new_n309), .A2(new_n310), .ZN(new_n682));
  INV_X1    g496(.A(new_n374), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n615), .A4(new_n677), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  INV_X1    g499(.A(new_n570), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n675), .A2(new_n686), .A3(new_n676), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n667), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n640), .A2(new_n688), .A3(new_n641), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NOR3_X1   g504(.A1(new_n605), .A2(new_n569), .A3(new_n519), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n677), .A2(new_n613), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT108), .B(G472), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n576), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n275), .B1(new_n277), .B2(new_n304), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n290), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n683), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n532), .ZN(G24));
  AND2_X1   g513(.A1(new_n694), .A2(new_n696), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n663), .A2(new_n665), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n675), .A2(new_n604), .A3(new_n676), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n622), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  NAND3_X1  g518(.A1(new_n485), .A2(new_n488), .A3(new_n486), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n443), .A2(new_n312), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n444), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n425), .A2(new_n709), .ZN(new_n710));
  AOI211_X1 g524(.A(KEYINPUT109), .B(new_n407), .C1(new_n424), .C2(new_n402), .ZN(new_n711));
  OAI211_X1 g525(.A(G469), .B(new_n428), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n448), .B(new_n705), .C1(new_n708), .C2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n701), .A2(new_n639), .A3(new_n683), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n640), .A2(new_n641), .A3(new_n683), .A4(new_n713), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT110), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n715), .B(new_n720), .C1(new_n716), .C2(new_n717), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  NAND3_X1  g537(.A1(new_n375), .A2(new_n645), .A3(new_n713), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n580), .B1(new_n576), .B2(G472), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n628), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n596), .A2(new_n519), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n622), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n726), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n705), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n582), .A2(KEYINPUT44), .A3(new_n622), .A4(new_n731), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT113), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n733), .A2(new_n735), .A3(new_n738), .A4(new_n734), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n426), .A2(new_n430), .A3(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(KEYINPUT45), .B(new_n428), .C1(new_n710), .C2(new_n711), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(G469), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n707), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n444), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(KEYINPUT111), .A3(new_n444), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  INV_X1    g563(.A(new_n743), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(new_n706), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n449), .A3(new_n649), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(KEYINPUT112), .A3(new_n449), .A4(new_n649), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n737), .A2(new_n739), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  NAND3_X1  g573(.A1(new_n701), .A2(new_n374), .A3(new_n734), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n682), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n449), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT47), .B1(new_n752), .B2(new_n449), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n761), .B(KEYINPUT114), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  INV_X1    g584(.A(new_n489), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n664), .A3(new_n613), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT117), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT117), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n612), .A3(new_n613), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n584), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n633), .A2(new_n777), .A3(new_n574), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n692), .A2(new_n697), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n640), .A2(new_n641), .A3(new_n683), .A4(new_n677), .ZN(new_n780));
  INV_X1    g594(.A(new_n607), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n689), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n615), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT116), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n698), .B1(new_n682), .B2(new_n688), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n678), .A2(new_n786), .A3(new_n684), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n778), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n705), .A2(new_n599), .A3(new_n568), .A4(new_n644), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n682), .A2(new_n642), .A3(new_n631), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n700), .A2(new_n701), .A3(new_n622), .A4(new_n713), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n647), .A2(new_n703), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n691), .A2(new_n643), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n622), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n448), .B1(new_n708), .B2(new_n712), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n655), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(KEYINPUT52), .A3(new_n669), .A4(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n669), .A2(new_n647), .A3(new_n798), .A4(new_n703), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n793), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n789), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n789), .A2(new_n803), .A3(new_n804), .A4(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(KEYINPUT118), .A3(new_n806), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n523), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n731), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n677), .A2(new_n734), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n374), .B1(new_n295), .B2(new_n308), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT48), .Z(new_n819));
  NOR2_X1   g633(.A1(new_n814), .A2(new_n697), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n702), .ZN(new_n821));
  OR4_X1    g635(.A1(new_n374), .A2(new_n655), .A3(new_n815), .A4(new_n523), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n520), .B(new_n821), .C1(new_n822), .C2(new_n600), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n622), .A3(new_n700), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT120), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n822), .A2(new_n599), .A3(new_n596), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n763), .A2(new_n764), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n674), .A2(new_n449), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n734), .B(new_n820), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n601), .A2(new_n820), .A3(new_n657), .A4(new_n677), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT119), .B(KEYINPUT50), .Z(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(KEYINPUT119), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n828), .A2(new_n831), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n824), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n678), .A2(new_n786), .A3(new_n684), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n724), .A2(KEYINPUT53), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n778), .A2(new_n841), .A3(new_n842), .A4(new_n718), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n805), .A2(new_n806), .B1(new_n843), .B2(new_n803), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n812), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(G952), .B2(G953), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n374), .A2(new_n448), .A3(new_n601), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT115), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n674), .A2(KEYINPUT49), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n674), .A2(KEYINPUT49), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n656), .A2(new_n851), .A3(new_n852), .A4(new_n729), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n848), .B1(new_n655), .B2(new_n854), .ZN(G75));
  NOR2_X1   g669(.A1(new_n263), .A2(G952), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n844), .A2(new_n312), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n484), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n477), .A2(new_n479), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(new_n480), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT56), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n857), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n858), .A2(G210), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n866), .B2(new_n863), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n867), .ZN(G51));
  XNOR2_X1  g682(.A(new_n706), .B(KEYINPUT121), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT57), .Z(new_n870));
  NAND2_X1  g684(.A1(new_n843), .A2(new_n803), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n807), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n844), .A2(new_n845), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n442), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n858), .A2(new_n750), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n856), .B1(new_n876), .B2(new_n877), .ZN(G54));
  AND2_X1   g692(.A1(KEYINPUT58), .A2(G475), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n858), .A2(new_n514), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n514), .B1(new_n858), .B2(new_n879), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n856), .ZN(G60));
  AND2_X1   g696(.A1(new_n588), .A2(new_n590), .ZN(new_n883));
  NAND2_X1  g697(.A1(G478), .A2(G902), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT59), .Z(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n873), .B2(new_n874), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n857), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n812), .A2(new_n846), .ZN(new_n889));
  INV_X1    g703(.A(new_n885), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n888), .B1(new_n883), .B2(new_n891), .ZN(G63));
  NAND2_X1  g706(.A1(G217), .A2(G902), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT60), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n872), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n364), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n856), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n894), .B1(new_n807), .B2(new_n871), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n620), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(KEYINPUT122), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n857), .B1(new_n900), .B2(new_n364), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n872), .A2(new_n620), .A3(new_n895), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n902), .A2(new_n907), .ZN(G66));
  INV_X1    g722(.A(G224), .ZN(new_n909));
  OAI21_X1  g723(.A(G953), .B1(new_n524), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n789), .B2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n860), .B1(G898), .B2(new_n263), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G69));
  NAND3_X1  g727(.A1(new_n237), .A2(new_n257), .A3(new_n259), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(new_n507), .Z(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n794), .A2(new_n669), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n817), .A2(new_n691), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n755), .B2(new_n756), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n769), .A2(new_n758), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n917), .B1(new_n922), .B2(new_n804), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n769), .A2(new_n758), .A3(new_n921), .ZN(new_n924));
  INV_X1    g738(.A(new_n804), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT126), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n263), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n664), .A2(new_n612), .A3(KEYINPUT124), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT124), .B1(new_n664), .B2(new_n612), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n734), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n650), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n375), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n769), .A2(new_n758), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n660), .A2(new_n647), .A3(new_n669), .A4(new_n703), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT62), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n263), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(G900), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n936), .A2(KEYINPUT123), .B1(new_n937), .B2(G953), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n916), .B1(new_n927), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n404), .B2(new_n937), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n936), .A2(new_n942), .A3(new_n916), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n939), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n941), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n937), .A2(G953), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n922), .A2(new_n917), .A3(new_n804), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT126), .B1(new_n924), .B2(new_n925), .ZN(new_n951));
  AOI21_X1  g765(.A(G953), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n915), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n946), .B1(new_n953), .B2(new_n943), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n945), .A2(new_n954), .ZN(G72));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n789), .A3(new_n951), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n296), .A2(new_n312), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n267), .B(new_n297), .C1(new_n956), .C2(new_n960), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n933), .A2(new_n935), .ZN(new_n962));
  INV_X1    g776(.A(new_n789), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n964), .A2(new_n267), .A3(new_n297), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n260), .A2(new_n270), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n959), .B1(new_n299), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n810), .A2(new_n811), .A3(new_n967), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n961), .A2(new_n965), .A3(new_n968), .A4(new_n856), .ZN(G57));
endmodule


