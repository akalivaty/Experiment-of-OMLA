

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X2 U554 ( .A1(n654), .A2(n653), .ZN(n655) );
  BUF_X1 U555 ( .A(n604), .Z(n605) );
  NOR2_X2 U556 ( .A1(G2105), .A2(n528), .ZN(n600) );
  XOR2_X1 U557 ( .A(KEYINPUT100), .B(n726), .Z(n521) );
  INV_X1 U558 ( .A(KEYINPUT98), .ZN(n703) );
  XNOR2_X1 U559 ( .A(n704), .B(n703), .ZN(n716) );
  NOR2_X1 U560 ( .A1(n556), .A2(G651), .ZN(n793) );
  INV_X1 U561 ( .A(KEYINPUT104), .ZN(n762) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n791) );
  XNOR2_X1 U563 ( .A(n762), .B(KEYINPUT40), .ZN(n763) );
  XNOR2_X1 U564 ( .A(n764), .B(n763), .ZN(G329) );
  XNOR2_X1 U565 ( .A(n533), .B(KEYINPUT85), .ZN(G164) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U568 ( .A(n523), .B(n522), .ZN(n604) );
  NAND2_X1 U569 ( .A1(n604), .A2(G138), .ZN(n524) );
  XNOR2_X1 U570 ( .A(n524), .B(KEYINPUT84), .ZN(n526) );
  XOR2_X1 U571 ( .A(G2104), .B(KEYINPUT64), .Z(n528) );
  NAND2_X1 U572 ( .A1(n600), .A2(G102), .ZN(n525) );
  AND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n532) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U575 ( .A1(G114), .A2(n885), .ZN(n527) );
  XNOR2_X1 U576 ( .A(KEYINPUT83), .B(n527), .ZN(n530) );
  AND2_X1 U577 ( .A1(G2105), .A2(n528), .ZN(n884) );
  AND2_X1 U578 ( .A1(G126), .A2(n884), .ZN(n529) );
  NOR2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G113), .A2(n885), .ZN(n535) );
  NAND2_X1 U582 ( .A1(G137), .A2(n604), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U584 ( .A(KEYINPUT66), .B(n536), .ZN(n538) );
  AND2_X1 U585 ( .A1(n884), .A2(G125), .ZN(n537) );
  NOR2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n541) );
  NAND2_X1 U587 ( .A1(G101), .A2(n600), .ZN(n539) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  AND2_X1 U589 ( .A1(n541), .A2(n540), .ZN(G160) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n556) );
  NAND2_X1 U591 ( .A1(G47), .A2(n793), .ZN(n542) );
  XNOR2_X1 U592 ( .A(n542), .B(KEYINPUT68), .ZN(n551) );
  NAND2_X1 U593 ( .A1(G85), .A2(n791), .ZN(n545) );
  INV_X1 U594 ( .A(G651), .ZN(n546) );
  NOR2_X1 U595 ( .A1(G543), .A2(n546), .ZN(n543) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n543), .Z(n669) );
  NAND2_X1 U597 ( .A1(G60), .A2(n669), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n549) );
  NOR2_X1 U599 ( .A1(n556), .A2(n546), .ZN(n796) );
  NAND2_X1 U600 ( .A1(G72), .A2(n796), .ZN(n547) );
  XNOR2_X1 U601 ( .A(KEYINPUT67), .B(n547), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U604 ( .A(KEYINPUT69), .B(n552), .Z(G290) );
  NAND2_X1 U605 ( .A1(G49), .A2(n793), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G74), .A2(G651), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U608 ( .A1(n669), .A2(n555), .ZN(n558) );
  NAND2_X1 U609 ( .A1(n556), .A2(G87), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n558), .A2(n557), .ZN(G288) );
  NAND2_X1 U611 ( .A1(G65), .A2(n669), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G53), .A2(n793), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U614 ( .A1(G78), .A2(n796), .ZN(n562) );
  NAND2_X1 U615 ( .A1(G91), .A2(n791), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n563) );
  OR2_X1 U617 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G52), .A2(n793), .ZN(n565) );
  XOR2_X1 U619 ( .A(KEYINPUT70), .B(n565), .Z(n572) );
  NAND2_X1 U620 ( .A1(G77), .A2(n796), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G90), .A2(n791), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U623 ( .A(n568), .B(KEYINPUT9), .ZN(n570) );
  NAND2_X1 U624 ( .A1(G64), .A2(n669), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U626 ( .A1(n572), .A2(n571), .ZN(G171) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(n791), .A2(G89), .ZN(n573) );
  XNOR2_X1 U629 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U630 ( .A1(G76), .A2(n796), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U632 ( .A(n576), .B(KEYINPUT5), .ZN(n582) );
  NAND2_X1 U633 ( .A1(n669), .A2(G63), .ZN(n577) );
  XNOR2_X1 U634 ( .A(n577), .B(KEYINPUT76), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G51), .A2(n793), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U637 ( .A(KEYINPUT6), .B(n580), .Z(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U639 ( .A(n583), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U641 ( .A1(G75), .A2(n796), .ZN(n585) );
  NAND2_X1 U642 ( .A1(G88), .A2(n791), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U644 ( .A1(G62), .A2(n669), .ZN(n587) );
  NAND2_X1 U645 ( .A1(G50), .A2(n793), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U647 ( .A1(n589), .A2(n588), .ZN(G166) );
  XOR2_X1 U648 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U649 ( .A1(G61), .A2(n669), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G48), .A2(n793), .ZN(n590) );
  NAND2_X1 U651 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U652 ( .A1(G73), .A2(n796), .ZN(n592) );
  XOR2_X1 U653 ( .A(KEYINPUT2), .B(n592), .Z(n593) );
  NOR2_X1 U654 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U655 ( .A1(n791), .A2(G86), .ZN(n595) );
  NAND2_X1 U656 ( .A1(n596), .A2(n595), .ZN(G305) );
  NOR2_X1 U657 ( .A1(G164), .A2(G1384), .ZN(n658) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n640) );
  NOR2_X1 U659 ( .A1(n658), .A2(n640), .ZN(n752) );
  NAND2_X1 U660 ( .A1(G129), .A2(n884), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G117), .A2(n885), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(KEYINPUT92), .B(n599), .ZN(n603) );
  NAND2_X1 U664 ( .A1(G105), .A2(n600), .ZN(n601) );
  XOR2_X1 U665 ( .A(KEYINPUT38), .B(n601), .Z(n602) );
  NOR2_X1 U666 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U667 ( .A1(n605), .A2(G141), .ZN(n606) );
  NAND2_X1 U668 ( .A1(n607), .A2(n606), .ZN(n881) );
  NOR2_X1 U669 ( .A1(G1996), .A2(n881), .ZN(n983) );
  NAND2_X1 U670 ( .A1(n884), .A2(G119), .ZN(n608) );
  XOR2_X1 U671 ( .A(KEYINPUT89), .B(n608), .Z(n610) );
  NAND2_X1 U672 ( .A1(n885), .A2(G107), .ZN(n609) );
  NAND2_X1 U673 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U674 ( .A(KEYINPUT90), .B(n611), .Z(n615) );
  NAND2_X1 U675 ( .A1(n600), .A2(G95), .ZN(n613) );
  NAND2_X1 U676 ( .A1(G131), .A2(n605), .ZN(n612) );
  AND2_X1 U677 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U678 ( .A1(n615), .A2(n614), .ZN(n877) );
  NAND2_X1 U679 ( .A1(G1991), .A2(n877), .ZN(n616) );
  XNOR2_X1 U680 ( .A(n616), .B(KEYINPUT91), .ZN(n618) );
  AND2_X1 U681 ( .A1(G1996), .A2(n881), .ZN(n617) );
  NOR2_X1 U682 ( .A1(n618), .A2(n617), .ZN(n993) );
  XNOR2_X1 U683 ( .A(KEYINPUT93), .B(n752), .ZN(n619) );
  NOR2_X1 U684 ( .A1(n993), .A2(n619), .ZN(n753) );
  NOR2_X1 U685 ( .A1(G1986), .A2(G290), .ZN(n620) );
  NOR2_X1 U686 ( .A1(G1991), .A2(n877), .ZN(n987) );
  NOR2_X1 U687 ( .A1(n620), .A2(n987), .ZN(n621) );
  NOR2_X1 U688 ( .A1(n753), .A2(n621), .ZN(n622) );
  NOR2_X1 U689 ( .A1(n983), .A2(n622), .ZN(n623) );
  XNOR2_X1 U690 ( .A(n623), .B(KEYINPUT39), .ZN(n635) );
  NAND2_X1 U691 ( .A1(G104), .A2(n600), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G140), .A2(n605), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U694 ( .A(KEYINPUT34), .B(n626), .ZN(n632) );
  NAND2_X1 U695 ( .A1(G128), .A2(n884), .ZN(n628) );
  NAND2_X1 U696 ( .A1(G116), .A2(n885), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U698 ( .A(KEYINPUT35), .B(n629), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT87), .B(n630), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U701 ( .A(n633), .B(KEYINPUT36), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(KEYINPUT88), .ZN(n876) );
  XNOR2_X1 U703 ( .A(G2067), .B(KEYINPUT37), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n876), .A2(n636), .ZN(n979) );
  NAND2_X1 U705 ( .A1(n752), .A2(n979), .ZN(n754) );
  NAND2_X1 U706 ( .A1(n635), .A2(n754), .ZN(n637) );
  NAND2_X1 U707 ( .A1(n876), .A2(n636), .ZN(n988) );
  NAND2_X1 U708 ( .A1(n637), .A2(n988), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n752), .A2(n638), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n639), .B(KEYINPUT103), .ZN(n761) );
  NAND2_X1 U711 ( .A1(G1976), .A2(G288), .ZN(n923) );
  INV_X1 U712 ( .A(KEYINPUT28), .ZN(n646) );
  INV_X1 U713 ( .A(n640), .ZN(n656) );
  NAND2_X1 U714 ( .A1(n658), .A2(n656), .ZN(n705) );
  NAND2_X1 U715 ( .A1(G1956), .A2(n705), .ZN(n641) );
  XNOR2_X1 U716 ( .A(KEYINPUT96), .B(n641), .ZN(n644) );
  AND2_X1 U717 ( .A1(n658), .A2(n656), .ZN(n689) );
  NAND2_X1 U718 ( .A1(n689), .A2(G2072), .ZN(n642) );
  XOR2_X1 U719 ( .A(KEYINPUT27), .B(n642), .Z(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G299), .A2(n647), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(n686) );
  NOR2_X1 U723 ( .A1(G299), .A2(n647), .ZN(n684) );
  NAND2_X1 U724 ( .A1(G92), .A2(n791), .ZN(n649) );
  NAND2_X1 U725 ( .A1(G66), .A2(n669), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U727 ( .A(KEYINPUT74), .B(n650), .ZN(n654) );
  NAND2_X1 U728 ( .A1(G79), .A2(n796), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G54), .A2(n793), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U731 ( .A(KEYINPUT15), .B(n655), .Z(n920) );
  NAND2_X1 U732 ( .A1(n705), .A2(G1348), .ZN(n660) );
  AND2_X1 U733 ( .A1(G2067), .A2(n656), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(KEYINPUT97), .ZN(n680) );
  OR2_X1 U737 ( .A1(n920), .A2(n680), .ZN(n679) );
  AND2_X1 U738 ( .A1(n689), .A2(G1996), .ZN(n662) );
  XOR2_X1 U739 ( .A(n662), .B(KEYINPUT26), .Z(n677) );
  AND2_X1 U740 ( .A1(n705), .A2(G1341), .ZN(n675) );
  XNOR2_X1 U741 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n791), .A2(G81), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n663), .B(KEYINPUT12), .ZN(n665) );
  NAND2_X1 U744 ( .A1(G68), .A2(n796), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n666), .B(KEYINPUT13), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n669), .A2(G56), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT14), .B(n670), .Z(n671) );
  NOR2_X1 U750 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n793), .A2(G43), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n925) );
  NOR2_X1 U753 ( .A1(n675), .A2(n925), .ZN(n676) );
  AND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U756 ( .A1(n680), .A2(n920), .ZN(n681) );
  NAND2_X1 U757 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U758 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U760 ( .A(KEYINPUT29), .B(n687), .Z(n693) );
  XNOR2_X1 U761 ( .A(G2078), .B(KEYINPUT25), .ZN(n688) );
  XNOR2_X1 U762 ( .A(n688), .B(KEYINPUT95), .ZN(n1009) );
  NOR2_X1 U763 ( .A1(n1009), .A2(n705), .ZN(n691) );
  NOR2_X1 U764 ( .A1(n689), .A2(G1961), .ZN(n690) );
  NOR2_X1 U765 ( .A1(n691), .A2(n690), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n697), .A2(G301), .ZN(n692) );
  NOR2_X1 U767 ( .A1(n693), .A2(n692), .ZN(n702) );
  NAND2_X1 U768 ( .A1(G8), .A2(n705), .ZN(n746) );
  NOR2_X1 U769 ( .A1(G1966), .A2(n746), .ZN(n718) );
  NOR2_X1 U770 ( .A1(G2084), .A2(n705), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n718), .A2(n715), .ZN(n694) );
  NAND2_X1 U772 ( .A1(G8), .A2(n694), .ZN(n695) );
  XNOR2_X1 U773 ( .A(KEYINPUT30), .B(n695), .ZN(n696) );
  NOR2_X1 U774 ( .A1(G168), .A2(n696), .ZN(n699) );
  AND2_X1 U775 ( .A1(G301), .A2(n697), .ZN(n698) );
  NOR2_X1 U776 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U777 ( .A(n700), .B(KEYINPUT31), .ZN(n701) );
  NAND2_X1 U778 ( .A1(n716), .A2(G286), .ZN(n713) );
  INV_X1 U779 ( .A(G8), .ZN(n711) );
  NOR2_X1 U780 ( .A1(G1971), .A2(n746), .ZN(n707) );
  NOR2_X1 U781 ( .A1(G2090), .A2(n705), .ZN(n706) );
  NOR2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U783 ( .A(KEYINPUT99), .B(n708), .Z(n709) );
  NAND2_X1 U784 ( .A1(n709), .A2(G303), .ZN(n710) );
  OR2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U787 ( .A(KEYINPUT32), .B(n714), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G8), .A2(n715), .ZN(n720) );
  INV_X1 U789 ( .A(n716), .ZN(n717) );
  NOR2_X1 U790 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n744) );
  NOR2_X1 U793 ( .A1(G1971), .A2(G303), .ZN(n723) );
  NOR2_X1 U794 ( .A1(G1976), .A2(G288), .ZN(n922) );
  NOR2_X1 U795 ( .A1(n723), .A2(n922), .ZN(n724) );
  NAND2_X1 U796 ( .A1(n744), .A2(n724), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n923), .A2(n725), .ZN(n726) );
  INV_X1 U798 ( .A(n746), .ZN(n729) );
  INV_X1 U799 ( .A(KEYINPUT33), .ZN(n734) );
  NAND2_X1 U800 ( .A1(n922), .A2(n729), .ZN(n727) );
  NOR2_X1 U801 ( .A1(n734), .A2(n727), .ZN(n728) );
  XNOR2_X1 U802 ( .A(n728), .B(KEYINPUT101), .ZN(n733) );
  AND2_X1 U803 ( .A1(n729), .A2(n733), .ZN(n731) );
  XNOR2_X1 U804 ( .A(G1981), .B(G305), .ZN(n939) );
  INV_X1 U805 ( .A(n939), .ZN(n730) );
  AND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U807 ( .A1(n521), .A2(n732), .ZN(n751) );
  INV_X1 U808 ( .A(n733), .ZN(n735) );
  OR2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U810 ( .A1(n939), .A2(n736), .ZN(n741) );
  NOR2_X1 U811 ( .A1(G1981), .A2(G305), .ZN(n737) );
  XOR2_X1 U812 ( .A(n737), .B(KEYINPUT24), .Z(n738) );
  NOR2_X1 U813 ( .A1(n746), .A2(n738), .ZN(n739) );
  XNOR2_X1 U814 ( .A(n739), .B(KEYINPUT94), .ZN(n740) );
  NOR2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n749) );
  NOR2_X1 U816 ( .A1(G2090), .A2(G303), .ZN(n742) );
  NAND2_X1 U817 ( .A1(G8), .A2(n742), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n747), .B(KEYINPUT102), .ZN(n748) );
  AND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n750) );
  AND2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n759) );
  XNOR2_X1 U823 ( .A(G1986), .B(G290), .ZN(n936) );
  NAND2_X1 U824 ( .A1(n752), .A2(n936), .ZN(n757) );
  INV_X1 U825 ( .A(n753), .ZN(n755) );
  AND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U828 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U829 ( .A1(n761), .A2(n760), .ZN(n764) );
  AND2_X1 U830 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U831 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n766) );
  NAND2_X1 U832 ( .A1(G123), .A2(n884), .ZN(n765) );
  XNOR2_X1 U833 ( .A(n766), .B(n765), .ZN(n770) );
  NAND2_X1 U834 ( .A1(G111), .A2(n885), .ZN(n768) );
  NAND2_X1 U835 ( .A1(G99), .A2(n600), .ZN(n767) );
  NAND2_X1 U836 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U837 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U838 ( .A1(n605), .A2(G135), .ZN(n771) );
  NAND2_X1 U839 ( .A1(n772), .A2(n771), .ZN(n980) );
  XNOR2_X1 U840 ( .A(G2096), .B(n980), .ZN(n773) );
  OR2_X1 U841 ( .A1(G2100), .A2(n773), .ZN(G156) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U846 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U847 ( .A(G223), .ZN(n827) );
  NAND2_X1 U848 ( .A1(n827), .A2(G567), .ZN(n775) );
  XNOR2_X1 U849 ( .A(n775), .B(KEYINPUT11), .ZN(n776) );
  XNOR2_X1 U850 ( .A(KEYINPUT71), .B(n776), .ZN(G234) );
  INV_X1 U851 ( .A(G860), .ZN(n782) );
  OR2_X1 U852 ( .A1(n925), .A2(n782), .ZN(G153) );
  NOR2_X1 U853 ( .A1(n920), .A2(G868), .ZN(n777) );
  XNOR2_X1 U854 ( .A(n777), .B(KEYINPUT75), .ZN(n779) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n778) );
  NAND2_X1 U856 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U857 ( .A(G868), .ZN(n811) );
  NOR2_X1 U858 ( .A1(G286), .A2(n811), .ZN(n781) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n780) );
  NOR2_X1 U860 ( .A1(n781), .A2(n780), .ZN(G297) );
  NAND2_X1 U861 ( .A1(n782), .A2(G559), .ZN(n783) );
  NAND2_X1 U862 ( .A1(n783), .A2(n920), .ZN(n784) );
  XNOR2_X1 U863 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U864 ( .A1(G868), .A2(n925), .ZN(n785) );
  XOR2_X1 U865 ( .A(KEYINPUT77), .B(n785), .Z(n788) );
  NAND2_X1 U866 ( .A1(G868), .A2(n920), .ZN(n786) );
  NOR2_X1 U867 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U868 ( .A1(n788), .A2(n787), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G559), .A2(n920), .ZN(n789) );
  XOR2_X1 U870 ( .A(n925), .B(n789), .Z(n808) );
  XNOR2_X1 U871 ( .A(KEYINPUT79), .B(n808), .ZN(n790) );
  NOR2_X1 U872 ( .A1(G860), .A2(n790), .ZN(n802) );
  NAND2_X1 U873 ( .A1(G93), .A2(n791), .ZN(n792) );
  XNOR2_X1 U874 ( .A(n792), .B(KEYINPUT80), .ZN(n801) );
  NAND2_X1 U875 ( .A1(G67), .A2(n669), .ZN(n795) );
  NAND2_X1 U876 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U877 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U878 ( .A1(G80), .A2(n796), .ZN(n797) );
  XNOR2_X1 U879 ( .A(KEYINPUT81), .B(n797), .ZN(n798) );
  NOR2_X1 U880 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U881 ( .A1(n801), .A2(n800), .ZN(n810) );
  XOR2_X1 U882 ( .A(n802), .B(n810), .Z(G145) );
  XNOR2_X1 U883 ( .A(G166), .B(KEYINPUT19), .ZN(n807) );
  XOR2_X1 U884 ( .A(G305), .B(G290), .Z(n803) );
  XNOR2_X1 U885 ( .A(n810), .B(n803), .ZN(n804) );
  XNOR2_X1 U886 ( .A(n804), .B(G288), .ZN(n805) );
  XNOR2_X1 U887 ( .A(n805), .B(G299), .ZN(n806) );
  XNOR2_X1 U888 ( .A(n807), .B(n806), .ZN(n897) );
  XNOR2_X1 U889 ( .A(n897), .B(n808), .ZN(n809) );
  NAND2_X1 U890 ( .A1(n809), .A2(G868), .ZN(n813) );
  NAND2_X1 U891 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U892 ( .A1(n813), .A2(n812), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2078), .A2(G2084), .ZN(n814) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(n814), .Z(n815) );
  NAND2_X1 U895 ( .A1(G2090), .A2(n815), .ZN(n816) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n816), .ZN(n817) );
  NAND2_X1 U897 ( .A1(n817), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U898 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U899 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U900 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U901 ( .A1(G108), .A2(n819), .ZN(n834) );
  NAND2_X1 U902 ( .A1(n834), .A2(G567), .ZN(n825) );
  NOR2_X1 U903 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U905 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G96), .A2(n822), .ZN(n833) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n833), .ZN(n823) );
  XNOR2_X1 U908 ( .A(KEYINPUT82), .B(n823), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n825), .A2(n824), .ZN(n835) );
  NAND2_X1 U910 ( .A1(G661), .A2(G483), .ZN(n826) );
  NOR2_X1 U911 ( .A1(n835), .A2(n826), .ZN(n832) );
  NAND2_X1 U912 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n827), .ZN(G217) );
  INV_X1 U914 ( .A(G661), .ZN(n829) );
  NAND2_X1 U915 ( .A1(G2), .A2(G15), .ZN(n828) );
  NOR2_X1 U916 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U917 ( .A(KEYINPUT108), .B(n830), .Z(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n835), .ZN(G319) );
  XNOR2_X1 U927 ( .A(G1991), .B(G2474), .ZN(n845) );
  XOR2_X1 U928 ( .A(G1956), .B(G1966), .Z(n837) );
  XNOR2_X1 U929 ( .A(G1996), .B(G1981), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U931 ( .A(G1986), .B(G1961), .Z(n839) );
  XNOR2_X1 U932 ( .A(G1976), .B(G1971), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U935 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U937 ( .A(n845), .B(n844), .ZN(G229) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2072), .ZN(n846) );
  XNOR2_X1 U939 ( .A(n846), .B(KEYINPUT109), .ZN(n856) );
  XOR2_X1 U940 ( .A(KEYINPUT110), .B(G2100), .Z(n848) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U943 ( .A(G2096), .B(G2090), .Z(n850) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2084), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U946 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U947 ( .A(KEYINPUT43), .B(G2678), .ZN(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U949 ( .A(n856), .B(n855), .ZN(G227) );
  NAND2_X1 U950 ( .A1(G112), .A2(n885), .ZN(n858) );
  NAND2_X1 U951 ( .A1(G136), .A2(n605), .ZN(n857) );
  NAND2_X1 U952 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U953 ( .A1(n884), .A2(G124), .ZN(n859) );
  XNOR2_X1 U954 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U955 ( .A1(G100), .A2(n600), .ZN(n860) );
  NAND2_X1 U956 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U957 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n865) );
  XNOR2_X1 U959 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n865), .B(n864), .ZN(n874) );
  NAND2_X1 U961 ( .A1(G130), .A2(n884), .ZN(n867) );
  NAND2_X1 U962 ( .A1(G118), .A2(n885), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U964 ( .A1(G106), .A2(n600), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G142), .A2(n605), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(n870), .B(KEYINPUT45), .Z(n871) );
  NOR2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U969 ( .A(n874), .B(n873), .Z(n875) );
  XNOR2_X1 U970 ( .A(G162), .B(n875), .ZN(n879) );
  XNOR2_X1 U971 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U972 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U973 ( .A(n980), .B(n880), .ZN(n883) );
  XOR2_X1 U974 ( .A(n881), .B(G164), .Z(n882) );
  XNOR2_X1 U975 ( .A(n883), .B(n882), .ZN(n895) );
  NAND2_X1 U976 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U977 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U978 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U979 ( .A(n888), .B(KEYINPUT47), .ZN(n890) );
  NAND2_X1 U980 ( .A1(G103), .A2(n600), .ZN(n889) );
  NAND2_X1 U981 ( .A1(n890), .A2(n889), .ZN(n893) );
  NAND2_X1 U982 ( .A1(G139), .A2(n605), .ZN(n891) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(n891), .ZN(n892) );
  NOR2_X1 U984 ( .A1(n893), .A2(n892), .ZN(n973) );
  XOR2_X1 U985 ( .A(n973), .B(G160), .Z(n894) );
  XNOR2_X1 U986 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U987 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n925), .B(n897), .ZN(n899) );
  XNOR2_X1 U989 ( .A(G171), .B(n920), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U991 ( .A(n900), .B(G286), .ZN(n901) );
  NOR2_X1 U992 ( .A1(G37), .A2(n901), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2443), .B(KEYINPUT106), .Z(n903) );
  XNOR2_X1 U994 ( .A(G2451), .B(G2427), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U996 ( .A(n904), .B(G2430), .Z(n906) );
  XNOR2_X1 U997 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U998 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U999 ( .A(KEYINPUT107), .B(G2438), .Z(n908) );
  XNOR2_X1 U1000 ( .A(G2435), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1002 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1003 ( .A(G2446), .B(KEYINPUT105), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .Z(n946) );
  XNOR2_X1 U1016 ( .A(n920), .B(G1348), .ZN(n934) );
  XNOR2_X1 U1017 ( .A(G1961), .B(G171), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n921), .B(KEYINPUT122), .ZN(n929) );
  INV_X1 U1019 ( .A(n922), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(G1341), .B(n925), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G1956), .B(G299), .Z(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT123), .B(n930), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n944) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G303), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(n935), .B(KEYINPUT124), .ZN(n937) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n942) );
  XOR2_X1 U1031 ( .A(G1966), .B(G168), .Z(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1033 ( .A(KEYINPUT57), .B(n940), .Z(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(KEYINPUT125), .B(n947), .ZN(n1004) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G21), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(G5), .B(G1961), .ZN(n948) );
  NOR2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n960) );
  XNOR2_X1 U1041 ( .A(G1981), .B(G6), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1044 ( .A(KEYINPUT126), .B(G4), .Z(n953) );
  XNOR2_X1 U1045 ( .A(G1348), .B(KEYINPUT59), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n953), .B(n952), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G20), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1050 ( .A(KEYINPUT60), .B(n958), .Z(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n968) );
  XNOR2_X1 U1052 ( .A(G1976), .B(G23), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(G1986), .B(G24), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n963), .B(KEYINPUT127), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT61), .B(n969), .ZN(n971) );
  INV_X1 U1061 ( .A(G16), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G11), .ZN(n1002) );
  XNOR2_X1 U1064 ( .A(G164), .B(G2078), .ZN(n976) );
  XOR2_X1 U1065 ( .A(G2072), .B(n973), .Z(n974) );
  XNOR2_X1 U1066 ( .A(KEYINPUT117), .B(n974), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n977), .B(KEYINPUT50), .ZN(n995) );
  XOR2_X1 U1069 ( .A(G160), .B(G2084), .Z(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n991) );
  XOR2_X1 U1072 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1074 ( .A(KEYINPUT116), .B(n984), .Z(n985) );
  XOR2_X1 U1075 ( .A(KEYINPUT51), .B(n985), .Z(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1081 ( .A(KEYINPUT52), .B(n996), .Z(n997) );
  NOR2_X1 U1082 ( .A1(KEYINPUT55), .A2(n997), .ZN(n998) );
  XOR2_X1 U1083 ( .A(KEYINPUT118), .B(n998), .Z(n999) );
  NAND2_X1 U1084 ( .A1(n999), .A2(G29), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(KEYINPUT119), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1086 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1087 ( .A1(n1004), .A2(n1003), .ZN(n1026) );
  XOR2_X1 U1088 ( .A(G2072), .B(G33), .Z(n1005) );
  NAND2_X1 U1089 ( .A1(n1005), .A2(G28), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G26), .B(G2067), .ZN(n1006) );
  NOR2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1016) );
  XNOR2_X1 U1092 ( .A(G1991), .B(G25), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(n1008), .B(KEYINPUT120), .ZN(n1014) );
  XNOR2_X1 U1094 ( .A(G1996), .B(G32), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(n1009), .B(G27), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(KEYINPUT121), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1099 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(n1017), .B(KEYINPUT53), .ZN(n1020) );
  XOR2_X1 U1101 ( .A(G2084), .B(G34), .Z(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT54), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1104 ( .A(G35), .B(G2090), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT55), .B(n1023), .Z(n1024) );
  NOR2_X1 U1107 ( .A1(G29), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(n1027), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

