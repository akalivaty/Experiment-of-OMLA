

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n451), .B(n450), .ZN(n527) );
  XOR2_X2 U322 ( .A(KEYINPUT41), .B(n383), .Z(n546) );
  XOR2_X1 U323 ( .A(n352), .B(n351), .Z(n289) );
  NOR2_X1 U324 ( .A1(n551), .A2(n388), .ZN(n389) );
  XNOR2_X1 U325 ( .A(n321), .B(KEYINPUT10), .ZN(n322) );
  NOR2_X1 U326 ( .A1(n516), .A2(n413), .ZN(n414) );
  XNOR2_X1 U327 ( .A(n323), .B(n322), .ZN(n327) );
  NAND2_X1 U328 ( .A1(n452), .A2(n527), .ZN(n563) );
  XNOR2_X1 U329 ( .A(KEYINPUT78), .B(n555), .ZN(n536) );
  XNOR2_X1 U330 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n291) );
  XNOR2_X1 U333 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U335 ( .A(KEYINPUT89), .B(n292), .Z(n431) );
  XOR2_X1 U336 ( .A(G57GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U337 ( .A(G141GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U339 ( .A(G85GAT), .B(G162GAT), .Z(n296) );
  XNOR2_X1 U340 ( .A(G29GAT), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n311) );
  XOR2_X1 U343 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n300) );
  XNOR2_X1 U344 ( .A(KEYINPUT92), .B(KEYINPUT94), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n302) );
  XNOR2_X1 U347 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U350 ( .A(G113GAT), .B(G1GAT), .Z(n364) );
  XOR2_X1 U351 ( .A(G134GAT), .B(KEYINPUT0), .Z(n435) );
  XOR2_X1 U352 ( .A(n435), .B(KEYINPUT1), .Z(n306) );
  NAND2_X1 U353 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n364), .B(n307), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n431), .B(n312), .ZN(n516) );
  XOR2_X1 U359 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n314) );
  NAND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  XOR2_X1 U361 ( .A(n314), .B(n313), .Z(n316) );
  XNOR2_X1 U362 ( .A(G36GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n315), .B(G218GAT), .ZN(n403) );
  XNOR2_X1 U364 ( .A(n316), .B(n403), .ZN(n320) );
  XOR2_X1 U365 ( .A(G29GAT), .B(G43GAT), .Z(n318) );
  XNOR2_X1 U366 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n367) );
  XNOR2_X1 U368 ( .A(n367), .B(G134GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n323) );
  XOR2_X1 U370 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XOR2_X1 U371 ( .A(n426), .B(KEYINPUT9), .Z(n321) );
  XOR2_X1 U372 ( .A(KEYINPUT75), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G92GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U375 ( .A(G106GAT), .B(n326), .Z(n349) );
  XNOR2_X1 U376 ( .A(n327), .B(n349), .ZN(n555) );
  XNOR2_X1 U377 ( .A(KEYINPUT36), .B(n536), .ZN(n486) );
  XOR2_X1 U378 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n329) );
  NAND2_X1 U379 ( .A1(G231GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U381 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U385 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XOR2_X1 U386 ( .A(KEYINPUT80), .B(G64GAT), .Z(n335) );
  XNOR2_X1 U387 ( .A(G1GAT), .B(G78GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n439), .B(n336), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XOR2_X1 U392 ( .A(KEYINPUT13), .B(G57GAT), .Z(n350) );
  XOR2_X1 U393 ( .A(n396), .B(n350), .Z(n340) );
  XNOR2_X1 U394 ( .A(G71GAT), .B(G211GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(n342), .B(n341), .Z(n344) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G155GAT), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n551) );
  NAND2_X1 U399 ( .A1(n486), .A2(n551), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n345), .B(KEYINPUT45), .ZN(n346) );
  XNOR2_X1 U401 ( .A(KEYINPUT65), .B(n346), .ZN(n381) );
  XOR2_X1 U402 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n348) );
  XNOR2_X1 U403 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n360) );
  XOR2_X1 U405 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XNOR2_X1 U406 ( .A(n436), .B(n349), .ZN(n358) );
  XOR2_X1 U407 ( .A(KEYINPUT77), .B(n350), .Z(n352) );
  XOR2_X1 U408 ( .A(G176GAT), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U409 ( .A(G204GAT), .B(n399), .ZN(n351) );
  XNOR2_X1 U410 ( .A(G78GAT), .B(KEYINPUT74), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n353), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U412 ( .A(n418), .B(KEYINPUT76), .ZN(n355) );
  AND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n289), .B(n356), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n383) );
  BUF_X1 U418 ( .A(n383), .Z(n572) );
  XOR2_X1 U419 ( .A(KEYINPUT70), .B(G197GAT), .Z(n362) );
  XNOR2_X1 U420 ( .A(G36GAT), .B(G50GAT), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U422 ( .A(n363), .B(G15GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(n364), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U425 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XOR2_X1 U426 ( .A(n367), .B(n427), .Z(n369) );
  NAND2_X1 U427 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U429 ( .A(n371), .B(n370), .Z(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n373) );
  XNOR2_X1 U431 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U433 ( .A(G8GAT), .B(KEYINPUT67), .Z(n375) );
  XNOR2_X1 U434 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n567) );
  INV_X1 U438 ( .A(n567), .ZN(n544) );
  NOR2_X1 U439 ( .A1(n572), .A2(n544), .ZN(n380) );
  AND2_X1 U440 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n382), .B(KEYINPUT113), .ZN(n391) );
  INV_X1 U442 ( .A(n555), .ZN(n387) );
  XNOR2_X1 U443 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n385) );
  INV_X1 U444 ( .A(n546), .ZN(n560) );
  NOR2_X1 U445 ( .A1(n567), .A2(n560), .ZN(n384) );
  XOR2_X1 U446 ( .A(n385), .B(n384), .Z(n386) );
  NAND2_X1 U447 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U448 ( .A(KEYINPUT47), .B(n389), .ZN(n390) );
  NAND2_X1 U449 ( .A1(n391), .A2(n390), .ZN(n393) );
  XNOR2_X1 U450 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n392) );
  XNOR2_X2 U451 ( .A(n393), .B(n392), .ZN(n540) );
  XOR2_X1 U452 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n395) );
  XNOR2_X1 U453 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n443) );
  XNOR2_X1 U455 ( .A(G92GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n397), .B(KEYINPUT96), .ZN(n398) );
  XOR2_X1 U457 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U460 ( .A(n402), .B(KEYINPUT97), .Z(n405) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT98), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n443), .B(n406), .ZN(n410) );
  XOR2_X1 U464 ( .A(G204GAT), .B(G211GAT), .Z(n408) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n419) );
  INV_X1 U467 ( .A(n419), .ZN(n409) );
  XOR2_X1 U468 ( .A(n410), .B(n409), .Z(n478) );
  INV_X1 U469 ( .A(n478), .ZN(n518) );
  NAND2_X1 U470 ( .A1(n540), .A2(n518), .ZN(n412) );
  XOR2_X1 U471 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(KEYINPUT64), .ZN(n566) );
  XOR2_X1 U474 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n416) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U477 ( .A(n417), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U480 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n423) );
  XNOR2_X1 U481 ( .A(G218GAT), .B(G106GAT), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U483 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n470) );
  NAND2_X1 U487 ( .A1(n566), .A2(n470), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n432), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U489 ( .A(G183GAT), .B(G176GAT), .Z(n434) );
  XNOR2_X1 U490 ( .A(G113GAT), .B(G99GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n451) );
  XOR2_X1 U492 ( .A(G190GAT), .B(n435), .Z(n438) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n449) );
  XOR2_X1 U496 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n442) );
  XNOR2_X1 U497 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U499 ( .A(n443), .B(KEYINPUT20), .Z(n445) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U504 ( .A(n563), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n453), .A2(n536), .ZN(n455) );
  NOR2_X1 U506 ( .A1(n567), .A2(n563), .ZN(n458) );
  XNOR2_X1 U507 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n456) );
  XNOR2_X1 U508 ( .A(n456), .B(G169GAT), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(G1348GAT) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n460) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(n477) );
  INV_X1 U513 ( .A(n516), .ZN(n475) );
  NOR2_X1 U514 ( .A1(n567), .A2(n572), .ZN(n490) );
  NAND2_X1 U515 ( .A1(n527), .A2(n518), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n470), .A2(n461), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n462), .ZN(n467) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n518), .ZN(n469) );
  NOR2_X1 U519 ( .A1(n527), .A2(n470), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT26), .B(n463), .Z(n464) );
  XNOR2_X1 U521 ( .A(KEYINPUT99), .B(n464), .ZN(n565) );
  NAND2_X1 U522 ( .A1(n469), .A2(n565), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT100), .B(n465), .Z(n466) );
  NOR2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n468), .A2(n516), .ZN(n472) );
  AND2_X1 U526 ( .A1(n516), .A2(n469), .ZN(n541) );
  XNOR2_X1 U527 ( .A(KEYINPUT28), .B(n470), .ZN(n498) );
  NAND2_X1 U528 ( .A1(n541), .A2(n498), .ZN(n529) );
  NOR2_X1 U529 ( .A1(n529), .A2(n527), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n487) );
  INV_X1 U531 ( .A(n551), .ZN(n578) );
  NOR2_X1 U532 ( .A1(n536), .A2(n578), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U534 ( .A1(n487), .A2(n474), .ZN(n503) );
  NAND2_X1 U535 ( .A1(n490), .A2(n503), .ZN(n484) );
  NOR2_X1 U536 ( .A1(n475), .A2(n484), .ZN(n476) );
  XOR2_X1 U537 ( .A(n477), .B(n476), .Z(G1324GAT) );
  NOR2_X1 U538 ( .A1(n478), .A2(n484), .ZN(n479) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  INV_X1 U540 ( .A(n527), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n480), .A2(n484), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U544 ( .A(G15GAT), .B(n483), .Z(G1326GAT) );
  NOR2_X1 U545 ( .A1(n498), .A2(n484), .ZN(n485) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NOR2_X1 U548 ( .A1(n551), .A2(n487), .ZN(n488) );
  NAND2_X1 U549 ( .A1(n486), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT37), .ZN(n513) );
  NAND2_X1 U551 ( .A1(n490), .A2(n513), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT38), .B(n491), .Z(n499) );
  NAND2_X1 U553 ( .A1(n499), .A2(n516), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n499), .A2(n518), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n527), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  XOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT105), .Z(n501) );
  INV_X1 U562 ( .A(n498), .ZN(n522) );
  NAND2_X1 U563 ( .A1(n499), .A2(n522), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U565 ( .A1(n544), .A2(n560), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT106), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n503), .A2(n514), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT107), .B(n504), .ZN(n509) );
  NAND2_X1 U569 ( .A1(n516), .A2(n509), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n518), .A2(n509), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n527), .A2(n509), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U577 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(KEYINPUT109), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n527), .A2(n523), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT115), .Z(n531) );
  NAND2_X1 U594 ( .A1(n527), .A2(n540), .ZN(n528) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n537), .A2(n544), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U599 ( .A1(n537), .A2(n546), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n537), .A2(n551), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  INV_X1 U607 ( .A(n540), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n565), .ZN(n542) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n554), .A2(n544), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U614 ( .A1(n554), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT117), .Z(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT118), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n559) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n560), .A2(n563), .ZN(n561) );
  XOR2_X1 U627 ( .A(n562), .B(n561), .Z(G1349GAT) );
  NOR2_X1 U628 ( .A1(n578), .A2(n563), .ZN(n564) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n564), .Z(G1350GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n567), .A2(n577), .ZN(n569) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  INV_X1 U636 ( .A(n577), .ZN(n580) );
  AND2_X1 U637 ( .A1(n580), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NAND2_X1 U644 ( .A1(n486), .A2(n580), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XOR2_X1 U646 ( .A(n582), .B(KEYINPUT126), .Z(n584) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1355GAT) );
endmodule

