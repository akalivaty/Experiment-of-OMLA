

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U324 ( .A(n330), .B(n329), .Z(n291) );
  INV_X1 U325 ( .A(KEYINPUT111), .ZN(n384) );
  XNOR2_X1 U326 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n349) );
  XNOR2_X1 U327 ( .A(n384), .B(KEYINPUT47), .ZN(n385) );
  XNOR2_X1 U328 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U329 ( .A(n341), .B(n324), .ZN(n325) );
  XNOR2_X1 U330 ( .A(n331), .B(n291), .ZN(n332) );
  XOR2_X1 U331 ( .A(n357), .B(n356), .Z(n466) );
  XNOR2_X1 U332 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U333 ( .A(KEYINPUT124), .B(n447), .Z(n583) );
  NOR2_X1 U334 ( .A1(n539), .A2(n455), .ZN(n575) );
  XOR2_X1 U335 ( .A(n566), .B(KEYINPUT77), .Z(n574) );
  XNOR2_X1 U336 ( .A(n448), .B(KEYINPUT126), .ZN(n449) );
  XNOR2_X1 U337 ( .A(n457), .B(G176GAT), .ZN(n458) );
  XNOR2_X1 U338 ( .A(n450), .B(n449), .ZN(G1354GAT) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U340 ( .A(G78GAT), .B(G211GAT), .Z(n293) );
  XNOR2_X1 U341 ( .A(G127GAT), .B(G155GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U343 ( .A(G71GAT), .B(KEYINPUT13), .Z(n342) );
  XOR2_X1 U344 ( .A(G8GAT), .B(KEYINPUT78), .Z(n321) );
  XOR2_X1 U345 ( .A(n342), .B(n321), .Z(n295) );
  NAND2_X1 U346 ( .A1(G231GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U348 ( .A(G64GAT), .B(KEYINPUT15), .Z(n297) );
  XNOR2_X1 U349 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U351 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U352 ( .A(G22GAT), .B(G15GAT), .Z(n366) );
  XOR2_X1 U353 ( .A(KEYINPUT14), .B(G57GAT), .Z(n301) );
  XNOR2_X1 U354 ( .A(G1GAT), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n366), .B(n302), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(n306), .B(n305), .Z(n494) );
  XOR2_X1 U359 ( .A(G176GAT), .B(G64GAT), .Z(n352) );
  XNOR2_X1 U360 ( .A(G204GAT), .B(n352), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n307), .B(KEYINPUT90), .ZN(n310) );
  XOR2_X1 U362 ( .A(G92GAT), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n326) );
  XOR2_X1 U365 ( .A(n310), .B(n326), .Z(n319) );
  XOR2_X1 U366 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n312) );
  XNOR2_X1 U367 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(n313), .B(KEYINPUT19), .Z(n315) );
  XNOR2_X1 U370 ( .A(G169GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n416) );
  XOR2_X1 U372 ( .A(G211GAT), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n404) );
  XNOR2_X1 U375 ( .A(n416), .B(n404), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U377 ( .A(n321), .B(n320), .Z(n323) );
  NAND2_X1 U378 ( .A1(G226GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n471) );
  XNOR2_X1 U380 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n390) );
  XOR2_X1 U381 ( .A(KEYINPUT36), .B(KEYINPUT98), .Z(n339) );
  XOR2_X1 U382 ( .A(G99GAT), .B(G106GAT), .Z(n341) );
  AND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n324) );
  INV_X1 U384 ( .A(KEYINPUT76), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U386 ( .A(G50GAT), .B(G162GAT), .Z(n400) );
  XNOR2_X1 U387 ( .A(n400), .B(KEYINPUT75), .ZN(n331) );
  XOR2_X1 U388 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n330) );
  XNOR2_X1 U389 ( .A(KEYINPUT74), .B(KEYINPUT11), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT7), .B(G43GAT), .Z(n335) );
  XNOR2_X1 U391 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n368) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(G134GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n336), .B(G85GAT), .ZN(n435) );
  XNOR2_X1 U395 ( .A(n368), .B(n435), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n566) );
  XNOR2_X1 U397 ( .A(n339), .B(n574), .ZN(n582) );
  NOR2_X1 U398 ( .A1(n494), .A2(n582), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n340), .B(KEYINPUT45), .ZN(n377) );
  XOR2_X1 U400 ( .A(n342), .B(n341), .Z(n344) );
  XOR2_X1 U401 ( .A(G204GAT), .B(G78GAT), .Z(n399) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G57GAT), .Z(n439) );
  XNOR2_X1 U403 ( .A(n399), .B(n439), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n357) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n346) );
  XNOR2_X1 U406 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n348) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n351) );
  XOR2_X1 U410 ( .A(n349), .B(KEYINPUT33), .Z(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U412 ( .A(n353), .B(n352), .Z(n355) );
  XNOR2_X1 U413 ( .A(G85GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(KEYINPUT67), .B(G8GAT), .Z(n359) );
  XNOR2_X1 U416 ( .A(G169GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n361) );
  XNOR2_X1 U419 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n375) );
  XOR2_X1 U422 ( .A(G197GAT), .B(G50GAT), .Z(n365) );
  XNOR2_X1 U423 ( .A(G29GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U425 ( .A(n367), .B(n366), .Z(n373) );
  XOR2_X1 U426 ( .A(n368), .B(KEYINPUT68), .Z(n370) );
  NAND2_X1 U427 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U429 ( .A(G113GAT), .B(G1GAT), .Z(n441) );
  XNOR2_X1 U430 ( .A(n371), .B(n441), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n569) );
  INV_X1 U433 ( .A(n569), .ZN(n578) );
  AND2_X1 U434 ( .A1(n466), .A2(n578), .ZN(n376) );
  AND2_X1 U435 ( .A1(n377), .A2(n376), .ZN(n378) );
  XOR2_X1 U436 ( .A(KEYINPUT112), .B(n378), .Z(n388) );
  XNOR2_X1 U437 ( .A(KEYINPUT41), .B(n466), .ZN(n456) );
  NAND2_X1 U438 ( .A1(n456), .A2(n569), .ZN(n380) );
  INV_X1 U439 ( .A(KEYINPUT46), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  INV_X1 U441 ( .A(n494), .ZN(n571) );
  NOR2_X1 U442 ( .A1(n381), .A2(n571), .ZN(n382) );
  XOR2_X1 U443 ( .A(n382), .B(KEYINPUT110), .Z(n383) );
  NOR2_X1 U444 ( .A1(n566), .A2(n383), .ZN(n386) );
  NAND2_X1 U445 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n537) );
  NAND2_X1 U447 ( .A1(n471), .A2(n537), .ZN(n392) );
  XOR2_X1 U448 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n453) );
  XOR2_X1 U450 ( .A(KEYINPUT3), .B(G148GAT), .Z(n394) );
  XNOR2_X1 U451 ( .A(G141GAT), .B(G155GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U453 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n430) );
  XOR2_X1 U455 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n398) );
  XNOR2_X1 U456 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n411) );
  XOR2_X1 U458 ( .A(G106GAT), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U461 ( .A(n403), .B(KEYINPUT24), .Z(n409) );
  XOR2_X1 U462 ( .A(n404), .B(KEYINPUT87), .Z(n406) );
  NAND2_X1 U463 ( .A1(G228GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U465 ( .A(G22GAT), .B(n407), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n412) );
  XNOR2_X1 U468 ( .A(n430), .B(n412), .ZN(n473) );
  XOR2_X1 U469 ( .A(G120GAT), .B(KEYINPUT20), .Z(n414) );
  XNOR2_X1 U470 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n427) );
  XNOR2_X1 U473 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n417), .B(KEYINPUT0), .ZN(n440) );
  XOR2_X1 U475 ( .A(G134GAT), .B(n440), .Z(n419) );
  XNOR2_X1 U476 ( .A(G43GAT), .B(G190GAT), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n420), .B(G99GAT), .Z(n425) );
  XOR2_X1 U479 ( .A(G176GAT), .B(G71GAT), .Z(n422) );
  NAND2_X1 U480 ( .A1(G227GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U482 ( .A(G113GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n539) );
  NAND2_X1 U485 ( .A1(n473), .A2(n539), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n428), .B(KEYINPUT92), .ZN(n429) );
  XNOR2_X1 U487 ( .A(KEYINPUT26), .B(n429), .ZN(n555) );
  INV_X1 U488 ( .A(n430), .ZN(n434) );
  XOR2_X1 U489 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n432) );
  XNOR2_X1 U490 ( .A(G162GAT), .B(KEYINPUT6), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n445) );
  XOR2_X1 U493 ( .A(n435), .B(KEYINPUT1), .Z(n437) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U496 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n479) );
  XNOR2_X1 U500 ( .A(KEYINPUT89), .B(n479), .ZN(n526) );
  INV_X1 U501 ( .A(n526), .ZN(n451) );
  NOR2_X1 U502 ( .A1(n555), .A2(n451), .ZN(n446) );
  AND2_X1 U503 ( .A1(n453), .A2(n446), .ZN(n447) );
  NOR2_X1 U504 ( .A1(n494), .A2(n583), .ZN(n450) );
  INV_X1 U505 ( .A(G211GAT), .ZN(n448) );
  NOR2_X1 U506 ( .A1(n451), .A2(n473), .ZN(n452) );
  AND2_X1 U507 ( .A1(n453), .A2(n452), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n575), .A2(n456), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  INV_X1 U511 ( .A(G204GAT), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n466), .A2(n583), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(G1353GAT) );
  XOR2_X1 U516 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n465) );
  XNOR2_X1 U517 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(n486) );
  NAND2_X1 U519 ( .A1(n466), .A2(n569), .ZN(n467) );
  XNOR2_X1 U520 ( .A(n467), .B(KEYINPUT73), .ZN(n498) );
  XNOR2_X1 U521 ( .A(n473), .B(KEYINPUT28), .ZN(n542) );
  XOR2_X1 U522 ( .A(n471), .B(KEYINPUT27), .Z(n470) );
  NOR2_X1 U523 ( .A1(n470), .A2(n526), .ZN(n538) );
  NAND2_X1 U524 ( .A1(n539), .A2(n538), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n542), .A2(n468), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT91), .B(n469), .Z(n481) );
  NOR2_X1 U527 ( .A1(n470), .A2(n555), .ZN(n477) );
  INV_X1 U528 ( .A(n471), .ZN(n528) );
  NOR2_X1 U529 ( .A1(n539), .A2(n528), .ZN(n472) );
  NOR2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT93), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT25), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U535 ( .A1(n481), .A2(n480), .ZN(n493) );
  NOR2_X1 U536 ( .A1(n494), .A2(n574), .ZN(n482) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n482), .Z(n483) );
  NOR2_X1 U538 ( .A1(n493), .A2(n483), .ZN(n513) );
  NAND2_X1 U539 ( .A1(n498), .A2(n513), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT94), .B(n484), .ZN(n491) );
  NOR2_X1 U541 ( .A1(n491), .A2(n526), .ZN(n485) );
  XOR2_X1 U542 ( .A(n486), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n491), .A2(n528), .ZN(n488) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  NOR2_X1 U547 ( .A1(n539), .A2(n491), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  INV_X1 U549 ( .A(n542), .ZN(n534) );
  NOR2_X1 U550 ( .A1(n534), .A2(n491), .ZN(n492) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n492), .Z(G1327GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT37), .B(KEYINPUT99), .Z(n497) );
  NOR2_X1 U553 ( .A1(n493), .A2(n582), .ZN(n495) );
  NAND2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n525) );
  NAND2_X1 U556 ( .A1(n498), .A2(n525), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(KEYINPUT100), .ZN(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT38), .B(n500), .ZN(n509) );
  NOR2_X1 U559 ( .A1(n526), .A2(n509), .ZN(n502) );
  XNOR2_X1 U560 ( .A(KEYINPUT39), .B(KEYINPUT101), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U562 ( .A(G29GAT), .B(n503), .Z(G1328GAT) );
  NOR2_X1 U563 ( .A1(n528), .A2(n509), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT102), .B(n504), .Z(n505) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  NOR2_X1 U566 ( .A1(n539), .A2(n509), .ZN(n507) );
  XNOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n534), .A2(n509), .ZN(n510) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U572 ( .A(KEYINPUT104), .B(n511), .ZN(G1331GAT) );
  INV_X1 U573 ( .A(n456), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n569), .A2(n512), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n513), .A2(n524), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n526), .A2(n519), .ZN(n515) );
  XNOR2_X1 U577 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n528), .A2(n519), .ZN(n517) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n539), .A2(n519), .ZN(n518) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n518), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n534), .ZN(n523) );
  XOR2_X1 U585 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n521) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n533) );
  NOR2_X1 U590 ( .A1(n526), .A2(n533), .ZN(n527) );
  XOR2_X1 U591 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n533), .ZN(n529) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n539), .A2(n533), .ZN(n530) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n532) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n536) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U600 ( .A(n536), .B(n535), .Z(G1339GAT) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n554) );
  NOR2_X1 U603 ( .A1(n539), .A2(n554), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(KEYINPUT113), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n569), .A2(n551), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n546) );
  NAND2_X1 U609 ( .A1(n551), .A2(n456), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT115), .Z(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  NAND2_X1 U613 ( .A1(n571), .A2(n551), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT50), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n574), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n558) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT117), .B(n556), .Z(n567) );
  NAND2_X1 U622 ( .A1(n569), .A2(n567), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n560) );
  XNOR2_X1 U625 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n564) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n567), .A2(n456), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n571), .A2(n567), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n575), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U638 ( .A1(n575), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT58), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(n577), .ZN(G1351GAT) );
  NOR2_X1 U643 ( .A1(n583), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

