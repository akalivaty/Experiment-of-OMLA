//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n194), .A4(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n194), .B1(new_n191), .B2(new_n193), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n196), .A2(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n207), .A3(new_n210), .A4(new_n205), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(G134), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n210), .B1(new_n205), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n192), .A2(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n190), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G128), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n190), .A2(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n191), .A3(new_n193), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n214), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n201), .A2(new_n212), .B1(new_n223), .B2(new_n211), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT2), .B(G113), .Z(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G119), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT66), .A3(G116), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n226), .B2(G119), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n225), .A2(new_n227), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n227), .A3(new_n229), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n206), .A2(G134), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n203), .A2(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n221), .A2(new_n191), .A3(new_n193), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n220), .A2(new_n190), .A3(G143), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n221), .B2(new_n193), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n211), .B(new_n242), .C1(new_n243), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n212), .A2(new_n201), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n216), .A2(new_n218), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n222), .A2(new_n249), .A3(new_n244), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(KEYINPUT65), .A3(new_n211), .A4(new_n242), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT30), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n201), .A2(new_n212), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n253), .A2(KEYINPUT30), .A3(new_n246), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n239), .B1(new_n255), .B2(new_n236), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT31), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(G101), .ZN(new_n260));
  INV_X1    g074(.A(G210), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n261), .A2(G237), .A3(G953), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n260), .B(new_n262), .Z(new_n263));
  NAND4_X1  g077(.A1(new_n256), .A2(new_n257), .A3(new_n258), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n246), .A2(new_n247), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n253), .A2(new_n251), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n224), .A2(KEYINPUT30), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n236), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(new_n258), .A3(new_n238), .A4(new_n263), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n238), .A3(new_n263), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n238), .A2(KEYINPUT28), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n224), .A2(new_n276), .A3(new_n237), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n236), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n263), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n274), .A2(KEYINPUT31), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(KEYINPUT68), .B(new_n189), .C1(new_n273), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n287), .B2(new_n188), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n187), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n270), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n281), .B1(new_n290), .B2(new_n239), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n276), .B1(new_n224), .B2(new_n237), .ZN(new_n292));
  AND4_X1   g106(.A1(new_n276), .A2(new_n253), .A3(new_n237), .A4(new_n246), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n263), .B(new_n279), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n278), .A2(KEYINPUT69), .A3(new_n263), .A4(new_n279), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n291), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT70), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n278), .B1(new_n237), .B2(new_n224), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n302), .B2(new_n263), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n291), .A2(new_n296), .A3(new_n304), .A4(new_n297), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n299), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n189), .B1(new_n273), .B2(new_n282), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n306), .A2(G472), .B1(new_n307), .B2(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n289), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G140), .ZN(new_n310));
  INV_X1    g124(.A(G953), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G227), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G104), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(new_n315), .B2(G107), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G104), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(G107), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G101), .ZN(new_n322));
  INV_X1    g136(.A(G101), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n316), .A2(new_n319), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n326), .A3(G101), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n201), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n318), .A3(G104), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT78), .B1(new_n318), .B2(G104), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n315), .A2(G107), .ZN(new_n332));
  OAI211_X1 g146(.A(G101), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(new_n324), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT10), .A4(new_n250), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n250), .A2(new_n324), .A3(new_n333), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n328), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n212), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n212), .B(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n314), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n313), .B1(new_n341), .B2(new_n345), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT83), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n313), .C1(new_n341), .C2(new_n345), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n334), .A2(new_n250), .ZN(new_n354));
  INV_X1    g168(.A(new_n250), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n333), .A2(new_n324), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n354), .A2(new_n357), .B1(new_n209), .B2(new_n211), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(KEYINPUT12), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n250), .B1(new_n324), .B2(new_n333), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n212), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT12), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(KEYINPUT82), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n365), .A3(KEYINPUT12), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT12), .B(new_n212), .C1(new_n360), .C2(new_n361), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n359), .A2(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n347), .B1(new_n352), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G469), .ZN(new_n371));
  INV_X1    g185(.A(G902), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(new_n372), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n314), .B1(new_n369), .B2(new_n346), .ZN(new_n376));
  INV_X1    g190(.A(new_n348), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n342), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G469), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G214), .B1(G237), .B2(G902), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT84), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n201), .A2(G125), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n250), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT7), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(KEYINPUT87), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n311), .A2(G224), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n387), .A2(new_n390), .B1(KEYINPUT7), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(KEYINPUT7), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n393), .B(new_n389), .C1(new_n384), .C2(new_n386), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n325), .A2(new_n236), .A3(new_n327), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n228), .A3(G116), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n398), .A2(KEYINPUT85), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n231), .A2(new_n229), .A3(KEYINPUT5), .A4(new_n227), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(KEYINPUT85), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n399), .A2(new_n400), .A3(G113), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n334), .A2(new_n402), .A3(new_n232), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G122), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n404), .B(KEYINPUT8), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n232), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n356), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n395), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n396), .A2(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(new_n404), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n405), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n391), .B(KEYINPUT86), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n387), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n419), .A3(new_n414), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n423), .A3(new_n421), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n383), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT9), .B(G234), .Z(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G221), .B1(new_n429), .B2(G902), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n380), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n311), .A2(G952), .ZN(new_n432));
  NAND2_X1  g246(.A1(G234), .A2(G237), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT21), .B(G898), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n433), .A2(G902), .A3(G953), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n220), .A2(G143), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n203), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n220), .A2(G143), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n192), .A2(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n442), .B1(new_n445), .B2(new_n440), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n444), .A3(new_n203), .ZN(new_n447));
  XNOR2_X1  g261(.A(G116), .B(G122), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G107), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n448), .A2(new_n318), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n446), .B(new_n447), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G217), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n429), .A2(new_n453), .A3(G953), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT95), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT94), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n443), .A2(new_n444), .A3(new_n203), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n203), .B1(new_n443), .B2(new_n444), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G134), .B1(new_n215), .B2(new_n441), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT94), .A3(new_n447), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n226), .A2(KEYINPUT14), .A3(G122), .ZN(new_n463));
  OAI211_X1 g277(.A(G107), .B(new_n463), .C1(new_n449), .C2(KEYINPUT14), .ZN(new_n464));
  INV_X1    g278(.A(new_n450), .ZN(new_n465));
  AND4_X1   g279(.A1(new_n455), .A2(new_n462), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n450), .B1(new_n459), .B2(new_n461), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n455), .B1(new_n467), .B2(new_n464), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n452), .B(new_n454), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT96), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT95), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n455), .A3(new_n464), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n454), .B1(new_n475), .B2(new_n452), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n452), .B1(new_n466), .B2(new_n468), .ZN(new_n478));
  INV_X1    g292(.A(new_n454), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(KEYINPUT96), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G478), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n482), .A2(KEYINPUT97), .A3(new_n372), .A4(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G113), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(new_n315), .ZN(new_n488));
  NOR2_X1   g302(.A1(KEYINPUT88), .A2(G143), .ZN(new_n489));
  INV_X1    g303(.A(G237), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(G214), .A3(new_n490), .A4(new_n311), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT88), .B(G143), .ZN(new_n492));
  INV_X1    g306(.A(G214), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n493), .A2(G237), .A3(G953), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n210), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n311), .A3(G214), .ZN(new_n498));
  NAND2_X1  g312(.A1(KEYINPUT88), .A2(G143), .ZN(new_n499));
  OR2_X1    g313(.A1(KEYINPUT88), .A2(G143), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(G131), .A3(new_n491), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n210), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT17), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G125), .B(G140), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT16), .ZN(new_n507));
  OR3_X1    g321(.A1(new_n385), .A2(KEYINPUT16), .A3(G140), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(G146), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G146), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n502), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n505), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n506), .A2(new_n190), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n190), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n190), .B2(new_n506), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n495), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n502), .A2(new_n522), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n496), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n488), .B1(new_n515), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n502), .A2(new_n497), .ZN(new_n528));
  AOI21_X1  g342(.A(G131), .B1(new_n501), .B2(new_n491), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n504), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT90), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT72), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n507), .A2(new_n534), .A3(G146), .A4(new_n508), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n506), .B(KEYINPUT19), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n190), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n503), .A2(new_n539), .A3(new_n504), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n532), .A2(new_n536), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n488), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n525), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n527), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n527), .A2(new_n543), .A3(new_n547), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n478), .A2(new_n479), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n470), .A3(new_n469), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT97), .A3(new_n372), .A4(new_n480), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n484), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n554));
  OR3_X1    g368(.A1(new_n515), .A2(new_n526), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n515), .B2(new_n526), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n372), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT91), .B(G475), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n486), .A2(new_n549), .A3(new_n553), .A4(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n431), .A2(new_n439), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G110), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n228), .A2(G128), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(G119), .B2(new_n220), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n228), .A2(KEYINPUT23), .A3(G128), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n562), .B(new_n563), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n220), .A2(G119), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT23), .B1(new_n228), .B2(G128), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n564), .A2(new_n220), .A3(G119), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n574), .A2(new_n575), .B1(new_n228), .B2(G128), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT71), .A3(new_n562), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n533), .A3(new_n520), .A4(new_n535), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n571), .A2(new_n572), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n576), .A2(new_n562), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(new_n581), .C1(new_n510), .C2(new_n511), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n584));
  NAND2_X1  g398(.A1(G221), .A2(G234), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT22), .B1(new_n585), .B2(G953), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT22), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n587), .A2(new_n311), .A3(G221), .A4(G234), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n586), .A2(G137), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G137), .B1(new_n586), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n206), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n588), .A3(G137), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT74), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n579), .A2(new_n582), .A3(new_n594), .A4(new_n593), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n583), .A2(KEYINPUT75), .A3(new_n597), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n372), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT75), .B1(new_n583), .B2(new_n597), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n599), .B(new_n596), .C1(new_n579), .C2(new_n582), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(new_n372), .A3(new_n601), .A4(new_n604), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n453), .B1(G234), .B2(new_n372), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n609), .A2(new_n601), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n611), .A2(G902), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT77), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n309), .A2(new_n561), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT98), .B(G101), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G3));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n287), .B2(new_n372), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n287), .A2(new_n188), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT68), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n307), .A2(new_n284), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n380), .A2(new_n430), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n381), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n425), .B2(new_n426), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n439), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n627), .A2(new_n618), .A3(new_n629), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n551), .A2(new_n480), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n550), .A2(KEYINPUT33), .A3(new_n469), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(G478), .A3(new_n372), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n551), .A2(new_n480), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n483), .B1(new_n640), .B2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n549), .A2(new_n559), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT34), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  AOI21_X1  g461(.A(KEYINPUT100), .B1(new_n546), .B2(new_n548), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n545), .B2(KEYINPUT20), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n486), .A2(new_n553), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n559), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n634), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT35), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n583), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n615), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n612), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n560), .A2(new_n660), .A3(new_n439), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n627), .A3(new_n427), .A4(new_n629), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n562), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G12));
  XNOR2_X1  g479(.A(new_n434), .B(KEYINPUT102), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n438), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n648), .B2(new_n650), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n653), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n660), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n628), .A2(new_n632), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n309), .A2(new_n672), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n669), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n629), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n425), .A2(new_n426), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n630), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n679), .A2(new_n652), .A3(new_n643), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n307), .A2(KEYINPUT32), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n224), .A2(new_n237), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n281), .B1(new_n239), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n274), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(KEYINPUT103), .B2(new_n687), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n690), .B2(G902), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n289), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n660), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n192), .ZN(G45));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n696), .A2(new_n642), .A3(new_n643), .A4(new_n670), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n639), .A2(new_n641), .B1(new_n549), .B2(new_n559), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n698), .B2(new_n670), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n309), .A3(new_n673), .A4(new_n674), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NAND2_X1  g516(.A1(new_n370), .A2(new_n372), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n704), .A2(new_n373), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n430), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n644), .A2(new_n632), .A3(new_n439), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n309), .A2(new_n618), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT41), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G113), .ZN(G15));
  NOR2_X1   g525(.A1(new_n653), .A2(new_n651), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n617), .A2(new_n439), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n430), .A2(new_n631), .A3(new_n373), .A4(new_n704), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n309), .A2(new_n712), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  AOI21_X1  g530(.A(KEYINPUT32), .B1(new_n625), .B2(new_n626), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n306), .A2(G472), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n685), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n661), .B(new_n714), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  AND4_X1   g535(.A1(new_n652), .A2(new_n705), .A3(new_n430), .A4(new_n643), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n264), .A2(new_n272), .B1(new_n281), .B2(new_n300), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n189), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n623), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n723), .B1(new_n727), .B2(new_n618), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n623), .A2(new_n726), .A3(KEYINPUT105), .A4(new_n617), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n633), .B(new_n722), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR3_X1   g545(.A1(new_n623), .A2(new_n660), .A3(new_n726), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n700), .A2(new_n714), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND2_X1  g548(.A1(new_n624), .A2(new_n187), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n617), .B1(new_n308), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n377), .A2(new_n737), .A3(new_n342), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT106), .B1(new_n343), .B2(new_n348), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n376), .A2(new_n740), .A3(G469), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n373), .A2(new_n375), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n430), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n680), .A2(new_n630), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n700), .A2(new_n736), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n742), .A3(new_n430), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n617), .B(new_n746), .C1(new_n289), .C2(new_n308), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n697), .A2(new_n699), .A3(KEYINPUT42), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n745), .A2(KEYINPUT42), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n672), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND3_X1  g566(.A1(new_n642), .A2(new_n549), .A3(new_n559), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(G902), .B1(new_n273), .B2(new_n282), .ZN(new_n756));
  OAI22_X1  g570(.A1(new_n283), .A2(new_n288), .B1(new_n622), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n757), .A3(new_n673), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n376), .A2(new_n378), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n376), .A2(new_n740), .A3(KEYINPUT45), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(G469), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n375), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n375), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n373), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n430), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n677), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n758), .A2(new_n759), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n760), .A2(new_n772), .A3(new_n744), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  AND3_X1   g589(.A1(new_n770), .A2(KEYINPUT47), .A3(new_n430), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT47), .B1(new_n770), .B2(new_n430), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n309), .A2(new_n697), .A3(new_n699), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n617), .A3(new_n744), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NAND2_X1  g597(.A1(new_n755), .A2(new_n666), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n755), .A2(new_n786), .A3(new_n666), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n728), .A2(new_n729), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n682), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n381), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n788), .A2(new_n707), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT50), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n789), .B1(new_n785), .B2(new_n787), .ZN(new_n797));
  INV_X1    g611(.A(new_n795), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n707), .A3(new_n798), .A4(new_n792), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n744), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n776), .A2(new_n778), .A3(KEYINPUT112), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT112), .B1(new_n776), .B2(new_n778), .ZN(new_n803));
  INV_X1    g617(.A(new_n430), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n705), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n744), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n706), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n788), .A2(new_n732), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n692), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n618), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n435), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n642), .A2(new_n643), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n800), .A2(new_n807), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n797), .A2(new_n714), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n796), .A2(new_n799), .B1(new_n814), .B2(new_n815), .ZN(new_n821));
  INV_X1    g635(.A(new_n805), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n801), .B1(new_n780), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n788), .A2(new_n736), .A3(new_n809), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n825), .B(KEYINPUT115), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(KEYINPUT48), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n819), .A2(new_n820), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n812), .A2(new_n644), .A3(new_n813), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n617), .B1(new_n289), .B2(new_n308), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n757), .A2(new_n431), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n834), .A2(new_n561), .B1(new_n835), .B2(new_n661), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n643), .A2(new_n641), .A3(new_n639), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n439), .B(new_n383), .C1(new_n425), .C2(new_n426), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n837), .A2(new_n560), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n627), .A3(new_n618), .A4(new_n629), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n836), .A2(new_n730), .A3(new_n720), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n718), .A2(new_n735), .A3(new_n685), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT104), .B1(new_n644), .B2(new_n669), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n698), .A2(new_n696), .A3(new_n670), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n618), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT42), .B1(new_n845), .B2(new_n746), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n747), .A2(new_n748), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n709), .A2(new_n715), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n841), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n628), .B(new_n632), .C1(new_n289), .C2(new_n308), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n673), .C1(new_n672), .C2(new_n700), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n652), .A2(new_n643), .A3(new_n631), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n673), .A3(new_n669), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n692), .A2(new_n854), .A3(new_n743), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n733), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n701), .A2(new_n733), .A3(new_n855), .A4(new_n675), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n486), .A2(new_n553), .A3(new_n559), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n671), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT107), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n628), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT107), .B1(new_n671), .B2(new_n861), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n309), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n843), .A2(new_n844), .A3(new_n727), .A4(new_n743), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n660), .B(new_n808), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n751), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n868), .A2(KEYINPUT108), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT108), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n867), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n673), .A3(new_n744), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n873), .B2(new_n751), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n850), .B(new_n860), .C1(new_n870), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n619), .A2(new_n720), .A3(new_n840), .A4(new_n662), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n709), .A2(new_n715), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n749), .A2(new_n878), .A3(new_n730), .A4(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT108), .B1(new_n868), .B2(new_n869), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n871), .A3(new_n751), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(KEYINPUT53), .A3(new_n860), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n877), .A2(new_n884), .A3(KEYINPUT109), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n875), .A2(new_n876), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT53), .B1(new_n883), .B2(new_n860), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT109), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n877), .A2(new_n884), .A3(new_n885), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n833), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n895));
  OAI21_X1  g709(.A(G953), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n833), .B(new_n895), .C1(new_n887), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n432), .ZN(new_n898));
  INV_X1    g712(.A(new_n812), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n791), .A2(new_n804), .A3(new_n753), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n705), .B(KEYINPUT49), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n382), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n896), .A2(new_n898), .A3(new_n902), .ZN(G75));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n877), .A2(new_n884), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G902), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n261), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n416), .A2(new_n420), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n418), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT55), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n311), .A2(G952), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n907), .B2(new_n908), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n907), .B2(new_n908), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(G51));
  NAND2_X1  g731(.A1(new_n890), .A2(new_n892), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n374), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n375), .A2(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n370), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n906), .A2(new_n765), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n922), .B2(new_n923), .ZN(G54));
  NAND4_X1  g738(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n527), .A2(new_n543), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n914), .ZN(G60));
  NAND3_X1  g742(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n483), .A2(new_n372), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n929), .A2(new_n886), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n637), .A2(new_n638), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n890), .B2(new_n892), .ZN(new_n937));
  INV_X1    g751(.A(new_n935), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n914), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT118), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n936), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT119), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n877), .B2(new_n884), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n658), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT120), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n952), .A3(new_n658), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT121), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n914), .B1(new_n951), .B2(new_n953), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n949), .A2(new_n613), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n957), .B(new_n956), .C1(new_n954), .C2(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  AOI21_X1  g775(.A(new_n311), .B1(new_n436), .B2(G224), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n841), .A2(new_n849), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n964), .B2(new_n311), .ZN(new_n965));
  INV_X1    g779(.A(G898), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n909), .B1(new_n966), .B2(G953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  INV_X1    g782(.A(new_n853), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n772), .A2(new_n736), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n782), .A2(new_n774), .A3(new_n751), .A4(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n852), .A2(new_n733), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n749), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n972), .B1(new_n971), .B2(new_n975), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n977), .A3(new_n311), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n255), .B(new_n537), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(new_n979), .C1(new_n667), .C2(new_n311), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n694), .B2(new_n973), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n974), .B(KEYINPUT62), .C1(new_n693), .C2(new_n684), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n782), .A2(new_n774), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n678), .A2(new_n808), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n834), .A3(new_n560), .A4(new_n837), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT122), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n984), .A2(new_n990), .A3(new_n985), .A4(new_n987), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n980), .B1(new_n992), .B2(new_n979), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n994));
  AOI21_X1  g808(.A(G227), .B1(new_n979), .B2(KEYINPUT124), .ZN(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n995), .B2(new_n667), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n993), .B2(new_n994), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(G72));
  INV_X1    g813(.A(new_n914), .ZN(new_n1000));
  INV_X1    g814(.A(new_n256), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n989), .A2(new_n963), .A3(new_n991), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1001), .B(new_n263), .C1(new_n1002), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n256), .A2(new_n281), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT126), .Z(new_n1008));
  NAND3_X1  g822(.A1(new_n976), .A2(new_n977), .A3(new_n963), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1009), .A2(KEYINPUT125), .A3(new_n1004), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT125), .B1(new_n1009), .B2(new_n1004), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n291), .A2(new_n274), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n905), .A2(new_n1004), .A3(new_n1013), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n1000), .A2(new_n1006), .A3(new_n1012), .A4(new_n1014), .ZN(G57));
endmodule


