//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G250), .B1(G257), .B2(G264), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n207), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n206), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n204), .A2(G50), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(new_n217), .B2(KEYINPUT0), .ZN(new_n239));
  NAND3_X1  g0039(.A1(new_n218), .A2(new_n229), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g0040(.A(new_n240), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G358));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT66), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n225), .A2(G1698), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(new_n261), .C1(G226), .C2(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G97), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(new_n259), .A3(G274), .ZN(new_n270));
  INV_X1    g0070(.A(G238), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n259), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n264), .A2(new_n266), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n266), .B1(new_n264), .B2(new_n274), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G169), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  OR3_X1    g0079(.A1(new_n264), .A2(KEYINPUT70), .A3(new_n274), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT70), .B1(new_n264), .B2(new_n274), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(KEYINPUT13), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G179), .A3(new_n275), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(new_n284), .A3(G169), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n279), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT65), .B(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(new_n220), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n234), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT11), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n211), .A3(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n203), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n293), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(G68), .C1(G1), .C2(new_n211), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n296), .A2(new_n297), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n286), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n282), .A2(G190), .A3(new_n275), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n277), .B2(G200), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT71), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT71), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G222), .ZN(new_n317));
  INV_X1    g0117(.A(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(G223), .B1(new_n315), .B2(G77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G226), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n273), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G274), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n329), .B2(new_n269), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT9), .ZN(new_n334));
  OAI21_X1  g0134(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n287), .A2(G150), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n335), .B(new_n336), .C1(new_n290), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n293), .ZN(new_n339));
  INV_X1    g0139(.A(G50), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n210), .B2(G20), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n302), .A2(new_n341), .B1(new_n340), .B2(new_n299), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n332), .A2(new_n333), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n343), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n345), .A2(KEYINPUT9), .B1(new_n331), .B2(new_n346), .ZN(new_n347));
  OR3_X1    g0147(.A1(new_n344), .A2(new_n347), .A3(KEYINPUT10), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT10), .B1(new_n344), .B2(new_n347), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n332), .A2(G169), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n331), .A2(G179), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n351), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT68), .B1(new_n290), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n337), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n287), .B1(new_n233), .B2(G77), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n290), .A2(KEYINPUT68), .A3(new_n355), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n293), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n220), .B1(new_n210), .B2(G20), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n302), .A2(new_n362), .B1(new_n220), .B2(new_n299), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n316), .A2(G232), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT67), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n316), .A2(KEYINPUT67), .A3(G232), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n321), .A2(G238), .B1(new_n315), .B2(G107), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n259), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n270), .B1(new_n221), .B2(new_n273), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n364), .B1(new_n373), .B2(G190), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n333), .B2(new_n373), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(new_n364), .C1(G169), .C2(new_n373), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n312), .A2(new_n350), .A3(new_n354), .A4(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n337), .B1(new_n210), .B2(G20), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n302), .B1(new_n299), .B2(new_n337), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT7), .B1(new_n260), .B2(G20), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n315), .A2(new_n289), .A3(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n383), .A2(new_n385), .A3(G68), .ZN(new_n386));
  XNOR2_X1  g0186(.A(G58), .B(G68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n287), .A2(KEYINPUT72), .A3(G159), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT72), .B1(new_n287), .B2(G159), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n388), .B(KEYINPUT16), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n293), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT7), .B1(new_n233), .B2(new_n260), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n315), .A2(new_n384), .A3(new_n211), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(G68), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n391), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n389), .B1(new_n387), .B2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT16), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n382), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G223), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n318), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n326), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n313), .C2(new_n314), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n259), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n259), .A2(G232), .A3(new_n272), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n270), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(G169), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n324), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n270), .A2(new_n407), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n413), .B2(new_n376), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n400), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n400), .A2(KEYINPUT18), .A3(new_n414), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(KEYINPUT73), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n420), .A3(new_n416), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n382), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n396), .A2(new_n398), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n292), .A2(new_n234), .ZN(new_n427));
  INV_X1    g0227(.A(new_n392), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n383), .A2(new_n385), .A3(G68), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n423), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n411), .A2(new_n412), .A3(new_n346), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n333), .B1(new_n406), .B2(new_n408), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n434), .B(new_n382), .C1(new_n393), .C2(new_n399), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT74), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n426), .A2(new_n430), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT74), .A3(new_n382), .A4(new_n434), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n441), .B2(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n422), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n380), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n206), .B2(G33), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n293), .B1(new_n211), .B2(G116), .C1(new_n233), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT20), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n427), .B1(G20), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n233), .A2(new_n447), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n299), .A2(new_n451), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n298), .A2(G1), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n210), .A2(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n427), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n456), .B1(new_n460), .B2(new_n451), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n260), .A2(G264), .A3(G1698), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n260), .A2(G257), .A3(new_n318), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n315), .A2(G303), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n324), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n268), .A2(G1), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n324), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n470), .A2(new_n469), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n471), .A2(G270), .B1(new_n472), .B2(new_n329), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n463), .A2(G169), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n376), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n463), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n463), .A2(KEYINPUT21), .A3(G169), .A4(new_n474), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n461), .B1(new_n450), .B2(new_n454), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n468), .A2(new_n473), .A3(G190), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n468), .A2(new_n473), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(new_n333), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n474), .A2(G169), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n476), .B1(new_n486), .B2(new_n481), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n477), .A2(new_n463), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(new_n484), .A3(new_n488), .A4(new_n480), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(new_n318), .C1(new_n313), .C2(new_n314), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n318), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n494), .A2(new_n495), .A3(new_n446), .ZN(new_n496));
  OAI211_X1 g0296(.A(G250), .B(G1698), .C1(new_n313), .C2(new_n314), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT77), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n259), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n471), .A2(G257), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n472), .A2(new_n329), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT77), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n497), .B(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n495), .A3(new_n446), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n324), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n502), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(G179), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n394), .A2(G107), .A3(new_n395), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n208), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT75), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n208), .A2(KEYINPUT75), .A3(new_n516), .A4(new_n512), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n233), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n287), .A2(G77), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n511), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n293), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n299), .A2(new_n206), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n206), .C2(new_n460), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n510), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n492), .A2(new_n493), .B1(G33), .B2(G283), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n497), .A2(KEYINPUT77), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n497), .A2(KEYINPUT77), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n495), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n502), .B1(new_n533), .B2(new_n324), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G190), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n526), .B1(new_n521), .B2(new_n293), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n333), .C2(new_n534), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n230), .B(new_n232), .C1(new_n313), .C2(new_n314), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n203), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n263), .A2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n233), .A2(new_n542), .B1(G87), .B2(new_n208), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n230), .A2(new_n232), .A3(G33), .A4(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n541), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n289), .A2(new_n260), .A3(KEYINPUT79), .A4(G68), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n540), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n293), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n355), .A2(new_n299), .ZN(new_n549));
  INV_X1    g0349(.A(new_n460), .ZN(new_n550));
  INV_X1    g0350(.A(new_n355), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT80), .ZN(new_n554));
  OAI211_X1 g0354(.A(G244), .B(G1698), .C1(new_n313), .C2(new_n314), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n260), .A2(KEYINPUT78), .A3(G244), .A4(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G116), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n260), .A2(G238), .A3(new_n318), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n324), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n259), .B1(G250), .B2(new_n469), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n268), .A2(G1), .A3(G274), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(G179), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G169), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n561), .B2(new_n324), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT80), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n548), .A2(new_n571), .A3(new_n549), .A4(new_n552), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n554), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n550), .A2(G87), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n548), .A2(new_n549), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n562), .A2(new_n566), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n569), .A2(G190), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n529), .A2(new_n537), .A3(new_n573), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n457), .A2(G20), .A3(new_n207), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT25), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT84), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(KEYINPUT84), .A3(new_n582), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(new_n550), .B2(G107), .ZN(new_n587));
  INV_X1    g0387(.A(G87), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT22), .B1(new_n539), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n289), .A2(new_n260), .A3(new_n590), .A4(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G20), .B2(new_n559), .ZN(new_n594));
  NOR2_X1   g0394(.A1(KEYINPUT23), .A2(G107), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT82), .B1(new_n289), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n233), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n592), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT83), .B1(new_n605), .B2(new_n293), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n592), .A2(new_n600), .A3(new_n603), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n592), .B2(new_n600), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT83), .B(new_n293), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n587), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n260), .A2(G257), .A3(G1698), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n260), .A2(G250), .A3(new_n318), .ZN(new_n613));
  INV_X1    g0413(.A(G33), .ZN(new_n614));
  INV_X1    g0414(.A(G294), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n324), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT85), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n471), .A2(G264), .B1(new_n472), .B2(new_n329), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n616), .A2(new_n620), .A3(new_n324), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n619), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n622), .A2(G169), .B1(new_n624), .B2(G179), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n611), .A2(new_n626), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n622), .A2(G190), .B1(new_n624), .B2(G200), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n628), .B(new_n587), .C1(new_n606), .C2(new_n610), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n491), .A2(new_n580), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n445), .A2(new_n630), .ZN(G372));
  OAI21_X1  g0431(.A(new_n305), .B1(new_n311), .B2(new_n378), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n442), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n417), .A2(new_n418), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n353), .B1(new_n635), .B2(new_n350), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n487), .A2(new_n480), .A3(new_n488), .ZN(new_n637));
  INV_X1    g0437(.A(new_n587), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n293), .B1(new_n607), .B2(new_n608), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT83), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n609), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n637), .B1(new_n642), .B2(new_n625), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n333), .B1(new_n507), .B2(new_n508), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n528), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n535), .A2(new_n645), .B1(new_n510), .B2(new_n528), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n643), .A2(new_n629), .A3(new_n646), .A4(new_n579), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT86), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n499), .A2(new_n376), .A3(new_n502), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n568), .B1(new_n507), .B2(new_n508), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n503), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n528), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n570), .A2(new_n553), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n579), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n648), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n536), .B1(new_n503), .B2(new_n509), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n573), .A2(new_n658), .A3(KEYINPUT26), .A4(new_n579), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n647), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n636), .B1(new_n445), .B2(new_n662), .ZN(G369));
  NAND2_X1  g0463(.A1(new_n289), .A2(new_n457), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n611), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n627), .A2(new_n670), .A3(new_n629), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n642), .A2(new_n625), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n669), .ZN(new_n674));
  INV_X1    g0474(.A(new_n669), .ZN(new_n675));
  NOR4_X1   g0475(.A1(new_n642), .A2(KEYINPUT87), .A3(new_n625), .A4(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n675), .A2(new_n481), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n491), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n487), .A2(new_n480), .A3(new_n488), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n627), .A2(new_n669), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n675), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n677), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(G399));
  NOR2_X1   g0492(.A1(new_n215), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n237), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT88), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n588), .A2(new_n206), .A3(new_n207), .A4(new_n451), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n693), .A2(new_n696), .A3(new_n210), .ZN(new_n697));
  MUX2_X1   g0497(.A(new_n695), .B(KEYINPUT88), .S(new_n697), .Z(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  INV_X1    g0499(.A(KEYINPUT89), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n471), .A2(G264), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n617), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n576), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n569), .A2(KEYINPUT89), .A3(new_n617), .A4(new_n701), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n477), .A3(new_n534), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n507), .A2(new_n508), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n708), .A2(new_n376), .A3(new_n474), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(KEYINPUT30), .A3(new_n703), .A4(new_n704), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n624), .A2(new_n483), .A3(G179), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n708), .A3(new_n576), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n669), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n716), .B(new_n717), .C1(new_n630), .C2(new_n669), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n661), .A2(new_n720), .A3(new_n675), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n536), .B1(new_n510), .B2(new_n649), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n579), .A3(new_n655), .A4(new_n653), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT26), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n573), .A2(new_n658), .A3(new_n648), .A4(new_n579), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n647), .A2(new_n655), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n726), .A2(new_n675), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n719), .B(new_n721), .C1(new_n727), .C2(new_n720), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n699), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(new_n693), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n233), .A2(new_n298), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(G1), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n234), .B1(G20), .B2(new_n568), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n215), .A2(new_n260), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n268), .B2(new_n694), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n256), .B2(new_n268), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n214), .A2(new_n260), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT90), .Z(new_n746));
  AOI22_X1  g0546(.A1(new_n746), .A2(G355), .B1(new_n451), .B2(new_n215), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n740), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n376), .A2(new_n333), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n233), .A2(G190), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n233), .B1(new_n346), .B2(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(G50), .B1(G97), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n289), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n376), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n233), .A2(G190), .A3(new_n757), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G77), .B1(G58), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n756), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(G179), .A3(new_n333), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT91), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT91), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n755), .B(new_n762), .C1(new_n767), .C2(new_n207), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n763), .A2(new_n753), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n756), .A2(new_n749), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G68), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT32), .B1(new_n770), .B2(new_n771), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n211), .A2(new_n346), .A3(new_n333), .A4(G179), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n315), .B1(new_n776), .B2(G87), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n772), .A2(new_n774), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n750), .B(KEYINPUT92), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G326), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n767), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n776), .B(KEYINPUT93), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G303), .B1(new_n769), .B2(G329), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n761), .A2(G322), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n260), .B1(new_n759), .B2(G311), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n773), .A2(new_n788), .B1(G294), .B2(new_n754), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n768), .A2(new_n778), .B1(new_n783), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n734), .B(new_n748), .C1(new_n791), .C2(new_n738), .ZN(new_n792));
  INV_X1    g0592(.A(new_n737), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n684), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT94), .Z(new_n795));
  INV_X1    g0595(.A(G330), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n681), .A2(new_n796), .A3(new_n683), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n797), .A2(new_n685), .A3(new_n734), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  AND2_X1   g0600(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n767), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G283), .A2(new_n804), .B1(new_n805), .B2(G87), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n770), .A2(new_n807), .B1(new_n615), .B2(new_n760), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G107), .B2(new_n784), .ZN(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n758), .A2(new_n451), .B1(new_n810), .B2(new_n750), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n260), .B(new_n811), .C1(G97), .C2(new_n754), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n806), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n773), .A2(G150), .B1(G137), .B2(new_n751), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT97), .B(G143), .Z(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n771), .B2(new_n758), .C1(new_n760), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n805), .A2(G68), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n315), .B1(new_n754), .B2(G58), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n784), .A2(G50), .B1(new_n769), .B2(G132), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n813), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n738), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n738), .A2(new_n735), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT95), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n734), .B1(new_n828), .B2(new_n220), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n364), .A2(new_n669), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n375), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n378), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n378), .A2(new_n669), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n825), .B(new_n829), .C1(new_n836), .C2(new_n736), .ZN(new_n837));
  INV_X1    g0637(.A(new_n734), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n835), .B1(new_n662), .B2(new_n669), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n375), .A2(new_n378), .A3(new_n675), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n629), .A2(new_n646), .A3(new_n579), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n682), .B1(new_n611), .B2(new_n626), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n655), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n659), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n648), .B2(new_n723), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n838), .B1(new_n847), .B2(new_n719), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n847), .A2(new_n719), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n837), .B1(new_n849), .B2(new_n850), .ZN(G384));
  NOR2_X1   g0651(.A1(new_n732), .A2(new_n210), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n304), .B(new_n669), .C1(new_n311), .C2(new_n286), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n304), .A2(new_n669), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n305), .B(new_n854), .C1(new_n310), .C2(new_n309), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n718), .A2(new_n856), .A3(new_n836), .ZN(new_n857));
  INV_X1    g0657(.A(new_n415), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n431), .A2(new_n667), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n859), .A2(new_n438), .A3(new_n440), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT16), .B1(new_n429), .B2(new_n398), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n382), .B1(new_n393), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n667), .B(new_n409), .C1(new_n413), .C2(new_n376), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n438), .A2(new_n440), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n867), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT101), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n862), .B(KEYINPUT102), .C1(new_n868), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n667), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n422), .B2(new_n442), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n880), .B(new_n877), .C1(new_n872), .C2(new_n873), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n857), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n885));
  INV_X1    g0685(.A(new_n442), .ZN(new_n886));
  INV_X1    g0686(.A(new_n634), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n860), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n415), .A2(new_n436), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n889), .B2(new_n860), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n862), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  AND4_X1   g0694(.A1(KEYINPUT40), .A2(new_n718), .A3(new_n856), .A4(new_n836), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n444), .A2(new_n718), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n796), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT101), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n867), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT102), .B1(new_n905), .B2(new_n862), .ZN(new_n906));
  INV_X1    g0706(.A(new_n873), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n878), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n880), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n881), .B2(new_n892), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n305), .A2(new_n669), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n885), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n846), .A2(new_n834), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT100), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n846), .A2(new_n918), .A3(new_n834), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(new_n920), .A3(new_n856), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n887), .A2(new_n667), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n721), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n720), .B1(new_n726), .B2(new_n675), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n444), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n636), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n923), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n852), .B1(new_n900), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n900), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n236), .A2(new_n451), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT98), .Z(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT35), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT36), .Z(new_n938));
  AOI211_X1 g0738(.A(new_n220), .B(new_n237), .C1(G58), .C2(G68), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n939), .A2(KEYINPUT99), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n939), .A2(KEYINPUT99), .B1(new_n203), .B2(new_n201), .ZN(new_n941));
  OAI211_X1 g0741(.A(G1), .B(new_n298), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n930), .A2(new_n938), .A3(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n741), .A2(new_n248), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n740), .B1(new_n215), .B2(new_n551), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n734), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n575), .A2(new_n675), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n656), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n553), .A3(new_n570), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n805), .A2(G77), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n951), .B1(new_n771), .B2(new_n803), .C1(new_n779), .C2(new_n815), .ZN(new_n952));
  INV_X1    g0752(.A(G150), .ZN(new_n953));
  INV_X1    g0753(.A(new_n776), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n260), .B1(new_n760), .B2(new_n953), .C1(new_n954), .C2(new_n202), .ZN(new_n955));
  INV_X1    g0755(.A(new_n754), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n203), .ZN(new_n957));
  INV_X1    g0757(.A(G137), .ZN(new_n958));
  INV_X1    g0758(.A(new_n201), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n770), .A2(new_n958), .B1(new_n959), .B2(new_n758), .ZN(new_n960));
  NOR4_X1   g0760(.A1(new_n952), .A2(new_n955), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n767), .A2(new_n206), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n803), .A2(new_n615), .B1(new_n807), .B2(new_n779), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n954), .A2(new_n451), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n315), .B1(new_n810), .B2(new_n760), .C1(new_n964), .C2(KEYINPUT46), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n769), .A2(G317), .B1(G107), .B2(new_n754), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n784), .A2(KEYINPUT46), .A3(G116), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n782), .C2(new_n758), .ZN(new_n968));
  NOR4_X1   g0768(.A1(new_n962), .A2(new_n963), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  INV_X1    g0771(.A(new_n738), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n946), .B1(new_n793), .B2(new_n950), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT106), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n693), .B(KEYINPUT41), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n677), .A2(new_n690), .ZN(new_n976));
  INV_X1    g0776(.A(new_n688), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n646), .B1(new_n536), .B2(new_n675), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n722), .A2(new_n653), .A3(new_n669), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n691), .B2(new_n980), .ZN(new_n987));
  INV_X1    g0787(.A(new_n980), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n611), .A2(new_n626), .A3(new_n669), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT87), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n673), .A2(new_n672), .A3(new_n669), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n689), .B1(new_n992), .B2(new_n671), .ZN(new_n993));
  OAI211_X1 g0793(.A(KEYINPUT44), .B(new_n988), .C1(new_n993), .C2(new_n688), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n985), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n686), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n992), .A2(new_n671), .A3(new_n689), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n685), .B1(new_n999), .B2(new_n993), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n976), .A2(G330), .A3(new_n998), .A4(new_n684), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n1002), .A2(new_n728), .A3(KEYINPUT104), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n985), .A2(new_n687), .A3(new_n995), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT104), .B1(new_n1002), .B2(new_n728), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n997), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n975), .B1(new_n1006), .B2(new_n729), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT105), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(KEYINPUT105), .B(new_n975), .C1(new_n1006), .C2(new_n729), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n733), .A2(G1), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n980), .A2(new_n673), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n669), .B1(new_n1015), .B2(new_n529), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n993), .A2(new_n980), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(KEYINPUT42), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(KEYINPUT42), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT103), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n950), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n687), .A2(new_n988), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1019), .B(new_n1020), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1030), .A2(new_n1025), .A3(new_n1024), .A4(new_n1018), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n974), .B1(new_n1014), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT107), .ZN(G387));
  AND2_X1   g0836(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n678), .A2(new_n737), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n337), .A2(G50), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT109), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT108), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n268), .B1(new_n203), .B2(new_n220), .C1(new_n696), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n696), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1040), .A2(KEYINPUT50), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n741), .B1(new_n245), .B2(new_n268), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n746), .A2(new_n696), .B1(new_n207), .B2(new_n215), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(KEYINPUT110), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n739), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT110), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n838), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n754), .A2(new_n551), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n340), .B2(new_n760), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT111), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n773), .A2(new_n357), .B1(G159), .B2(new_n751), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n953), .B2(new_n770), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n260), .B1(new_n954), .B2(new_n220), .C1(new_n758), .C2(new_n203), .ZN(new_n1058));
  OR4_X1    g0858(.A1(new_n962), .A2(new_n1055), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n780), .A2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n759), .A2(G303), .B1(G317), .B2(new_n761), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n803), .C2(new_n807), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n956), .A2(new_n782), .B1(new_n954), .B2(new_n615), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n260), .B1(new_n769), .B2(G326), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n451), .C2(new_n767), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1059), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1052), .B1(new_n1072), .B2(new_n738), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1037), .A2(new_n1012), .B1(new_n1038), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1002), .A2(new_n728), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n693), .B1(new_n1002), .B2(new_n728), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1037), .A2(new_n729), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n693), .A3(new_n1075), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(KEYINPUT113), .A3(new_n1074), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(G393));
  AND3_X1   g0884(.A1(new_n985), .A2(new_n995), .A3(new_n687), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n687), .B1(new_n985), .B2(new_n995), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1006), .A2(new_n1087), .A3(new_n693), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT114), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n997), .A2(new_n1090), .A3(new_n1004), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1091), .A3(new_n1012), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n980), .A2(new_n793), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT115), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n253), .A2(new_n742), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n739), .B1(new_n206), .B2(new_n214), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n838), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n260), .B1(new_n954), .B2(new_n203), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n770), .A2(new_n815), .B1(new_n337), .B2(new_n758), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G77), .C2(new_n754), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n588), .B2(new_n767), .C1(new_n803), .C2(new_n959), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n953), .A2(new_n750), .B1(new_n760), .B2(new_n771), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  OAI21_X1  g0903(.A(new_n315), .B1(new_n954), .B2(new_n782), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n769), .B2(G322), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n759), .A2(G294), .B1(G116), .B2(new_n754), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n767), .C2(new_n207), .ZN(new_n1107));
  INV_X1    g0907(.A(G317), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n807), .A2(new_n760), .B1(new_n750), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n804), .A2(G303), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1101), .A2(new_n1103), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1097), .B1(new_n1114), .B2(new_n738), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1094), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1092), .A2(KEYINPUT117), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT117), .B1(new_n1092), .B2(new_n1116), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1088), .B1(new_n1118), .B2(new_n1119), .ZN(G390));
  NAND4_X1  g0920(.A1(new_n718), .A2(new_n856), .A3(G330), .A4(new_n836), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(KEYINPUT100), .B(new_n833), .C1(new_n661), .C2(new_n840), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n918), .B1(new_n846), .B2(new_n834), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n856), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n913), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n912), .A2(new_n910), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n726), .A2(new_n675), .A3(new_n832), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n856), .B1(new_n1129), .B2(new_n833), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n1126), .A3(new_n894), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1122), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT39), .B1(new_n885), .B2(new_n893), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n879), .A2(new_n881), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(KEYINPUT39), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n913), .B1(new_n920), .B2(new_n856), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1121), .B(new_n1131), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n444), .A2(G330), .A3(new_n718), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n926), .A2(new_n1139), .A3(new_n636), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n718), .A2(G330), .A3(new_n836), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n856), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1121), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n920), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1143), .A2(new_n834), .A3(new_n1121), .A4(new_n1128), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1140), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1133), .A2(new_n1138), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n693), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT118), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT118), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1151), .A3(new_n693), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1140), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1133), .A2(new_n1138), .A3(new_n1012), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n838), .B1(new_n827), .B2(new_n357), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G137), .A2(new_n804), .B1(new_n805), .B2(new_n201), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n769), .A2(G125), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G128), .A2(new_n751), .B1(new_n761), .B2(G132), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n758), .A2(new_n1164), .B1(new_n956), .B2(new_n771), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n954), .A2(new_n953), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT53), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n260), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1165), .B(new_n1168), .C1(new_n1167), .C2(new_n1166), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n761), .A2(G116), .B1(G77), .B2(new_n754), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT119), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n820), .B(new_n1172), .C1(new_n207), .C2(new_n803), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n260), .B1(new_n784), .B2(G87), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n769), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n206), .C2(new_n758), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1170), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1160), .B1(new_n1177), .B2(new_n738), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1136), .B2(new_n736), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1159), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1158), .A2(new_n1181), .ZN(G378));
  NOR2_X1   g0982(.A1(new_n260), .A2(G41), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G50), .B(new_n1183), .C1(new_n614), .C2(new_n267), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n805), .A2(G58), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n758), .A2(new_n355), .B1(new_n207), .B2(new_n760), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G97), .B2(new_n773), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n954), .B2(new_n220), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n957), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n769), .A2(G283), .B1(G116), .B2(new_n751), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n759), .A2(G137), .B1(G150), .B2(new_n754), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1164), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n773), .A2(G132), .B1(new_n776), .B2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G125), .A2(new_n751), .B1(new_n761), .B2(G128), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n771), .C2(new_n767), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1193), .B1(new_n1192), .B2(new_n1191), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n738), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n734), .B1(new_n959), .B2(new_n826), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n350), .A2(new_n354), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n345), .A2(new_n667), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1206), .B(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1204), .B(new_n1205), .C1(new_n1211), .C2(new_n736), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n914), .A2(new_n921), .A3(new_n922), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n796), .B1(new_n894), .B2(new_n895), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n884), .A2(new_n1210), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1210), .B1(new_n884), .B2(new_n1215), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1215), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT40), .B1(new_n915), .B2(new_n857), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1211), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n884), .A2(new_n1210), .A3(new_n1215), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n923), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1213), .B1(new_n1224), .B2(new_n1012), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1218), .A2(new_n1223), .A3(KEYINPUT121), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT121), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1221), .A2(new_n923), .A3(new_n1222), .A4(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(KEYINPUT57), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1148), .A2(new_n1155), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n693), .B1(new_n1232), .B2(KEYINPUT57), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1225), .B1(new_n1231), .B2(new_n1233), .ZN(G375));
  NAND2_X1  g1034(.A1(new_n1154), .A2(new_n1012), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n838), .B1(new_n827), .B2(G68), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n769), .A2(G128), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n953), .B2(new_n758), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G132), .B2(new_n751), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n260), .B1(new_n760), .B2(new_n958), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n956), .A2(new_n340), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(G159), .C2(new_n784), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n804), .A2(new_n1195), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1185), .A2(new_n1239), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n951), .A2(new_n315), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT123), .Z(new_n1246));
  NAND2_X1  g1046(.A1(new_n761), .A2(G283), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n784), .A2(G97), .B1(new_n769), .B2(G303), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1053), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n759), .A2(G107), .B1(G294), .B2(new_n751), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n803), .B2(new_n451), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1244), .B1(new_n1249), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1236), .B1(new_n1253), .B2(new_n738), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n736), .B2(new_n856), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1235), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n975), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1145), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1156), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G381));
  NAND3_X1  g1061(.A1(new_n1080), .A2(new_n799), .A3(new_n1083), .ZN(new_n1262));
  OR4_X1    g1062(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1262), .ZN(new_n1263));
  OR4_X1    g1063(.A1(G387), .A2(new_n1263), .A3(G378), .A4(G375), .ZN(G407));
  AOI22_X1  g1064(.A1(new_n1149), .A2(KEYINPUT118), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1180), .B1(new_n1265), .B2(new_n1152), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n668), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G375), .C2(new_n1267), .ZN(G409));
  AOI21_X1  g1068(.A(new_n799), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT107), .B1(new_n1270), .B2(new_n1262), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G390), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1262), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(new_n1269), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1092), .A2(new_n1116), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT117), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1117), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1274), .B1(new_n1278), .B2(new_n1088), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1035), .B1(new_n1272), .B2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1278), .B(new_n1088), .C1(new_n1274), .C2(KEYINPUT107), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1270), .A2(new_n1262), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G390), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1013), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1034), .B1(new_n1284), .B2(new_n1010), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n974), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1281), .A2(new_n1283), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1280), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n668), .A2(G213), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(G375), .A2(new_n1266), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT124), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1227), .A2(KEYINPUT124), .A3(new_n1229), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1012), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1213), .B1(new_n1232), .B2(new_n1258), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G378), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1290), .B1(new_n1291), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1259), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1156), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1301), .B2(new_n1156), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n693), .B1(new_n1259), .B2(new_n1300), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1299), .B1(new_n1306), .B2(new_n1256), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1257), .C1(new_n1308), .C2(new_n1303), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1290), .A2(KEYINPUT126), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1290), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1307), .A2(new_n1309), .A3(new_n1313), .A4(new_n1310), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1317), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1290), .B(new_n1319), .C1(new_n1291), .C2(new_n1297), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT62), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(KEYINPUT62), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1289), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1307), .A2(new_n1309), .A3(KEYINPUT63), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1290), .B(new_n1325), .C1(new_n1291), .C2(new_n1297), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1281), .A2(new_n1283), .A3(new_n1287), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1287), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1294), .A2(new_n1012), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1296), .B1(new_n1332), .B2(new_n1292), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1266), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1226), .A2(new_n1224), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT57), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n693), .A3(new_n1230), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(G378), .A2(new_n1338), .A3(new_n1225), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1312), .B1(new_n1334), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1331), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1330), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1320), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1289), .B1(new_n1340), .B2(new_n1325), .ZN(new_n1347));
  AND4_X1   g1147(.A1(KEYINPUT127), .A2(new_n1318), .A3(new_n1347), .A4(new_n1345), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1324), .B1(new_n1346), .B2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1266), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1339), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1319), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1351), .B(new_n1352), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1329), .ZN(G402));
endmodule


