//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n461), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n465), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OAI21_X1  g056(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(G126), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n466), .B2(new_n467), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(new_n485), .C1(new_n466), .C2(new_n467), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n462), .A2(new_n493), .A3(G138), .A4(new_n461), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT70), .B(G651), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(G651), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(KEYINPUT6), .C1(KEYINPUT70), .C2(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT71), .A3(G651), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n506), .A2(new_n500), .A3(G88), .A4(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n506), .A2(G50), .A3(G543), .A4(new_n508), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT72), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n500), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n498), .A2(KEYINPUT73), .A3(new_n499), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  AND3_X1   g095(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT6), .B1(KEYINPUT70), .B2(G651), .ZN(new_n522));
  OAI211_X1 g097(.A(G543), .B(new_n508), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n506), .A2(new_n500), .A3(new_n508), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(G168));
  AND2_X1   g107(.A1(new_n516), .A2(new_n517), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G64), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n503), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n527), .A2(new_n537), .B1(new_n538), .B2(new_n523), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n518), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n502), .B1(new_n543), .B2(KEYINPUT75), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n527), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT76), .B(G81), .ZN(new_n548));
  INV_X1    g123(.A(new_n523), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(G43), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n546), .A2(G860), .A3(new_n550), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n498), .A2(new_n499), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n547), .A2(G91), .B1(new_n559), .B2(G651), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n523), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(new_n524), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(G286));
  NAND2_X1  g145(.A1(new_n549), .A2(G49), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n506), .A2(new_n500), .A3(G87), .A4(new_n508), .ZN(new_n572));
  AOI21_X1  g147(.A(G74), .B1(new_n516), .B2(new_n517), .ZN(new_n573));
  INV_X1    g148(.A(G651), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(G288));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n498), .B2(new_n499), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n502), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n506), .A2(new_n500), .A3(G86), .A4(new_n508), .ZN(new_n580));
  INV_X1    g155(.A(G48), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n523), .ZN(G305));
  NAND2_X1  g157(.A1(new_n533), .A2(G60), .ZN(new_n583));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n503), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n527), .A2(new_n586), .B1(new_n587), .B2(new_n523), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  OR3_X1    g166(.A1(G171), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT77), .B1(G171), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n557), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n549), .B2(G54), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n527), .A2(KEYINPUT10), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT10), .B1(new_n527), .B2(new_n598), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n592), .B(new_n593), .C1(G868), .C2(new_n601), .ZN(G284));
  OAI211_X1 g177(.A(new_n592), .B(new_n593), .C1(G868), .C2(new_n601), .ZN(G321));
  NAND2_X1  g178(.A1(G299), .A2(new_n591), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n591), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n591), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n601), .B1(new_n607), .B2(G860), .ZN(G148));
  OAI21_X1  g183(.A(new_n550), .B1(new_n544), .B2(new_n545), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n607), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT78), .ZN(new_n611));
  MUX2_X1   g186(.A(new_n609), .B(new_n611), .S(G868), .Z(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n474), .A2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n476), .A2(G135), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n461), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT79), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT80), .B(G2096), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n462), .A2(new_n469), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2430), .Z(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n633), .B(new_n637), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(G14), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n639), .ZN(G401));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n659), .A2(KEYINPUT20), .A3(new_n662), .ZN(new_n668));
  OAI221_X1 g243(.A(new_n664), .B1(new_n662), .B2(new_n663), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT84), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(G6), .B(G305), .S(G16), .Z(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  NAND2_X1  g266(.A1(G166), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G16), .B2(G22), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n687), .B(new_n690), .C1(new_n691), .C2(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n694), .A2(KEYINPUT34), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n474), .A2(G119), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n476), .A2(G131), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n461), .A2(G107), .ZN(new_n699));
  OAI21_X1  g274(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n681), .A2(G24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n589), .B2(new_n681), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT85), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n696), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT34), .B1(new_n694), .B2(new_n695), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  MUX2_X1   g293(.A(G19), .B(new_n609), .S(G16), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT89), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1341), .Z(new_n721));
  NOR2_X1   g296(.A1(G5), .A2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT92), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G301), .B2(new_n681), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n681), .A2(G20), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT23), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G299), .B2(G16), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1956), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n681), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n681), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1966), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n727), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT25), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n462), .A2(G127), .ZN(new_n740));
  NAND2_X1  g315(.A1(G115), .A2(G2104), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n461), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n739), .B(new_n742), .C1(G139), .C2(new_n476), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(new_n736), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G2072), .Z(new_n745));
  AND2_X1   g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n736), .B1(KEYINPUT24), .B2(G34), .ZN(new_n747));
  OAI22_X1  g322(.A1(G160), .A2(new_n736), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G2084), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  AND2_X1   g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  INV_X1    g326(.A(G28), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(KEYINPUT30), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n736), .B1(new_n754), .B2(G28), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n749), .B1(new_n750), .B2(new_n751), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n619), .A2(new_n736), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n748), .A2(G2084), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n474), .A2(G128), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n476), .A2(G140), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n461), .A2(G116), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n736), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n745), .A2(new_n759), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(G29), .A2(G32), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n773));
  AND3_X1   g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(G105), .B2(new_n469), .ZN(new_n777));
  AOI22_X1  g352(.A1(G129), .A2(new_n474), .B1(new_n476), .B2(G141), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT91), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n736), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n736), .A2(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n736), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n681), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n601), .B2(new_n681), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n771), .A2(new_n783), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n781), .A2(new_n782), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n736), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n736), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT29), .Z(new_n794));
  INV_X1    g369(.A(G2090), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n794), .A2(new_n795), .B1(new_n724), .B2(new_n725), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n791), .B(new_n796), .C1(new_n795), .C2(new_n794), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G1966), .B2(new_n733), .ZN(new_n798));
  AND4_X1   g373(.A1(new_n721), .A2(new_n735), .A3(new_n790), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n717), .A2(new_n718), .A3(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  NAND2_X1  g376(.A1(new_n533), .A2(G67), .ZN(new_n802));
  NAND2_X1  g377(.A1(G80), .A2(G543), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n503), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT94), .B(G93), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n547), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n549), .A2(G55), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G860), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n546), .A2(new_n809), .A3(new_n814), .A4(new_n550), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n802), .A2(new_n803), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(new_n502), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n817), .A2(new_n814), .A3(new_n807), .A4(new_n806), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT95), .B1(new_n804), .B2(new_n808), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n609), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT38), .Z(new_n822));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n607), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT96), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n810), .B1(new_n826), .B2(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n813), .B1(new_n828), .B2(new_n829), .ZN(G145));
  XNOR2_X1  g405(.A(new_n764), .B(new_n496), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n701), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n474), .A2(G130), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n476), .A2(G142), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n461), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n623), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n743), .A2(new_n779), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n780), .B2(new_n743), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n619), .B(G160), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G162), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT98), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(G37), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n842), .A2(new_n844), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT99), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g426(.A1(new_n601), .A2(G299), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n823), .A2(new_n564), .A3(new_n560), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n855), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n858), .A2(KEYINPUT102), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n854), .A2(new_n855), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n821), .B(new_n611), .ZN(new_n866));
  MUX2_X1   g441(.A(new_n865), .B(new_n859), .S(new_n866), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n589), .B(G303), .ZN(new_n868));
  XNOR2_X1  g443(.A(G288), .B(G305), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT103), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT42), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G868), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(G868), .B2(new_n809), .ZN(G295));
  OAI21_X1  g450(.A(new_n874), .B1(G868), .B2(new_n809), .ZN(G331));
  XNOR2_X1  g451(.A(G171), .B(G168), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n821), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  XNOR2_X1  g454(.A(G171), .B(G286), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n815), .A3(new_n820), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n880), .A2(KEYINPUT104), .A3(new_n815), .A4(new_n820), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n859), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT105), .ZN(new_n886));
  INV_X1    g461(.A(new_n870), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n865), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n862), .B1(new_n882), .B2(new_n883), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n886), .A2(new_n887), .A3(new_n889), .A4(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI211_X1 g470(.A(KEYINPUT105), .B(new_n862), .C1(new_n882), .C2(new_n883), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n861), .A2(new_n864), .B1(new_n881), .B2(new_n878), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n887), .A4(new_n886), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n854), .A2(new_n857), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT41), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(KEYINPUT41), .B2(new_n859), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n884), .A2(new_n903), .B1(new_n862), .B2(new_n888), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n904), .B2(new_n870), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n887), .B1(new_n898), .B2(new_n886), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(G37), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n890), .A2(new_n891), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n913), .A2(new_n896), .A3(new_n897), .ZN(new_n914));
  OAI211_X1 g489(.A(KEYINPUT106), .B(new_n912), .C1(new_n914), .C2(new_n887), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n911), .A2(new_n900), .A3(KEYINPUT43), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n911), .A2(new_n900), .A3(new_n907), .A4(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n912), .B1(new_n914), .B2(new_n887), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n920), .A2(new_n909), .B1(new_n895), .B2(new_n899), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n907), .A4(new_n915), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n917), .B1(new_n925), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n496), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G125), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n473), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n464), .ZN(new_n933));
  OAI21_X1  g508(.A(G2105), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n471), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(G40), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n939), .A2(KEYINPUT46), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(KEYINPUT46), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n764), .B(new_n769), .ZN(new_n942));
  INV_X1    g517(.A(new_n779), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n940), .A2(new_n941), .B1(new_n937), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT47), .Z(new_n946));
  NOR2_X1   g521(.A1(new_n939), .A2(new_n780), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT109), .Z(new_n948));
  OAI21_X1  g523(.A(new_n942), .B1(new_n943), .B2(new_n938), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n701), .A2(new_n703), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n701), .A2(new_n703), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n937), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(G290), .A2(G1986), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n937), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT48), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n946), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n952), .B(KEYINPUT125), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n950), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(G2067), .B2(new_n764), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n937), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT123), .ZN(new_n964));
  INV_X1    g539(.A(G40), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n465), .A2(new_n965), .A3(new_n471), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n490), .B2(new_n495), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n495), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(G2084), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n936), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n972));
  AOI21_X1  g547(.A(G1966), .B1(new_n930), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G8), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  NOR2_X1   g550(.A1(G168), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT51), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G286), .A2(G8), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n979), .B2(KEYINPUT120), .ZN(new_n982));
  INV_X1    g557(.A(G1966), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n966), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n928), .A2(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(G2084), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n967), .A2(new_n968), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n966), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(G8), .B(new_n982), .C1(new_n992), .C2(G286), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n980), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n979), .B1(new_n987), .B2(new_n991), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT121), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(new_n995), .C1(new_n980), .C2(new_n993), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n997), .A2(new_n999), .A3(KEYINPUT62), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n928), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n972), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n691), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n969), .A2(new_n970), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n795), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1012), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT111), .A3(new_n1010), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1008), .A2(G8), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n967), .A2(new_n966), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G288), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n975), .B1(new_n967), .B2(new_n966), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(new_n1023), .C1(new_n1019), .C2(G288), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n549), .A2(G48), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1027), .A2(new_n670), .A3(new_n580), .A4(new_n579), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n1023), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1031), .A2(new_n1035), .A3(new_n1032), .A4(new_n1023), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1025), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1004), .A2(new_n691), .B1(new_n1006), .B2(new_n795), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(new_n975), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1016), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT117), .B1(new_n969), .B2(new_n970), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n988), .A2(new_n1043), .A3(new_n966), .A4(new_n990), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1044), .A3(new_n725), .ZN(new_n1045));
  INV_X1    g620(.A(G2078), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1001), .A2(new_n1003), .A3(new_n972), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n930), .A2(new_n972), .A3(KEYINPUT53), .A4(new_n1046), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1041), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n964), .B1(new_n1000), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n994), .A2(new_n996), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n998), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n994), .A2(KEYINPUT121), .A3(new_n996), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT123), .B(new_n1053), .C1(new_n1059), .C2(KEYINPUT62), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1039), .A2(new_n975), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1037), .A2(new_n1063), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n683), .A2(new_n1019), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1028), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n974), .A2(G286), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1016), .A2(new_n1040), .A3(new_n1037), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1072), .A2(KEYINPUT114), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1072), .B2(KEYINPUT114), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n564), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G299), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n560), .B(new_n564), .C1(new_n1077), .C2(KEYINPUT57), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1001), .A2(new_n1003), .A3(new_n972), .A4(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT115), .B(G1956), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n969), .B2(new_n970), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1081), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1042), .A2(new_n1044), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n967), .A2(new_n966), .A3(new_n769), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n823), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1081), .B1(new_n1086), .B2(new_n1083), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1088), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1087), .B2(new_n1097), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT119), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1102), .B(new_n1099), .C1(new_n1087), .C2(new_n1097), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1001), .A2(new_n1003), .A3(new_n972), .A4(new_n938), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1017), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n609), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT59), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1087), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT60), .B(new_n823), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1104), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT60), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT118), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1093), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1114), .A2(new_n1118), .A3(new_n823), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1098), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n997), .A2(new_n999), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n471), .A2(KEYINPUT122), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n471), .A2(KEYINPUT122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1046), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1124));
  NOR4_X1   g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n465), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n930), .A2(new_n984), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1045), .A2(new_n1049), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(KEYINPUT54), .C1(G171), .C2(new_n1051), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1016), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1045), .A2(new_n1049), .A3(G301), .A4(new_n1126), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1052), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1129), .B(new_n1130), .C1(new_n1132), .C2(KEYINPUT54), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1121), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1076), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1062), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n589), .A2(new_n672), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n937), .B1(new_n955), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n950), .A2(new_n1138), .A3(new_n953), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT124), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1142), .B(new_n1139), .C1(new_n1062), .C2(new_n1135), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n963), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT127), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1146), .B(new_n963), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g723(.A(G319), .ZN(new_n1150));
  NOR3_X1   g724(.A1(G401), .A2(new_n1150), .A3(G227), .ZN(new_n1151));
  OAI21_X1  g725(.A(new_n1151), .B1(new_n678), .B2(new_n679), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n849), .B2(new_n847), .ZN(new_n1153));
  AND2_X1   g727(.A1(new_n908), .A2(new_n916), .ZN(new_n1154));
  AND2_X1   g728(.A1(new_n1153), .A2(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(G225));
endmodule


