

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732;

  INV_X1 U370 ( .A(KEYINPUT46), .ZN(n348) );
  NOR2_X1 U371 ( .A1(n536), .A2(n547), .ZN(n540) );
  XNOR2_X1 U372 ( .A(n460), .B(n428), .ZN(n717) );
  INV_X1 U373 ( .A(G125), .ZN(n403) );
  XNOR2_X2 U374 ( .A(n500), .B(n360), .ZN(n505) );
  NAND2_X2 U375 ( .A1(n469), .A2(G214), .ZN(n630) );
  XNOR2_X2 U376 ( .A(n653), .B(n652), .ZN(n654) );
  AND2_X2 U377 ( .A1(n679), .A2(n582), .ZN(n546) );
  NOR2_X1 U378 ( .A1(n577), .A2(n347), .ZN(n580) );
  XNOR2_X2 U379 ( .A(n556), .B(n348), .ZN(n347) );
  OR2_X2 U380 ( .A1(n698), .A2(G902), .ZN(n437) );
  XNOR2_X2 U381 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X2 U382 ( .A(KEYINPUT34), .B(KEYINPUT83), .ZN(n362) );
  XOR2_X2 U383 ( .A(KEYINPUT76), .B(KEYINPUT22), .Z(n360) );
  NOR2_X2 U384 ( .A1(n608), .A2(KEYINPUT2), .ZN(n610) );
  NOR2_X1 U385 ( .A1(n679), .A2(n581), .ZN(n635) );
  INV_X1 U386 ( .A(n549), .ZN(n625) );
  INV_X1 U387 ( .A(G953), .ZN(n459) );
  XNOR2_X2 U388 ( .A(n599), .B(n598), .ZN(n686) );
  AND2_X2 U389 ( .A1(n649), .A2(n651), .ZN(n388) );
  NAND2_X2 U390 ( .A1(n356), .A2(n389), .ZN(n651) );
  XNOR2_X2 U391 ( .A(n599), .B(n598), .ZN(n373) );
  NAND2_X1 U392 ( .A1(n505), .A2(n358), .ZN(n396) );
  NOR2_X1 U393 ( .A1(n560), .A2(n475), .ZN(n378) );
  AND2_X1 U394 ( .A1(n394), .A2(n391), .ZN(n356) );
  XNOR2_X1 U395 ( .A(n479), .B(n364), .ZN(n718) );
  INV_X1 U396 ( .A(KEYINPUT19), .ZN(n354) );
  BUF_X1 U397 ( .A(n412), .Z(n351) );
  NAND2_X1 U398 ( .A1(n363), .A2(n557), .ZN(n353) );
  XNOR2_X1 U399 ( .A(n514), .B(KEYINPUT31), .ZN(n412) );
  NOR2_X1 U400 ( .A1(n376), .A2(n566), .ZN(n457) );
  NOR2_X1 U401 ( .A1(n376), .A2(n549), .ZN(n513) );
  NOR2_X1 U402 ( .A1(n519), .A2(n352), .ZN(n520) );
  BUF_X1 U403 ( .A(n619), .Z(n352) );
  XNOR2_X1 U404 ( .A(n368), .B(KEYINPUT1), .ZN(n619) );
  NOR2_X1 U405 ( .A1(n535), .A2(n474), .ZN(n475) );
  XNOR2_X1 U406 ( .A(n458), .B(G134), .ZN(n479) );
  XNOR2_X1 U407 ( .A(KEYINPUT67), .B(G101), .ZN(n446) );
  INV_X1 U408 ( .A(KEYINPUT4), .ZN(n409) );
  XOR2_X1 U409 ( .A(KEYINPUT91), .B(KEYINPUT0), .Z(n361) );
  NAND2_X1 U410 ( .A1(n541), .A2(n630), .ZN(n366) );
  NAND2_X1 U411 ( .A1(n525), .A2(n526), .ZN(n371) );
  XNOR2_X1 U412 ( .A(n524), .B(KEYINPUT89), .ZN(n525) );
  NAND2_X1 U413 ( .A1(n510), .A2(n509), .ZN(n526) );
  NAND2_X1 U414 ( .A1(n350), .A2(n517), .ZN(n521) );
  NAND2_X1 U415 ( .A1(n410), .A2(n411), .ZN(n350) );
  XNOR2_X2 U416 ( .A(n353), .B(KEYINPUT35), .ZN(n730) );
  XNOR2_X2 U417 ( .A(n569), .B(n354), .ZN(n560) );
  XNOR2_X2 U418 ( .A(n366), .B(KEYINPUT90), .ZN(n569) );
  XNOR2_X1 U419 ( .A(n601), .B(n603), .ZN(n604) );
  AND2_X1 U420 ( .A1(n649), .A2(n651), .ZN(n355) );
  NAND2_X2 U421 ( .A1(n511), .A2(n499), .ZN(n500) );
  AND2_X1 U422 ( .A1(n568), .A2(n679), .ZN(n583) );
  XNOR2_X1 U423 ( .A(n457), .B(n370), .ZN(n407) );
  INV_X1 U424 ( .A(KEYINPUT33), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n435), .B(KEYINPUT25), .ZN(n436) );
  INV_X1 U426 ( .A(KEYINPUT65), .ZN(n393) );
  XNOR2_X1 U427 ( .A(KEYINPUT10), .B(G140), .ZN(n428) );
  XOR2_X1 U428 ( .A(G140), .B(KEYINPUT80), .Z(n419) );
  XNOR2_X1 U429 ( .A(n408), .B(n414), .ZN(n364) );
  XNOR2_X1 U430 ( .A(G131), .B(KEYINPUT69), .ZN(n414) );
  XNOR2_X1 U431 ( .A(n409), .B(G137), .ZN(n408) );
  AND2_X1 U432 ( .A1(n392), .A2(n615), .ZN(n391) );
  NAND2_X1 U433 ( .A1(n503), .A2(n393), .ZN(n392) );
  XNOR2_X1 U434 ( .A(n549), .B(n456), .ZN(n566) );
  NOR2_X1 U435 ( .A1(n729), .A2(n732), .ZN(n556) );
  XNOR2_X1 U436 ( .A(G143), .B(G104), .ZN(n490) );
  XOR2_X1 U437 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n491) );
  XNOR2_X1 U438 ( .A(G113), .B(G131), .ZN(n489) );
  XNOR2_X1 U439 ( .A(n384), .B(KEYINPUT81), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n718), .B(G146), .ZN(n452) );
  INV_X1 U441 ( .A(n407), .ZN(n369) );
  XNOR2_X1 U442 ( .A(n668), .B(n404), .ZN(n581) );
  INV_X1 U443 ( .A(KEYINPUT101), .ZN(n404) );
  XNOR2_X1 U444 ( .A(n544), .B(n543), .ZN(n582) );
  NOR2_X1 U445 ( .A1(n559), .A2(n553), .ZN(n544) );
  INV_X1 U446 ( .A(KEYINPUT107), .ZN(n367) );
  XNOR2_X1 U447 ( .A(n402), .B(n401), .ZN(n411) );
  INV_X1 U448 ( .A(KEYINPUT99), .ZN(n401) );
  XNOR2_X1 U449 ( .A(n496), .B(n405), .ZN(n516) );
  XNOR2_X1 U450 ( .A(G475), .B(KEYINPUT13), .ZN(n405) );
  XNOR2_X1 U451 ( .A(G119), .B(G137), .ZN(n423) );
  NOR2_X1 U452 ( .A1(n722), .A2(G952), .ZN(n701) );
  XNOR2_X1 U453 ( .A(KEYINPUT36), .B(KEYINPUT110), .ZN(n571) );
  XNOR2_X1 U454 ( .A(n406), .B(n362), .ZN(n363) );
  NAND2_X1 U455 ( .A1(n390), .A2(n393), .ZN(n389) );
  INV_X1 U456 ( .A(n411), .ZN(n669) );
  OR2_X1 U457 ( .A1(n643), .A2(n642), .ZN(n357) );
  AND2_X1 U458 ( .A1(n502), .A2(n566), .ZN(n358) );
  NOR2_X1 U459 ( .A1(n638), .A2(n369), .ZN(n359) );
  NOR2_X2 U460 ( .A1(n515), .A2(n516), .ZN(n668) );
  NAND2_X1 U461 ( .A1(n730), .A2(KEYINPUT44), .ZN(n523) );
  NAND2_X1 U462 ( .A1(n365), .A2(n407), .ZN(n406) );
  NAND2_X1 U463 ( .A1(n365), .A2(n513), .ZN(n514) );
  NAND2_X1 U464 ( .A1(n365), .A2(n512), .ZN(n402) );
  XNOR2_X2 U465 ( .A(n476), .B(n361), .ZN(n365) );
  XNOR2_X2 U466 ( .A(n374), .B(n375), .ZN(n541) );
  XNOR2_X1 U467 ( .A(n368), .B(n367), .ZN(n552) );
  NAND2_X1 U468 ( .A1(n620), .A2(n368), .ZN(n536) );
  XNOR2_X2 U469 ( .A(n422), .B(G469), .ZN(n368) );
  OR2_X1 U470 ( .A1(n629), .A2(n369), .ZN(n644) );
  XNOR2_X1 U471 ( .A(n500), .B(n360), .ZN(n372) );
  NAND2_X2 U472 ( .A1(n597), .A2(n611), .ZN(n599) );
  XNOR2_X1 U473 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U474 ( .A(G128), .B(G110), .ZN(n426) );
  NOR2_X2 U475 ( .A1(n600), .A2(n528), .ZN(n374) );
  NAND2_X1 U476 ( .A1(n469), .A2(G210), .ZN(n375) );
  NAND2_X1 U477 ( .A1(n620), .A2(n619), .ZN(n376) );
  NOR2_X2 U478 ( .A1(n615), .A2(n616), .ZN(n620) );
  XNOR2_X1 U479 ( .A(n718), .B(G146), .ZN(n377) );
  NOR2_X2 U480 ( .A1(n560), .A2(n475), .ZN(n476) );
  BUF_X1 U481 ( .A(n649), .Z(n379) );
  NAND2_X1 U482 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U483 ( .A(n371), .B(KEYINPUT45), .ZN(n380) );
  XNOR2_X1 U484 ( .A(n527), .B(KEYINPUT45), .ZN(n707) );
  XNOR2_X1 U485 ( .A(n378), .B(n361), .ZN(n511) );
  XNOR2_X1 U486 ( .A(n382), .B(n381), .ZN(n462) );
  XNOR2_X1 U487 ( .A(n460), .B(n458), .ZN(n381) );
  XNOR2_X1 U488 ( .A(n385), .B(n383), .ZN(n382) );
  NAND2_X1 U489 ( .A1(n459), .A2(G224), .ZN(n384) );
  XNOR2_X1 U490 ( .A(n387), .B(n386), .ZN(n385) );
  XNOR2_X2 U491 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n386) );
  XNOR2_X2 U492 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n387) );
  NAND2_X1 U493 ( .A1(n388), .A2(n506), .ZN(n508) );
  NAND2_X1 U494 ( .A1(n355), .A2(KEYINPUT44), .ZN(n509) );
  INV_X1 U495 ( .A(n372), .ZN(n390) );
  NAND2_X1 U496 ( .A1(n505), .A2(n395), .ZN(n394) );
  AND2_X1 U497 ( .A1(n504), .A2(KEYINPUT65), .ZN(n395) );
  XNOR2_X2 U498 ( .A(n396), .B(KEYINPUT32), .ZN(n649) );
  XNOR2_X1 U499 ( .A(n397), .B(n647), .ZN(G75) );
  NAND2_X1 U500 ( .A1(n398), .A2(n722), .ZN(n397) );
  XNOR2_X1 U501 ( .A(n400), .B(n399), .ZN(n398) );
  INV_X1 U502 ( .A(KEYINPUT118), .ZN(n399) );
  NAND2_X1 U503 ( .A1(n646), .A2(n645), .ZN(n400) );
  XNOR2_X2 U504 ( .A(n403), .B(G146), .ZN(n460) );
  XNOR2_X2 U505 ( .A(G143), .B(G128), .ZN(n458) );
  NAND2_X1 U506 ( .A1(n372), .A2(n520), .ZN(n648) );
  INV_X1 U507 ( .A(n412), .ZN(n410) );
  NAND2_X1 U508 ( .A1(n351), .A2(n679), .ZN(n680) );
  NAND2_X1 U509 ( .A1(n351), .A2(n668), .ZN(n682) );
  XOR2_X1 U510 ( .A(n427), .B(n426), .Z(n413) );
  INV_X1 U511 ( .A(KEYINPUT86), .ZN(n529) );
  XNOR2_X1 U512 ( .A(n530), .B(n529), .ZN(n591) );
  INV_X1 U513 ( .A(KEYINPUT48), .ZN(n578) );
  XNOR2_X1 U514 ( .A(n578), .B(KEYINPUT70), .ZN(n579) );
  XNOR2_X1 U515 ( .A(G478), .B(KEYINPUT100), .ZN(n485) );
  XNOR2_X1 U516 ( .A(KEYINPUT75), .B(KEYINPUT39), .ZN(n543) );
  XNOR2_X1 U517 ( .A(G107), .B(G104), .ZN(n416) );
  XNOR2_X1 U518 ( .A(G110), .B(KEYINPUT93), .ZN(n415) );
  XNOR2_X1 U519 ( .A(n416), .B(n415), .ZN(n702) );
  XNOR2_X1 U520 ( .A(n446), .B(KEYINPUT74), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n702), .B(n417), .ZN(n461) );
  BUF_X2 U522 ( .A(n459), .Z(n722) );
  NAND2_X1 U523 ( .A1(G227), .A2(n722), .ZN(n418) );
  XOR2_X1 U524 ( .A(n419), .B(n418), .Z(n420) );
  XNOR2_X1 U525 ( .A(n461), .B(n420), .ZN(n421) );
  XNOR2_X1 U526 ( .A(n452), .B(n421), .ZN(n690) );
  INV_X1 U527 ( .A(G902), .ZN(n453) );
  NAND2_X1 U528 ( .A1(n690), .A2(n453), .ZN(n422) );
  XNOR2_X1 U529 ( .A(n423), .B(KEYINPUT23), .ZN(n432) );
  XOR2_X1 U530 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n425) );
  NAND2_X1 U531 ( .A1(G234), .A2(n722), .ZN(n424) );
  XNOR2_X1 U532 ( .A(n425), .B(n424), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n482), .A2(G221), .ZN(n430) );
  XOR2_X1 U534 ( .A(KEYINPUT79), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U535 ( .A(n717), .B(n413), .ZN(n429) );
  XNOR2_X1 U536 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U537 ( .A(n432), .B(n431), .ZN(n698) );
  XNOR2_X1 U538 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n433) );
  XNOR2_X1 U539 ( .A(n433), .B(G902), .ZN(n592) );
  NAND2_X1 U540 ( .A1(n592), .A2(G234), .ZN(n434) );
  XNOR2_X1 U541 ( .A(KEYINPUT20), .B(n434), .ZN(n438) );
  NAND2_X1 U542 ( .A1(G217), .A2(n438), .ZN(n435) );
  XNOR2_X2 U543 ( .A(n437), .B(n436), .ZN(n615) );
  XOR2_X1 U544 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n440) );
  NAND2_X1 U545 ( .A1(n438), .A2(G221), .ZN(n439) );
  XNOR2_X1 U546 ( .A(n440), .B(n439), .ZN(n616) );
  XNOR2_X1 U547 ( .A(KEYINPUT3), .B(G119), .ZN(n442) );
  XNOR2_X1 U548 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n442), .B(n441), .ZN(n445) );
  XNOR2_X1 U550 ( .A(G116), .B(G113), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n443), .B(KEYINPUT94), .ZN(n444) );
  XNOR2_X1 U552 ( .A(n445), .B(n444), .ZN(n465) );
  NOR2_X1 U553 ( .A1(G953), .A2(G237), .ZN(n487) );
  NAND2_X1 U554 ( .A1(n487), .A2(G210), .ZN(n447) );
  XNOR2_X1 U555 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U556 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n448) );
  XNOR2_X1 U557 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U558 ( .A(n465), .B(n450), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n377), .B(n451), .ZN(n653) );
  NAND2_X1 U560 ( .A1(n653), .A2(n453), .ZN(n455) );
  INV_X1 U561 ( .A(G472), .ZN(n454) );
  XNOR2_X2 U562 ( .A(n455), .B(n454), .ZN(n549) );
  INV_X1 U563 ( .A(KEYINPUT6), .ZN(n456) );
  XNOR2_X1 U564 ( .A(n462), .B(n461), .ZN(n466) );
  XNOR2_X1 U565 ( .A(KEYINPUT16), .B(G122), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n463), .B(KEYINPUT77), .ZN(n464) );
  XNOR2_X1 U567 ( .A(n465), .B(n464), .ZN(n704) );
  XNOR2_X1 U568 ( .A(n466), .B(n704), .ZN(n600) );
  INV_X1 U569 ( .A(n592), .ZN(n528) );
  NOR2_X1 U570 ( .A1(G237), .A2(G902), .ZN(n468) );
  INV_X1 U571 ( .A(KEYINPUT78), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U573 ( .A1(G234), .A2(G237), .ZN(n470) );
  XNOR2_X1 U574 ( .A(n470), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U575 ( .A1(n473), .A2(G952), .ZN(n471) );
  XOR2_X1 U576 ( .A(KEYINPUT95), .B(n471), .Z(n643) );
  NOR2_X1 U577 ( .A1(n643), .A2(G953), .ZN(n535) );
  NOR2_X1 U578 ( .A1(G898), .A2(n722), .ZN(n472) );
  XOR2_X1 U579 ( .A(KEYINPUT96), .B(n472), .Z(n705) );
  NAND2_X1 U580 ( .A1(G902), .A2(n473), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n705), .A2(n531), .ZN(n474) );
  XNOR2_X1 U582 ( .A(G116), .B(G122), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n477), .B(KEYINPUT7), .ZN(n478) );
  XOR2_X1 U584 ( .A(n478), .B(KEYINPUT9), .Z(n481) );
  XNOR2_X1 U585 ( .A(n479), .B(G107), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n484) );
  NAND2_X1 U587 ( .A1(G217), .A2(n482), .ZN(n483) );
  XOR2_X1 U588 ( .A(n484), .B(n483), .Z(n694) );
  NOR2_X1 U589 ( .A1(G902), .A2(n694), .ZN(n486) );
  XNOR2_X2 U590 ( .A(n486), .B(n485), .ZN(n515) );
  NAND2_X1 U591 ( .A1(G214), .A2(n487), .ZN(n488) );
  XNOR2_X1 U592 ( .A(n717), .B(n488), .ZN(n495) );
  XNOR2_X1 U593 ( .A(n489), .B(G122), .ZN(n493) );
  XNOR2_X1 U594 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U595 ( .A(n493), .B(n492), .Z(n494) );
  XNOR2_X1 U596 ( .A(n495), .B(n494), .ZN(n660) );
  NOR2_X1 U597 ( .A1(G902), .A2(n660), .ZN(n496) );
  INV_X1 U598 ( .A(n516), .ZN(n497) );
  NOR2_X1 U599 ( .A1(n515), .A2(n497), .ZN(n557) );
  INV_X1 U600 ( .A(n730), .ZN(n506) );
  NAND2_X1 U601 ( .A1(n515), .A2(n497), .ZN(n633) );
  NOR2_X1 U602 ( .A1(n633), .A2(n616), .ZN(n498) );
  XNOR2_X1 U603 ( .A(n498), .B(KEYINPUT102), .ZN(n499) );
  NAND2_X1 U604 ( .A1(n352), .A2(n615), .ZN(n501) );
  XNOR2_X1 U605 ( .A(n501), .B(KEYINPUT103), .ZN(n502) );
  OR2_X1 U606 ( .A1(n352), .A2(n625), .ZN(n503) );
  INV_X1 U607 ( .A(n503), .ZN(n504) );
  INV_X1 U608 ( .A(KEYINPUT44), .ZN(n507) );
  NAND2_X1 U609 ( .A1(n508), .A2(n507), .ZN(n510) );
  NOR2_X1 U610 ( .A1(n625), .A2(n536), .ZN(n512) );
  AND2_X1 U611 ( .A1(n516), .A2(n515), .ZN(n679) );
  XNOR2_X1 U612 ( .A(KEYINPUT85), .B(n635), .ZN(n517) );
  INV_X1 U613 ( .A(n615), .ZN(n518) );
  NAND2_X1 U614 ( .A1(n566), .A2(n518), .ZN(n519) );
  AND2_X1 U615 ( .A1(n521), .A2(n648), .ZN(n522) );
  NAND2_X1 U616 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n707), .A2(n528), .ZN(n530) );
  OR2_X1 U618 ( .A1(n722), .A2(n531), .ZN(n532) );
  XNOR2_X1 U619 ( .A(KEYINPUT104), .B(n532), .ZN(n533) );
  NOR2_X1 U620 ( .A1(G900), .A2(n533), .ZN(n534) );
  NOR2_X1 U621 ( .A1(n535), .A2(n534), .ZN(n547) );
  NAND2_X1 U622 ( .A1(n625), .A2(n630), .ZN(n538) );
  XOR2_X1 U623 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n537) );
  XNOR2_X1 U624 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U625 ( .A1(n540), .A2(n539), .ZN(n559) );
  BUF_X1 U626 ( .A(n541), .Z(n542) );
  XNOR2_X1 U627 ( .A(n542), .B(KEYINPUT38), .ZN(n553) );
  XNOR2_X1 U628 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n545) );
  XNOR2_X1 U629 ( .A(n546), .B(n545), .ZN(n729) );
  NOR2_X1 U630 ( .A1(n547), .A2(n616), .ZN(n548) );
  NAND2_X1 U631 ( .A1(n615), .A2(n548), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n567), .A2(n549), .ZN(n550) );
  XNOR2_X1 U633 ( .A(KEYINPUT28), .B(n550), .ZN(n551) );
  NAND2_X1 U634 ( .A1(n552), .A2(n551), .ZN(n561) );
  INV_X1 U635 ( .A(n553), .ZN(n631) );
  NAND2_X1 U636 ( .A1(n631), .A2(n630), .ZN(n634) );
  NOR2_X1 U637 ( .A1(n633), .A2(n634), .ZN(n554) );
  XNOR2_X1 U638 ( .A(n554), .B(KEYINPUT41), .ZN(n629) );
  NOR2_X1 U639 ( .A1(n561), .A2(n629), .ZN(n555) );
  XNOR2_X1 U640 ( .A(n555), .B(KEYINPUT42), .ZN(n732) );
  NAND2_X1 U641 ( .A1(n557), .A2(n542), .ZN(n558) );
  NOR2_X1 U642 ( .A1(n559), .A2(n558), .ZN(n676) );
  NOR2_X1 U643 ( .A1(n561), .A2(n560), .ZN(n677) );
  NOR2_X1 U644 ( .A1(KEYINPUT47), .A2(KEYINPUT85), .ZN(n562) );
  XNOR2_X1 U645 ( .A(n562), .B(n635), .ZN(n563) );
  NAND2_X1 U646 ( .A1(n677), .A2(n563), .ZN(n565) );
  OR2_X1 U647 ( .A1(n677), .A2(KEYINPUT47), .ZN(n564) );
  NAND2_X1 U648 ( .A1(n565), .A2(n564), .ZN(n574) );
  NOR2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U650 ( .A(KEYINPUT109), .B(n583), .ZN(n570) );
  NOR2_X1 U651 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n573), .A2(n352), .ZN(n684) );
  NAND2_X1 U653 ( .A1(n574), .A2(n684), .ZN(n575) );
  NOR2_X1 U654 ( .A1(n676), .A2(n575), .ZN(n576) );
  XNOR2_X1 U655 ( .A(KEYINPUT71), .B(n576), .ZN(n577) );
  XNOR2_X1 U656 ( .A(n580), .B(n579), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n685) );
  NAND2_X1 U658 ( .A1(n583), .A2(n630), .ZN(n584) );
  XOR2_X1 U659 ( .A(KEYINPUT105), .B(n584), .Z(n585) );
  NOR2_X1 U660 ( .A1(n352), .A2(n585), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n586), .B(KEYINPUT43), .ZN(n587) );
  OR2_X1 U662 ( .A1(n587), .A2(n542), .ZN(n650) );
  NAND2_X1 U663 ( .A1(n685), .A2(n650), .ZN(n588) );
  OR2_X2 U664 ( .A1(n589), .A2(n588), .ZN(n720) );
  INV_X1 U665 ( .A(n720), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT88), .B(n592), .Z(n593) );
  NAND2_X1 U668 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U670 ( .A(n380), .ZN(n596) );
  NOR2_X2 U671 ( .A1(n596), .A2(n720), .ZN(n608) );
  NAND2_X1 U672 ( .A1(n608), .A2(KEYINPUT2), .ZN(n611) );
  INV_X1 U673 ( .A(KEYINPUT64), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n686), .A2(G210), .ZN(n605) );
  BUF_X1 U675 ( .A(n600), .Z(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n602) );
  XOR2_X1 U677 ( .A(n602), .B(KEYINPUT120), .Z(n603) );
  XNOR2_X1 U678 ( .A(n605), .B(n604), .ZN(n606) );
  NOR2_X2 U679 ( .A1(n606), .A2(n701), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U681 ( .A(KEYINPUT84), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U684 ( .A(KEYINPUT87), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n614), .B(n613), .ZN(n646) );
  XOR2_X1 U686 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n618) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(n623) );
  NOR2_X1 U689 ( .A1(n620), .A2(n352), .ZN(n621) );
  XOR2_X1 U690 ( .A(KEYINPUT50), .B(n621), .Z(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U692 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U693 ( .A1(n513), .A2(n626), .ZN(n627) );
  XOR2_X1 U694 ( .A(KEYINPUT51), .B(n627), .Z(n628) );
  NOR2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n639) );
  NOR2_X1 U696 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n637) );
  NOR2_X1 U698 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U699 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U700 ( .A1(n639), .A2(n359), .ZN(n640) );
  XOR2_X1 U701 ( .A(n640), .B(KEYINPUT117), .Z(n641) );
  XNOR2_X1 U702 ( .A(KEYINPUT52), .B(n641), .ZN(n642) );
  AND2_X1 U703 ( .A1(n644), .A2(n357), .ZN(n645) );
  XNOR2_X1 U704 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n647) );
  XNOR2_X1 U705 ( .A(n648), .B(G101), .ZN(G3) );
  XNOR2_X1 U706 ( .A(n379), .B(G119), .ZN(G21) );
  XNOR2_X1 U707 ( .A(n650), .B(G140), .ZN(G42) );
  XNOR2_X1 U708 ( .A(n651), .B(G110), .ZN(G12) );
  NAND2_X1 U709 ( .A1(n373), .A2(G472), .ZN(n655) );
  XNOR2_X1 U710 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n652) );
  XNOR2_X1 U711 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U712 ( .A1(n656), .A2(n701), .ZN(n658) );
  XOR2_X1 U713 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n657) );
  XNOR2_X1 U714 ( .A(n658), .B(n657), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n373), .A2(G475), .ZN(n662) );
  XNOR2_X1 U716 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n659) );
  XNOR2_X1 U717 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X2 U718 ( .A1(n663), .A2(n701), .ZN(n665) );
  XNOR2_X1 U719 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n664) );
  XNOR2_X1 U720 ( .A(n665), .B(n664), .ZN(G60) );
  XOR2_X1 U721 ( .A(G104), .B(KEYINPUT113), .Z(n667) );
  NAND2_X1 U722 ( .A1(n669), .A2(n679), .ZN(n666) );
  XNOR2_X1 U723 ( .A(n667), .B(n666), .ZN(G6) );
  XNOR2_X1 U724 ( .A(G107), .B(KEYINPUT114), .ZN(n673) );
  XOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n671) );
  NAND2_X1 U726 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U728 ( .A(n673), .B(n672), .ZN(G9) );
  XOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U730 ( .A1(n677), .A2(n668), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n675), .B(n674), .ZN(G30) );
  XOR2_X1 U732 ( .A(G143), .B(n676), .Z(G45) );
  NAND2_X1 U733 ( .A1(n677), .A2(n679), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n678), .B(G146), .ZN(G48) );
  XOR2_X1 U735 ( .A(G113), .B(KEYINPUT115), .Z(n681) );
  XNOR2_X1 U736 ( .A(n681), .B(n680), .ZN(G15) );
  XNOR2_X1 U737 ( .A(n682), .B(G116), .ZN(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n683) );
  XNOR2_X1 U739 ( .A(n684), .B(n683), .ZN(G27) );
  XNOR2_X1 U740 ( .A(G134), .B(n685), .ZN(G36) );
  BUF_X1 U741 ( .A(n686), .Z(n697) );
  NAND2_X1 U742 ( .A1(n697), .A2(G469), .ZN(n692) );
  XOR2_X1 U743 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n688) );
  XNOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n701), .A2(n693), .ZN(G54) );
  NAND2_X1 U749 ( .A1(n697), .A2(G478), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U751 ( .A1(n701), .A2(n696), .ZN(G63) );
  NAND2_X1 U752 ( .A1(n697), .A2(G217), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n701), .A2(n700), .ZN(G66) );
  XNOR2_X1 U755 ( .A(n702), .B(G101), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n706), .A2(n705), .ZN(n715) );
  BUF_X1 U758 ( .A(n380), .Z(n708) );
  NAND2_X1 U759 ( .A1(n708), .A2(n722), .ZN(n713) );
  NAND2_X1 U760 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(KEYINPUT124), .ZN(n710) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U763 ( .A1(G898), .A2(n711), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U766 ( .A(KEYINPUT125), .B(n716), .ZN(G69) );
  XNOR2_X1 U767 ( .A(n717), .B(KEYINPUT126), .ZN(n719) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n724) );
  XNOR2_X1 U769 ( .A(KEYINPUT127), .B(n724), .ZN(n721) );
  XOR2_X1 U770 ( .A(n721), .B(n720), .Z(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(n722), .ZN(n728) );
  XNOR2_X1 U772 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(G72) );
  XOR2_X1 U776 ( .A(G131), .B(n729), .Z(G33) );
  BUF_X1 U777 ( .A(n730), .Z(n731) );
  XOR2_X1 U778 ( .A(n731), .B(G122), .Z(G24) );
  XOR2_X1 U779 ( .A(G137), .B(n732), .Z(G39) );
endmodule

