

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U320 ( .A(KEYINPUT107), .B(KEYINPUT47), .ZN(n288) );
  XOR2_X1 U321 ( .A(n338), .B(n337), .Z(n289) );
  XNOR2_X1 U322 ( .A(KEYINPUT48), .B(KEYINPUT108), .ZN(n496) );
  XNOR2_X1 U323 ( .A(n339), .B(n289), .ZN(n340) );
  XNOR2_X1 U324 ( .A(n497), .B(n496), .ZN(n531) );
  XNOR2_X1 U325 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U326 ( .A(KEYINPUT41), .B(n570), .Z(n550) );
  XOR2_X1 U327 ( .A(n427), .B(n396), .Z(n543) );
  XOR2_X1 U328 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n291) );
  XNOR2_X1 U329 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n290) );
  XNOR2_X1 U330 ( .A(n291), .B(n290), .ZN(n301) );
  XOR2_X1 U331 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n299) );
  XOR2_X1 U332 ( .A(G127GAT), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U333 ( .A(G113GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n383) );
  XNOR2_X1 U335 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n294), .B(KEYINPUT3), .ZN(n295) );
  XOR2_X1 U337 ( .A(n295), .B(KEYINPUT2), .Z(n297) );
  XNOR2_X1 U338 ( .A(G141GAT), .B(G155GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n416) );
  XNOR2_X1 U340 ( .A(n383), .B(n416), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n313) );
  NAND2_X1 U343 ( .A1(G225GAT), .A2(G233GAT), .ZN(n307) );
  XOR2_X1 U344 ( .A(G148GAT), .B(G120GAT), .Z(n303) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(G1GAT), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U347 ( .A(G162GAT), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U350 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n309) );
  XNOR2_X1 U351 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U353 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U354 ( .A(n313), .B(n312), .Z(n515) );
  INV_X1 U355 ( .A(n515), .ZN(n533) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G43GAT), .Z(n315) );
  XNOR2_X1 U357 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n314) );
  XNOR2_X1 U358 ( .A(n315), .B(n314), .ZN(n371) );
  XNOR2_X1 U359 ( .A(G22GAT), .B(G15GAT), .ZN(n316) );
  XNOR2_X1 U360 ( .A(n316), .B(G1GAT), .ZN(n359) );
  XNOR2_X1 U361 ( .A(n371), .B(n359), .ZN(n329) );
  XOR2_X1 U362 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n318) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U365 ( .A(n319), .B(KEYINPUT66), .Z(n327) );
  XOR2_X1 U366 ( .A(G141GAT), .B(G197GAT), .Z(n321) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G50GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U369 ( .A(G8GAT), .B(KEYINPUT67), .Z(n323) );
  XNOR2_X1 U370 ( .A(G169GAT), .B(G113GAT), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U374 ( .A(n329), .B(n328), .Z(n517) );
  INV_X1 U375 ( .A(n517), .ZN(n566) );
  XOR2_X1 U376 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n331) );
  NAND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U379 ( .A(n332), .B(KEYINPUT71), .Z(n336) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U381 ( .A(n333), .B(G148GAT), .ZN(n403) );
  XNOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n334), .B(KEYINPUT13), .ZN(n358) );
  XNOR2_X1 U384 ( .A(n403), .B(n358), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U386 ( .A(G120GAT), .B(G71GAT), .Z(n384) );
  XOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .Z(n375) );
  XNOR2_X1 U388 ( .A(n384), .B(n375), .ZN(n339) );
  XOR2_X1 U389 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n338) );
  XNOR2_X1 U390 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n337) );
  XOR2_X1 U391 ( .A(KEYINPUT70), .B(G64GAT), .Z(n343) );
  XNOR2_X1 U392 ( .A(G204GAT), .B(G92GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U394 ( .A(G176GAT), .B(n344), .Z(n420) );
  XNOR2_X1 U395 ( .A(n345), .B(n420), .ZN(n570) );
  INV_X1 U396 ( .A(n570), .ZN(n346) );
  NOR2_X1 U397 ( .A1(n566), .A2(n346), .ZN(n455) );
  XOR2_X1 U398 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n379) );
  XOR2_X1 U399 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n363) );
  XOR2_X1 U402 ( .A(G8GAT), .B(G183GAT), .Z(n417) );
  XOR2_X1 U403 ( .A(G211GAT), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U404 ( .A(G127GAT), .B(G155GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U406 ( .A(n417), .B(n351), .Z(n353) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U409 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U412 ( .A(n357), .B(n356), .Z(n361) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n574) );
  INV_X1 U416 ( .A(n574), .ZN(n525) );
  XOR2_X1 U417 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n365) );
  XNOR2_X1 U418 ( .A(G134GAT), .B(G106GAT), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n368) );
  XOR2_X1 U420 ( .A(G50GAT), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U421 ( .A(n408), .B(G92GAT), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n366), .B(KEYINPUT10), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT74), .B(G218GAT), .Z(n370) );
  XNOR2_X1 U425 ( .A(G36GAT), .B(G190GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n422) );
  XNOR2_X1 U427 ( .A(n371), .B(n422), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U429 ( .A(n375), .B(n374), .Z(n377) );
  NAND2_X1 U430 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XOR2_X1 U431 ( .A(n377), .B(n376), .Z(n527) );
  INV_X1 U432 ( .A(n527), .ZN(n560) );
  NAND2_X1 U433 ( .A1(n525), .A2(n560), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n442) );
  XOR2_X1 U435 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(G169GAT), .B(n382), .Z(n427) );
  XOR2_X1 U439 ( .A(n384), .B(n383), .Z(n386) );
  XNOR2_X1 U440 ( .A(G190GAT), .B(G99GAT), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U442 ( .A(KEYINPUT79), .B(KEYINPUT64), .Z(n388) );
  NAND2_X1 U443 ( .A1(G227GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U445 ( .A(n390), .B(n389), .Z(n395) );
  XOR2_X1 U446 ( .A(G183GAT), .B(KEYINPUT20), .Z(n392) );
  XNOR2_X1 U447 ( .A(G43GAT), .B(G15GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n393), .B(G176GAT), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  INV_X1 U451 ( .A(n543), .ZN(n548) );
  XOR2_X1 U452 ( .A(KEYINPUT24), .B(G204GAT), .Z(n398) );
  XNOR2_X1 U453 ( .A(KEYINPUT88), .B(KEYINPUT81), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U455 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n400) );
  XNOR2_X1 U456 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U458 ( .A(n402), .B(n401), .Z(n414) );
  XOR2_X1 U459 ( .A(n403), .B(G22GAT), .Z(n405) );
  NAND2_X1 U460 ( .A1(G228GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n412) );
  XOR2_X1 U462 ( .A(G211GAT), .B(KEYINPUT82), .Z(n407) );
  XNOR2_X1 U463 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n423) );
  XOR2_X1 U465 ( .A(KEYINPUT23), .B(n423), .Z(n410) );
  XNOR2_X1 U466 ( .A(G218GAT), .B(n408), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n535) );
  XOR2_X1 U471 ( .A(KEYINPUT28), .B(n535), .Z(n482) );
  AND2_X1 U472 ( .A1(n515), .A2(n482), .ZN(n429) );
  XNOR2_X1 U473 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n428) );
  XOR2_X1 U474 ( .A(KEYINPUT94), .B(n417), .Z(n419) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U477 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n530) );
  XNOR2_X1 U481 ( .A(n428), .B(n530), .ZN(n433) );
  NAND2_X1 U482 ( .A1(n429), .A2(n433), .ZN(n498) );
  XNOR2_X1 U483 ( .A(KEYINPUT96), .B(n498), .ZN(n430) );
  NOR2_X1 U484 ( .A1(n548), .A2(n430), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n431), .B(KEYINPUT97), .ZN(n441) );
  NAND2_X1 U486 ( .A1(n535), .A2(n543), .ZN(n432) );
  XOR2_X1 U487 ( .A(KEYINPUT26), .B(n432), .Z(n564) );
  NAND2_X1 U488 ( .A1(n564), .A2(n433), .ZN(n513) );
  XNOR2_X1 U489 ( .A(n513), .B(KEYINPUT98), .ZN(n438) );
  NOR2_X1 U490 ( .A1(n543), .A2(n530), .ZN(n434) );
  NOR2_X1 U491 ( .A1(n535), .A2(n434), .ZN(n435) );
  XOR2_X1 U492 ( .A(n435), .B(KEYINPUT99), .Z(n436) );
  XNOR2_X1 U493 ( .A(KEYINPUT25), .B(n436), .ZN(n437) );
  NAND2_X1 U494 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND2_X1 U495 ( .A1(n439), .A2(n533), .ZN(n440) );
  NAND2_X1 U496 ( .A1(n441), .A2(n440), .ZN(n452) );
  AND2_X1 U497 ( .A1(n442), .A2(n452), .ZN(n466) );
  NAND2_X1 U498 ( .A1(n455), .A2(n466), .ZN(n449) );
  NOR2_X1 U499 ( .A1(n533), .A2(n449), .ZN(n444) );
  XNOR2_X1 U500 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U502 ( .A(G1GAT), .B(n445), .Z(G1324GAT) );
  NOR2_X1 U503 ( .A1(n530), .A2(n449), .ZN(n446) );
  XOR2_X1 U504 ( .A(G8GAT), .B(n446), .Z(G1325GAT) );
  NOR2_X1 U505 ( .A1(n543), .A2(n449), .ZN(n448) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(G1326GAT) );
  NOR2_X1 U508 ( .A1(n482), .A2(n449), .ZN(n451) );
  XNOR2_X1 U509 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(G1327GAT) );
  XOR2_X1 U511 ( .A(n527), .B(KEYINPUT36), .Z(n578) );
  NAND2_X1 U512 ( .A1(n574), .A2(n452), .ZN(n453) );
  NOR2_X1 U513 ( .A1(n578), .A2(n453), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT37), .B(n454), .Z(n476) );
  NAND2_X1 U515 ( .A1(n476), .A2(n455), .ZN(n456) );
  XNOR2_X1 U516 ( .A(KEYINPUT38), .B(n456), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n464), .A2(n533), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n458) );
  XNOR2_X1 U519 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  NOR2_X1 U522 ( .A1(n464), .A2(n530), .ZN(n461) );
  XOR2_X1 U523 ( .A(G36GAT), .B(n461), .Z(G1329GAT) );
  NOR2_X1 U524 ( .A1(n543), .A2(n464), .ZN(n462) );
  XOR2_X1 U525 ( .A(KEYINPUT40), .B(n462), .Z(n463) );
  XNOR2_X1 U526 ( .A(G43GAT), .B(n463), .ZN(G1330GAT) );
  NOR2_X1 U527 ( .A1(n464), .A2(n482), .ZN(n465) );
  XOR2_X1 U528 ( .A(G50GAT), .B(n465), .Z(G1331GAT) );
  NOR2_X1 U529 ( .A1(n517), .A2(n550), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n475), .A2(n466), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n533), .A2(n471), .ZN(n467) );
  XOR2_X1 U532 ( .A(G57GAT), .B(n467), .Z(n468) );
  XNOR2_X1 U533 ( .A(KEYINPUT42), .B(n468), .ZN(G1332GAT) );
  NOR2_X1 U534 ( .A1(n530), .A2(n471), .ZN(n469) );
  XOR2_X1 U535 ( .A(G64GAT), .B(n469), .Z(G1333GAT) );
  NOR2_X1 U536 ( .A1(n543), .A2(n471), .ZN(n470) );
  XOR2_X1 U537 ( .A(G71GAT), .B(n470), .Z(G1334GAT) );
  NOR2_X1 U538 ( .A1(n482), .A2(n471), .ZN(n473) );
  XNOR2_X1 U539 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n472) );
  XNOR2_X1 U540 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U541 ( .A(G78GAT), .B(n474), .ZN(G1335GAT) );
  NAND2_X1 U542 ( .A1(n476), .A2(n475), .ZN(n481) );
  NOR2_X1 U543 ( .A1(n533), .A2(n481), .ZN(n478) );
  XNOR2_X1 U544 ( .A(G85GAT), .B(KEYINPUT105), .ZN(n477) );
  XNOR2_X1 U545 ( .A(n478), .B(n477), .ZN(G1336GAT) );
  NOR2_X1 U546 ( .A1(n530), .A2(n481), .ZN(n479) );
  XOR2_X1 U547 ( .A(G92GAT), .B(n479), .Z(G1337GAT) );
  NOR2_X1 U548 ( .A1(n543), .A2(n481), .ZN(n480) );
  XOR2_X1 U549 ( .A(G99GAT), .B(n480), .Z(G1338GAT) );
  NOR2_X1 U550 ( .A1(n482), .A2(n481), .ZN(n484) );
  XNOR2_X1 U551 ( .A(KEYINPUT44), .B(KEYINPUT106), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U553 ( .A(G106GAT), .B(n485), .Z(G1339GAT) );
  NOR2_X1 U554 ( .A1(n566), .A2(n550), .ZN(n486) );
  XNOR2_X1 U555 ( .A(n486), .B(KEYINPUT46), .ZN(n487) );
  NOR2_X1 U556 ( .A1(n487), .A2(n525), .ZN(n488) );
  AND2_X1 U557 ( .A1(n488), .A2(n560), .ZN(n489) );
  XNOR2_X1 U558 ( .A(n489), .B(n288), .ZN(n495) );
  NOR2_X1 U559 ( .A1(n574), .A2(n578), .ZN(n491) );
  XNOR2_X1 U560 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n490) );
  XNOR2_X1 U561 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U562 ( .A1(n570), .A2(n566), .ZN(n492) );
  NOR2_X1 U563 ( .A1(n493), .A2(n492), .ZN(n494) );
  NOR2_X1 U564 ( .A1(n495), .A2(n494), .ZN(n497) );
  NOR2_X1 U565 ( .A1(n531), .A2(n498), .ZN(n499) );
  NAND2_X1 U566 ( .A1(n548), .A2(n499), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(KEYINPUT109), .ZN(n510) );
  NAND2_X1 U568 ( .A1(n517), .A2(n510), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n501), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U570 ( .A(G120GAT), .B(KEYINPUT110), .Z(n503) );
  INV_X1 U571 ( .A(n550), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n510), .A2(n522), .ZN(n502) );
  XNOR2_X1 U573 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U574 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n504) );
  XNOR2_X1 U575 ( .A(n505), .B(n504), .ZN(G1341GAT) );
  XNOR2_X1 U576 ( .A(G127GAT), .B(KEYINPUT112), .ZN(n509) );
  XOR2_X1 U577 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n507) );
  NAND2_X1 U578 ( .A1(n510), .A2(n525), .ZN(n506) );
  XNOR2_X1 U579 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U580 ( .A(n509), .B(n508), .ZN(G1342GAT) );
  XOR2_X1 U581 ( .A(G134GAT), .B(KEYINPUT51), .Z(n512) );
  NAND2_X1 U582 ( .A1(n510), .A2(n527), .ZN(n511) );
  XNOR2_X1 U583 ( .A(n512), .B(n511), .ZN(G1343GAT) );
  NOR2_X1 U584 ( .A1(n531), .A2(n513), .ZN(n514) );
  NAND2_X1 U585 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n516), .Z(n528) );
  NAND2_X1 U587 ( .A1(n517), .A2(n528), .ZN(n518) );
  XNOR2_X1 U588 ( .A(G141GAT), .B(n518), .ZN(G1344GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n520) );
  XNOR2_X1 U590 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n519) );
  XNOR2_X1 U591 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U592 ( .A(KEYINPUT52), .B(n521), .Z(n524) );
  NAND2_X1 U593 ( .A1(n522), .A2(n528), .ZN(n523) );
  XNOR2_X1 U594 ( .A(n524), .B(n523), .ZN(G1345GAT) );
  NAND2_X1 U595 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n526), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n529), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(KEYINPUT54), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n563) );
  NOR2_X1 U602 ( .A1(n535), .A2(n563), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n540) );
  INV_X1 U605 ( .A(n540), .ZN(n539) );
  INV_X1 U606 ( .A(KEYINPUT55), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U608 ( .A1(KEYINPUT55), .A2(n540), .ZN(n541) );
  NAND2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n549) );
  NOR2_X1 U610 ( .A1(n566), .A2(n543), .ZN(n544) );
  AND2_X1 U611 ( .A1(n549), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G169GAT), .B(n547), .ZN(G1348GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n550), .A2(n559), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(KEYINPUT56), .B(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NOR2_X1 U622 ( .A1(n574), .A2(n559), .ZN(n556) );
  XOR2_X1 U623 ( .A(G183GAT), .B(n556), .Z(G1350GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n558) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(G1351GAT) );
  INV_X1 U629 ( .A(n563), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n566), .A2(n577), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n577), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(n575), .Z(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

