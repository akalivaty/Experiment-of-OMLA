//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n204), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(KEYINPUT66), .B1(new_n217), .B2(new_n218), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n206), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n210), .B(new_n215), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n221), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND3_X1  g0051(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n213), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n203), .B2(G20), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(new_n256), .B2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR3_X1   g0060(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n204), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT69), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n255), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n257), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n272), .A2(new_n203), .A3(G274), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G226), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1698), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G222), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G223), .A3(G1698), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n281), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G77), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n272), .B1(new_n291), .B2(new_n292), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n280), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(G190), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n270), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n270), .A2(new_n297), .A3(new_n301), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n269), .C1(G169), .C2(new_n295), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G68), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n266), .ZN(new_n310));
  INV_X1    g0110(.A(G77), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n255), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT11), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OR3_X1    g0115(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n317));
  AOI22_X1  g0117(.A1(G68), .A2(new_n256), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n315), .A2(new_n318), .A3(new_n322), .A4(new_n319), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n277), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n221), .A2(G1698), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n288), .C2(new_n281), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n272), .A2(G238), .A3(new_n278), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n276), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n327), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n272), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n276), .A2(new_n336), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT13), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n326), .B(G169), .C1(new_n338), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n335), .A2(new_n337), .A3(new_n327), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(G179), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n338), .A2(new_n341), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT14), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n325), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n342), .A2(new_n345), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n348), .B1(new_n343), .B2(new_n344), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n326), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT72), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n324), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n320), .B1(new_n347), .B2(G190), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n347), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n286), .B2(G20), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n308), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n220), .A2(new_n308), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G58), .A2(G68), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n259), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n360), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT7), .B1(new_n289), .B2(new_n204), .ZN(new_n371));
  NOR4_X1   g0171(.A1(new_n288), .A2(new_n281), .A3(new_n361), .A4(G20), .ZN(new_n372));
  OAI21_X1  g0172(.A(G68), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n369), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(KEYINPUT16), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n375), .A3(new_n255), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n268), .B1(G1), .B2(new_n204), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n264), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n252), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n264), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n265), .A2(new_n225), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G223), .A2(G1698), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n277), .B2(G1698), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n383), .B1(new_n385), .B2(new_n286), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(new_n272), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n277), .A2(G1698), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G223), .B2(G1698), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n389), .A2(new_n289), .B1(new_n265), .B2(new_n225), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(KEYINPUT74), .A3(new_n334), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n272), .A2(G232), .A3(new_n278), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n276), .A2(new_n392), .A3(new_n304), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n387), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n387), .A2(new_n391), .A3(KEYINPUT75), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n276), .A2(new_n392), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n272), .B2(new_n386), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n348), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n381), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT18), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n396), .A2(new_n397), .B1(new_n348), .B2(new_n400), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n381), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n400), .A2(new_n357), .ZN(new_n407));
  INV_X1    g0207(.A(G190), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n387), .A2(new_n391), .A3(new_n408), .A4(new_n399), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(new_n376), .A3(new_n380), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n410), .A2(new_n376), .A3(KEYINPUT17), .A4(new_n380), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n403), .A2(new_n406), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n284), .A2(G232), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n286), .A2(G238), .A3(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n289), .A2(G107), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n334), .ZN(new_n420));
  INV_X1    g0220(.A(new_n276), .ZN(new_n421));
  INV_X1    g0221(.A(new_n279), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(G244), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n426), .A2(new_n310), .B1(new_n204), .B2(new_n311), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT70), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n263), .B(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(new_n260), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n255), .B1(new_n311), .B2(new_n379), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT71), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n377), .B2(new_n311), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n256), .A2(KEYINPUT71), .A3(G77), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n420), .A2(new_n423), .A3(G190), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n425), .A2(new_n432), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n424), .A2(new_n348), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n379), .A2(new_n311), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n263), .B(KEYINPUT70), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n427), .B1(new_n441), .B2(new_n259), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n436), .B(new_n440), .C1(new_n442), .C2(new_n268), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n420), .A2(new_n423), .A3(new_n304), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n439), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n307), .A2(new_n359), .A3(new_n415), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n223), .A2(G1698), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(G257), .B2(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n286), .ZN(new_n450));
  INV_X1    g0250(.A(G303), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n289), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n452), .A3(new_n334), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n274), .A2(G1), .ZN(new_n454));
  AND2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  NOR2_X1   g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(KEYINPUT80), .A3(G270), .A4(new_n272), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(G274), .A3(new_n272), .A4(new_n454), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(G270), .A3(new_n272), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT81), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n460), .A4(new_n458), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n453), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n408), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n254), .A2(new_n213), .B1(G20), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n204), .C1(G33), .C2(new_n227), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT20), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n473), .A2(KEYINPUT83), .A3(new_n475), .A4(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n477), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n203), .A2(G33), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n268), .A2(new_n252), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT82), .B1(new_n252), .B2(G116), .ZN(new_n484));
  OR3_X1    g0284(.A1(new_n252), .A2(KEYINPUT82), .A3(G116), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n483), .A2(G116), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n453), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n463), .A2(new_n464), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n461), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(new_n467), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n488), .B1(new_n493), .B2(new_n357), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n470), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n487), .A2(G169), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n496), .B(new_n348), .C1(new_n481), .C2(new_n486), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n469), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(new_n467), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(G179), .A3(new_n453), .A4(new_n487), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n204), .B(G87), .C1(new_n288), .C2(new_n281), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n286), .A2(new_n507), .A3(new_n204), .A4(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G20), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n204), .B2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n222), .A2(KEYINPUT23), .A3(G20), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n509), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n255), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT25), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n252), .B2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n379), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n483), .A2(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n265), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n228), .A2(G1698), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G250), .B2(G1698), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n528), .B2(new_n289), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n334), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n457), .A2(G264), .A3(new_n272), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n408), .A3(new_n460), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G250), .A2(G1698), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n228), .B2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n525), .B1(new_n534), .B2(new_n286), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n460), .B(new_n531), .C1(new_n535), .C2(new_n272), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n532), .A2(KEYINPUT84), .B1(new_n357), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(KEYINPUT84), .A3(new_n357), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n519), .B(new_n523), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n348), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n530), .A2(new_n304), .A3(new_n460), .A4(new_n531), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n509), .A2(new_n516), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n268), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n523), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT85), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n539), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n457), .A2(G257), .A3(new_n272), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n460), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n328), .C1(new_n288), .C2(new_n281), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n328), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n474), .A4(new_n560), .ZN(new_n561));
  AOI211_X1 g0361(.A(new_n304), .B(new_n555), .C1(new_n561), .C2(new_n334), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n334), .ZN(new_n563));
  INV_X1    g0363(.A(new_n555), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n348), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n227), .A2(new_n222), .A3(KEYINPUT6), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n222), .A2(KEYINPUT76), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G107), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n566), .A2(new_n568), .A3(new_n570), .A4(new_n572), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n577));
  OAI21_X1  g0377(.A(G107), .B1(new_n371), .B2(new_n372), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n268), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n379), .A2(new_n227), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n268), .A2(new_n252), .A3(new_n482), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n227), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n562), .A2(new_n565), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  AND4_X1   g0383(.A1(new_n566), .A2(new_n568), .A3(new_n570), .A4(new_n572), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n566), .A2(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n585));
  OAI21_X1  g0385(.A(G20), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n259), .A2(G77), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n578), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n582), .B1(new_n588), .B2(new_n255), .ZN(new_n589));
  AOI211_X1 g0389(.A(G190), .B(new_n555), .C1(new_n561), .C2(new_n334), .ZN(new_n590));
  AOI21_X1  g0390(.A(G200), .B1(new_n563), .B2(new_n564), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(G244), .B(G1698), .C1(new_n288), .C2(new_n281), .ZN(new_n593));
  OAI211_X1 g0393(.A(G238), .B(new_n328), .C1(new_n288), .C2(new_n281), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n511), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n334), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT77), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n272), .A2(new_n597), .A3(G274), .A4(new_n454), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n272), .A2(G274), .A3(new_n454), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n454), .A2(new_n226), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n599), .A2(KEYINPUT77), .B1(new_n600), .B2(new_n272), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  NOR3_X1   g0403(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n604));
  INV_X1    g0404(.A(new_n332), .ZN(new_n605));
  AND2_X1   g0405(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n606));
  NOR2_X1   g0406(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n604), .B1(new_n608), .B2(new_n204), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n204), .B(G68), .C1(new_n288), .C2(new_n281), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n611));
  OR2_X1    g0411(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n612));
  NAND2_X1  g0412(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n255), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n426), .A2(new_n379), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n483), .A2(G87), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n599), .A2(KEYINPUT77), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n600), .A2(new_n272), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n598), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(G190), .A3(new_n596), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n603), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n426), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n483), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n616), .A2(new_n627), .A3(new_n617), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT79), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n623), .A2(new_n304), .A3(new_n596), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n602), .A2(new_n348), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT79), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n616), .A2(new_n627), .A3(new_n632), .A4(new_n617), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n583), .A2(new_n592), .A3(new_n625), .A4(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n447), .A2(new_n504), .A3(new_n553), .A4(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n563), .A2(new_n564), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G169), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n555), .B1(new_n561), .B2(new_n334), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G179), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n589), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT86), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n601), .A2(new_n643), .A3(new_n598), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n642), .A2(new_n644), .B1(new_n334), .B2(new_n595), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n624), .B(new_n619), .C1(new_n645), .C2(new_n357), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n628), .B(new_n630), .C1(new_n645), .C2(G169), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT87), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n641), .A2(new_n625), .A3(new_n634), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(new_n649), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT87), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n654), .A3(new_n649), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n647), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n539), .A2(new_n583), .A3(new_n592), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n646), .A2(new_n647), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n498), .A2(new_n500), .A3(new_n548), .A4(new_n502), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n447), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n413), .A2(new_n414), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n358), .A2(new_n444), .A3(new_n443), .A4(new_n439), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n355), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n403), .A2(new_n406), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n303), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n306), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT88), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(G213), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n488), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n503), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n500), .A2(new_n502), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n683), .B(new_n498), .C1(new_n470), .C2(new_n494), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(new_n681), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n546), .B2(new_n547), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n553), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n548), .B2(new_n680), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n548), .A2(new_n679), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n503), .A2(new_n680), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n553), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n207), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n604), .A2(new_n472), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n211), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n539), .A2(new_n583), .A3(new_n592), .ZN(new_n705));
  INV_X1    g0505(.A(new_n659), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n661), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n647), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n660), .A2(KEYINPUT89), .A3(new_n661), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n703), .B1(new_n714), .B2(new_n680), .ZN(new_n715));
  AOI211_X1 g0515(.A(KEYINPUT29), .B(new_n679), .C1(new_n656), .C2(new_n662), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n530), .A2(new_n453), .A3(G179), .A4(new_n531), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n602), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n501), .A2(new_n720), .A3(new_n639), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n644), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n643), .B1(new_n601), .B2(new_n598), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n596), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n536), .A2(new_n304), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n639), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n469), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n722), .B(new_n555), .C1(new_n561), .C2(new_n334), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n501), .A2(new_n730), .A3(new_n720), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n723), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n732), .B2(new_n679), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n553), .A2(new_n504), .A3(new_n635), .A4(new_n680), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n718), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n717), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n702), .B1(new_n740), .B2(G1), .ZN(G364));
  AND2_X1   g0541(.A1(new_n204), .A2(G13), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n203), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n697), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n686), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n685), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n696), .A2(new_n289), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n748), .A2(G355), .B1(new_n472), .B2(new_n696), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n247), .A2(new_n274), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n207), .A2(new_n289), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G45), .B2(new_n211), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n749), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT91), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n213), .B1(G20), .B2(new_n348), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n745), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n204), .B1(new_n765), .B2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n524), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n204), .A2(new_n408), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n357), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n204), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n765), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G303), .A2(new_n771), .B1(new_n774), .B2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n769), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n775), .B(new_n289), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n408), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n767), .B(new_n778), .C1(G326), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n304), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n772), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT92), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(KEYINPUT92), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n781), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n779), .A2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(KEYINPUT33), .B(G317), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n768), .A2(new_n783), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT95), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n788), .A2(new_n311), .B1(new_n220), .B2(new_n793), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n286), .B1(new_n777), .B2(new_n222), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n774), .A2(G159), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n801));
  INV_X1    g0601(.A(G50), .ZN(new_n802));
  INV_X1    g0602(.A(new_n780), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n799), .B(new_n804), .C1(G87), .C2(new_n771), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n766), .A2(new_n227), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n791), .A2(new_n308), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n800), .C2(new_n801), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n789), .A2(new_n796), .B1(new_n798), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n764), .B1(new_n811), .B2(new_n761), .ZN(new_n812));
  INV_X1    g0612(.A(new_n760), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n763), .B(new_n812), .C1(new_n685), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n747), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  AOI21_X1  g0616(.A(new_n679), .B1(new_n656), .B2(new_n662), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n679), .A2(new_n443), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n438), .A2(new_n445), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT98), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n445), .A2(new_n680), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT98), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n438), .A2(new_n445), .A3(new_n822), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT99), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n820), .A2(KEYINPUT99), .A3(new_n821), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n817), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n820), .A2(new_n823), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n679), .B(new_n831), .C1(new_n656), .C2(new_n662), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT100), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n829), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n738), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT101), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n835), .A2(new_n738), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(KEYINPUT101), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n764), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n761), .A2(new_n758), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n764), .B1(new_n311), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n289), .B1(new_n770), .B2(new_n222), .C1(new_n524), .C2(new_n793), .ZN(new_n843));
  INV_X1    g0643(.A(new_n788), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(G116), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n780), .A2(G303), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n807), .B1(new_n790), .B2(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n777), .A2(new_n225), .B1(new_n773), .B2(new_n782), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT96), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n793), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n851), .A2(G143), .B1(G137), .B2(new_n780), .ZN(new_n852));
  INV_X1    g0652(.A(G159), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n258), .B2(new_n791), .C1(new_n788), .C2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT34), .Z(new_n855));
  INV_X1    g0655(.A(new_n777), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(G68), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n773), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n289), .B(new_n859), .C1(G50), .C2(new_n771), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n220), .B2(new_n766), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n850), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT97), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n761), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(KEYINPUT97), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n842), .B1(new_n759), .B2(new_n824), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n840), .A2(new_n866), .ZN(G384));
  NAND2_X1  g0667(.A1(new_n214), .A2(G116), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n576), .B2(KEYINPUT35), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(KEYINPUT35), .B2(new_n576), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT36), .Z(new_n871));
  OAI211_X1 g0671(.A(new_n212), .B(G77), .C1(new_n220), .C2(new_n308), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n802), .A2(G68), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n203), .B(G13), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n447), .A2(new_n737), .ZN(new_n876));
  INV_X1    g0676(.A(new_n677), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n381), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n402), .A2(new_n411), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n881));
  NAND4_X1  g0681(.A1(new_n402), .A2(new_n411), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT104), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n880), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  INV_X1    g0686(.A(new_n878), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n415), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n415), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n415), .B2(new_n887), .ZN(new_n892));
  INV_X1    g0692(.A(new_n881), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n879), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n882), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n889), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(new_n723), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n728), .A2(new_n726), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n731), .B1(new_n899), .B2(new_n493), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n679), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT31), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n539), .A2(new_n548), .A3(new_n551), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n551), .B1(new_n539), .B2(new_n548), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n635), .B(new_n680), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n903), .B(new_n904), .C1(new_n907), .C2(new_n684), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n679), .A2(new_n321), .A3(new_n323), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n355), .A2(new_n358), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n346), .A2(new_n325), .A3(new_n349), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT72), .B1(new_n351), .B2(new_n353), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(new_n358), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n324), .A3(new_n679), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n916), .A3(new_n824), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n897), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n889), .ZN(new_n924));
  AND2_X1   g0724(.A1(KEYINPUT106), .A2(KEYINPUT40), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n919), .A2(KEYINPUT40), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n876), .B1(new_n927), .B2(new_n718), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT107), .ZN(new_n929));
  INV_X1    g0729(.A(new_n927), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n447), .A2(new_n908), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n404), .A2(new_n405), .A3(new_n381), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n405), .B1(new_n404), .B2(new_n381), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n877), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n445), .A2(new_n679), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n817), .B2(new_n830), .ZN(new_n938));
  INV_X1    g0738(.A(new_n916), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n922), .A2(new_n889), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n897), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n355), .A2(new_n679), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n447), .B1(new_n715), .B2(new_n716), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n670), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n932), .A2(new_n951), .B1(new_n203), .B2(new_n742), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n932), .A2(new_n951), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n875), .B1(new_n952), .B2(new_n953), .ZN(G367));
  NAND2_X1  g0754(.A1(new_n641), .A2(new_n679), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT108), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n583), .B(new_n592), .C1(new_n589), .C2(new_n680), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n693), .A2(new_n553), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n583), .B1(new_n959), .B2(new_n548), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n680), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n680), .A2(new_n619), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(new_n647), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n706), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n962), .A2(new_n964), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n691), .A2(new_n959), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n697), .B(KEYINPUT41), .Z(new_n975));
  OAI21_X1  g0775(.A(new_n960), .B1(new_n689), .B2(new_n693), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n686), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n740), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n694), .A2(new_n958), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT44), .Z(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n982), .B2(new_n690), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n694), .A2(new_n958), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT109), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n690), .A2(new_n982), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n979), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n975), .B1(new_n993), .B2(new_n740), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n974), .B1(new_n994), .B2(new_n744), .ZN(new_n995));
  INV_X1    g0795(.A(new_n752), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n762), .B1(new_n207), .B2(new_n426), .C1(new_n996), .C2(new_n242), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n745), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n844), .A2(G50), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n286), .B1(new_n793), .B2(new_n258), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G159), .B2(new_n790), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n766), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1002), .A2(G68), .B1(G143), .B2(new_n780), .ZN(new_n1003));
  INV_X1    g0803(.A(G137), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n777), .A2(new_n311), .B1(new_n773), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G58), .B2(new_n771), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n844), .A2(G283), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n770), .A2(new_n472), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT46), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G107), .B2(new_n1002), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1009), .A2(KEYINPUT46), .B1(G294), .B2(new_n790), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n289), .B1(new_n777), .B2(new_n227), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G317), .B2(new_n774), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n803), .A2(new_n782), .B1(new_n793), .B2(new_n451), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT111), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n998), .B1(new_n1019), .B2(new_n761), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n966), .A2(new_n967), .A3(new_n760), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n995), .A2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n977), .A2(new_n744), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n748), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1025), .A2(new_n699), .B1(G107), .B2(new_n207), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n430), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n699), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n996), .B1(new_n239), .B2(G45), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1026), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n762), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n745), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT112), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n844), .A2(G68), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n766), .A2(new_n426), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n286), .B1(new_n777), .B2(new_n227), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(G159), .C2(new_n780), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n264), .A2(new_n790), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n802), .A2(new_n793), .B1(new_n770), .B2(new_n311), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G150), .B2(new_n774), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n286), .B1(new_n774), .B2(G326), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n770), .A2(new_n524), .B1(new_n766), .B2(new_n776), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n851), .A2(G317), .B1(G311), .B2(new_n790), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n794), .B2(new_n803), .C1(new_n788), .C2(new_n451), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1044), .B1(new_n472), .B2(new_n777), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n761), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1035), .B(new_n1055), .C1(new_n689), .C2(new_n813), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n978), .A2(new_n697), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n740), .A2(new_n977), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1024), .B(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(G393));
  NAND2_X1  g0859(.A1(new_n959), .A2(new_n760), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n752), .A2(new_n250), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1033), .B1(G97), .B2(new_n696), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n851), .A2(G311), .B1(G317), .B2(new_n780), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n770), .A2(new_n776), .B1(new_n773), .B2(new_n794), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n286), .B(new_n1066), .C1(G107), .C2(new_n856), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n844), .A2(G294), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1002), .A2(G116), .B1(G303), .B2(new_n790), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G143), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n770), .A2(new_n308), .B1(new_n773), .B2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n844), .A2(new_n441), .B1(KEYINPUT113), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n286), .B1(new_n777), .B2(new_n225), .C1(new_n791), .C2(new_n802), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G77), .B2(new_n1002), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(KEYINPUT113), .C2(new_n1072), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n851), .A2(G159), .B1(G150), .B2(new_n780), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1070), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n764), .B(new_n1063), .C1(new_n1079), .C2(new_n761), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1060), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n989), .A2(new_n990), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n989), .A2(new_n990), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1084), .B2(new_n744), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n993), .A2(new_n697), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1084), .A2(new_n979), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(G390));
  NAND3_X1  g0888(.A1(new_n828), .A2(new_n908), .A3(G330), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n939), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n937), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n908), .A2(new_n916), .A3(G330), .A4(new_n824), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n714), .A2(new_n680), .A3(new_n830), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT115), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n916), .B1(new_n737), .B2(new_n824), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n908), .A2(G330), .A3(new_n824), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT115), .A3(new_n939), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n663), .A2(new_n680), .A3(new_n830), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1091), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1094), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n949), .A2(new_n670), .A3(new_n876), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1104), .A2(KEYINPUT116), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT116), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n916), .B1(new_n832), .B2(new_n937), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n945), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n944), .A2(new_n946), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n892), .A2(new_n895), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n891), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT38), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n889), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n939), .B1(new_n1093), .B2(new_n1091), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(KEYINPUT114), .B2(new_n1092), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1092), .A2(KEYINPUT114), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1110), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1109), .B1(new_n938), .B2(new_n939), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n946), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n894), .A2(new_n882), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n665), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n878), .B1(new_n935), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n890), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n921), .B1(new_n1126), .B2(new_n891), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n1127), .B2(new_n889), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1121), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1092), .A2(KEYINPUT114), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1093), .A2(new_n1091), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n916), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n945), .B1(new_n1127), .B2(new_n889), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1118), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1106), .A2(new_n1107), .B1(new_n1120), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n938), .B1(new_n1097), .B2(KEYINPUT115), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1099), .A2(new_n939), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n916), .B1(new_n737), .B2(new_n828), .ZN(new_n1141));
  AND4_X1   g0941(.A1(G330), .A2(new_n908), .A3(new_n916), .A4(new_n824), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1131), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1138), .A2(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n949), .A2(new_n670), .A3(new_n876), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1137), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1119), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1129), .A2(new_n1134), .A3(new_n1118), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1104), .A2(KEYINPUT116), .A3(new_n1105), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1136), .A2(new_n1151), .A3(new_n697), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n841), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n791), .A2(new_n1004), .B1(new_n793), .B2(new_n858), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n770), .A2(new_n258), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n803), .C1(new_n853), .C2(new_n766), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1154), .B(new_n1158), .C1(new_n844), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n286), .B1(new_n773), .B2(new_n1162), .C1(new_n802), .C2(new_n777), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n289), .B1(new_n770), .B2(new_n225), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n791), .A2(new_n222), .B1(new_n803), .B2(new_n776), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G77), .C2(new_n1002), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n857), .B1(new_n472), .B2(new_n793), .C1(new_n524), .C2(new_n773), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G97), .B2(new_n844), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1161), .A2(new_n1164), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n761), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n745), .B1(new_n264), .B2(new_n1153), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n944), .A2(new_n946), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n758), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n744), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1152), .A2(KEYINPUT118), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT118), .B1(new_n1152), .B2(new_n1176), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(G378));
  NAND2_X1  g0979(.A1(new_n877), .A2(new_n269), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT121), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n307), .B(new_n1181), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  XOR2_X1   g0983(.A(new_n1182), .B(new_n1183), .Z(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n927), .B2(new_n718), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1182), .B(new_n1183), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n924), .A2(new_n926), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n923), .B1(new_n897), .B2(new_n918), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(G330), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n948), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1185), .A2(new_n948), .A3(new_n1190), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n744), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n745), .B1(G50), .B2(new_n1153), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n289), .A2(new_n273), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n802), .C1(G33), .C2(G41), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n770), .A2(new_n311), .B1(new_n773), .B2(new_n776), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n791), .A2(new_n227), .B1(new_n803), .B2(new_n472), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G68), .C2(new_n1002), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n777), .A2(new_n220), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1197), .B(new_n1202), .C1(G107), .C2(new_n851), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n426), .C2(new_n788), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT58), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1205), .B2(new_n1204), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n788), .A2(new_n1004), .B1(new_n858), .B2(new_n791), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT119), .Z(new_n1209));
  OAI22_X1  g1009(.A1(new_n1157), .A2(new_n793), .B1(new_n770), .B2(new_n1159), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G150), .B2(new_n1002), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(new_n1162), .C2(new_n803), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n265), .B(new_n273), .C1(new_n777), .C2(new_n853), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G124), .B2(new_n774), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT59), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1207), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1196), .B1(new_n1220), .B2(new_n761), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1184), .B2(new_n759), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1195), .A2(KEYINPUT122), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT122), .B1(new_n1195), .B2(new_n1222), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1136), .A2(new_n1105), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1185), .A2(new_n948), .A3(new_n1190), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n948), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1229), .A3(KEYINPUT57), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n697), .B(new_n1230), .C1(new_n1231), .C2(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(KEYINPUT123), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1225), .B1(new_n1232), .B2(new_n1236), .ZN(G375));
  NOR2_X1   g1037(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n975), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT124), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n764), .B1(new_n308), .B2(new_n841), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n289), .B(new_n1202), .C1(G50), .C2(new_n1002), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1160), .A2(new_n790), .B1(G132), .B2(new_n780), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G159), .A2(new_n771), .B1(new_n774), .B2(G128), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n1004), .B2(new_n793), .C1(new_n788), .C2(new_n258), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G97), .A2(new_n771), .B1(new_n774), .B2(G303), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n776), .B2(new_n793), .C1(new_n788), .C2(new_n222), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n791), .A2(new_n472), .B1(new_n803), .B2(new_n524), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n289), .B1(new_n777), .B2(new_n311), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1252), .A2(new_n1037), .A3(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1247), .A2(new_n1249), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(KEYINPUT125), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n761), .B1(new_n1256), .B2(KEYINPUT125), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1244), .B1(new_n1257), .B2(new_n1258), .C1(new_n916), .C2(new_n759), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1145), .B2(new_n743), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1243), .A2(new_n1261), .ZN(G381));
  OR3_X1    g1062(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1152), .A2(new_n1176), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(G387), .A2(new_n1263), .A3(G390), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G375), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1261), .A4(new_n1243), .ZN(G407));
  NAND2_X1  g1068(.A1(new_n678), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1264), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(G213), .A3(new_n1271), .ZN(G409));
  XNOR2_X1  g1072(.A(G393), .B(new_n815), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n995), .A2(new_n1022), .A3(G390), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G390), .B1(new_n995), .B2(new_n1022), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1081), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n991), .A2(new_n992), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n743), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n978), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(new_n698), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n978), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1273), .A3(new_n1275), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1278), .A2(new_n1279), .A3(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1225), .C1(new_n1232), .C2(new_n1236), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1233), .A2(new_n975), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1195), .A2(new_n1222), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1264), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1240), .A2(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n697), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1238), .A2(KEYINPUT60), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1241), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(G384), .A3(new_n1261), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n866), .B(new_n840), .C1(new_n1298), .C2(new_n1260), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1294), .A2(new_n1269), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1289), .B1(new_n1305), .B2(KEYINPUT63), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1294), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1290), .A2(KEYINPUT126), .A3(new_n1293), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1308), .A2(new_n1269), .A3(new_n1309), .A4(new_n1303), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1308), .A2(new_n1313), .A3(new_n1269), .A4(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1270), .A2(G2897), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1302), .B(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1270), .B1(new_n1294), .B2(new_n1307), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1313), .B1(new_n1318), .B2(new_n1309), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1306), .B(new_n1312), .C1(new_n1317), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1278), .A2(new_n1288), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1294), .A2(new_n1269), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1316), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1321), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1327), .ZN(G405));
  NOR2_X1   g1128(.A1(new_n1267), .A2(new_n1265), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1290), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1303), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1290), .B(new_n1302), .C1(new_n1267), .C2(new_n1265), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1321), .ZN(G402));
endmodule


