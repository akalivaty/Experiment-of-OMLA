

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591;

  XNOR2_X1 U320 ( .A(n465), .B(KEYINPUT47), .ZN(n466) );
  INV_X1 U321 ( .A(KEYINPUT121), .ZN(n480) );
  XNOR2_X1 U322 ( .A(n467), .B(n466), .ZN(n473) );
  XNOR2_X1 U323 ( .A(n480), .B(KEYINPUT55), .ZN(n481) );
  AND2_X1 U324 ( .A1(G226GAT), .A2(G233GAT), .ZN(n288) );
  INV_X1 U325 ( .A(KEYINPUT96), .ZN(n398) );
  XNOR2_X1 U326 ( .A(n398), .B(KEYINPUT27), .ZN(n399) );
  XNOR2_X1 U327 ( .A(n397), .B(n399), .ZN(n439) );
  XNOR2_X1 U328 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n476) );
  XNOR2_X1 U329 ( .A(n392), .B(n288), .ZN(n393) );
  INV_X1 U330 ( .A(KEYINPUT19), .ZN(n289) );
  XNOR2_X1 U331 ( .A(n477), .B(n476), .ZN(n572) );
  XNOR2_X1 U332 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n389) );
  XOR2_X1 U336 ( .A(n346), .B(n345), .Z(n580) );
  INV_X1 U337 ( .A(G99GAT), .ZN(n451) );
  XNOR2_X1 U338 ( .A(KEYINPUT38), .B(n456), .ZN(n507) );
  XNOR2_X1 U339 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U340 ( .A(n451), .B(KEYINPUT112), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n457), .B(G43GAT), .ZN(n458) );
  XNOR2_X1 U342 ( .A(n487), .B(n486), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n453), .B(n452), .ZN(G1338GAT) );
  XNOR2_X1 U344 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n290) );
  XOR2_X1 U345 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n291) );
  XOR2_X1 U346 ( .A(G190GAT), .B(G99GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U349 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n296) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G176GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n304) );
  XOR2_X1 U353 ( .A(G127GAT), .B(KEYINPUT0), .Z(n300) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n405) );
  XOR2_X1 U356 ( .A(G120GAT), .B(G71GAT), .Z(n341) );
  XOR2_X1 U357 ( .A(n405), .B(n341), .Z(n302) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U361 ( .A(n389), .B(n305), .Z(n517) );
  INV_X1 U362 ( .A(n517), .ZN(n539) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n306), .B(G29GAT), .ZN(n307) );
  XOR2_X1 U365 ( .A(n307), .B(KEYINPUT8), .Z(n309) );
  XNOR2_X1 U366 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n382) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G1GAT), .Z(n351) );
  XOR2_X1 U369 ( .A(KEYINPUT73), .B(KEYINPUT68), .Z(n311) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G197GAT), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n351), .B(n312), .ZN(n314) );
  AND2_X1 U373 ( .A1(G229GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U375 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n316) );
  XNOR2_X1 U376 ( .A(KEYINPUT29), .B(KEYINPUT70), .ZN(n315) );
  XOR2_X1 U377 ( .A(n316), .B(n315), .Z(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n322) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(G22GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n319), .B(G141GAT), .ZN(n422) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G36GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(G8GAT), .ZN(n386) );
  XNOR2_X1 U383 ( .A(n422), .B(n386), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U385 ( .A(n382), .B(n323), .Z(n575) );
  INV_X1 U386 ( .A(G92GAT), .ZN(n324) );
  NAND2_X1 U387 ( .A1(G64GAT), .A2(n324), .ZN(n327) );
  INV_X1 U388 ( .A(G64GAT), .ZN(n325) );
  NAND2_X1 U389 ( .A1(n325), .A2(G92GAT), .ZN(n326) );
  NAND2_X1 U390 ( .A1(n327), .A2(n326), .ZN(n331) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n385) );
  XNOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n328), .B(KEYINPUT75), .ZN(n355) );
  INV_X1 U395 ( .A(n355), .ZN(n329) );
  NAND2_X1 U396 ( .A1(n385), .A2(n329), .ZN(n334) );
  XOR2_X1 U397 ( .A(n331), .B(n330), .Z(n332) );
  NAND2_X1 U398 ( .A1(n332), .A2(n355), .ZN(n333) );
  NAND2_X1 U399 ( .A1(n334), .A2(n333), .ZN(n338) );
  XNOR2_X1 U400 ( .A(G106GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n335), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n336), .B(KEYINPUT76), .ZN(n372) );
  XNOR2_X1 U404 ( .A(n429), .B(n372), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n340) );
  XNOR2_X1 U407 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n340), .B(n339), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n344) );
  AND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n580), .B(KEYINPUT41), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n347), .B(KEYINPUT64), .ZN(n460) );
  XNOR2_X1 U414 ( .A(n460), .B(KEYINPUT105), .ZN(n543) );
  NAND2_X1 U415 ( .A1(n575), .A2(n543), .ZN(n511) );
  XOR2_X1 U416 ( .A(G127GAT), .B(G71GAT), .Z(n349) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(G183GAT), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U419 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U420 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U422 ( .A(n354), .B(KEYINPUT83), .Z(n357) );
  XNOR2_X1 U423 ( .A(G8GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U425 ( .A(G64GAT), .B(G78GAT), .Z(n359) );
  XNOR2_X1 U426 ( .A(G155GAT), .B(G211GAT), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n361) );
  XNOR2_X1 U429 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U431 ( .A(n363), .B(n362), .Z(n364) );
  XOR2_X1 U432 ( .A(n365), .B(n364), .Z(n557) );
  XOR2_X1 U433 ( .A(G190GAT), .B(KEYINPUT81), .Z(n392) );
  XOR2_X1 U434 ( .A(KEYINPUT79), .B(G92GAT), .Z(n367) );
  XNOR2_X1 U435 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U437 ( .A(n392), .B(n368), .Z(n370) );
  NAND2_X1 U438 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U439 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U440 ( .A(n371), .B(KEYINPUT9), .Z(n374) );
  XNOR2_X1 U441 ( .A(G50GAT), .B(n372), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U443 ( .A(KEYINPUT80), .B(G106GAT), .Z(n376) );
  XNOR2_X1 U444 ( .A(G134GAT), .B(G162GAT), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U447 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n380) );
  XNOR2_X1 U448 ( .A(G36GAT), .B(KEYINPUT66), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n384), .B(n383), .ZN(n560) );
  XNOR2_X1 U452 ( .A(n560), .B(KEYINPUT36), .ZN(n589) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n391) );
  XOR2_X1 U455 ( .A(G211GAT), .B(KEYINPUT21), .Z(n388) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(G218GAT), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n388), .B(n387), .ZN(n430) );
  XNOR2_X1 U458 ( .A(n389), .B(n430), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n394) );
  XOR2_X1 U460 ( .A(n396), .B(n395), .Z(n397) );
  XOR2_X1 U461 ( .A(KEYINPUT93), .B(KEYINPUT90), .Z(n401) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U464 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n407) );
  XOR2_X1 U465 ( .A(KEYINPUT3), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U466 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U468 ( .A(KEYINPUT2), .B(n404), .Z(n433) );
  XNOR2_X1 U469 ( .A(n405), .B(n433), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n421) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XOR2_X1 U473 ( .A(G57GAT), .B(G148GAT), .Z(n411) );
  XNOR2_X1 U474 ( .A(G141GAT), .B(G120GAT), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U476 ( .A(G29GAT), .B(G85GAT), .Z(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n417) );
  XNOR2_X1 U480 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U483 ( .A(n421), .B(n420), .Z(n525) );
  NAND2_X1 U484 ( .A1(n439), .A2(n525), .ZN(n534) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(n422), .Z(n424) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U488 ( .A(G204GAT), .B(KEYINPUT23), .Z(n426) );
  XNOR2_X1 U489 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U491 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U494 ( .A(n434), .B(n433), .Z(n478) );
  XNOR2_X1 U495 ( .A(n478), .B(KEYINPUT67), .ZN(n435) );
  XOR2_X1 U496 ( .A(n435), .B(KEYINPUT28), .Z(n520) );
  INV_X1 U497 ( .A(n520), .ZN(n537) );
  NAND2_X1 U498 ( .A1(n537), .A2(n539), .ZN(n436) );
  NOR2_X1 U499 ( .A1(n534), .A2(n436), .ZN(n447) );
  XOR2_X1 U500 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n438) );
  NAND2_X1 U501 ( .A1(n478), .A2(n539), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n574) );
  INV_X1 U503 ( .A(n574), .ZN(n552) );
  NAND2_X1 U504 ( .A1(n439), .A2(n552), .ZN(n440) );
  XOR2_X1 U505 ( .A(KEYINPUT98), .B(n440), .Z(n444) );
  NOR2_X1 U506 ( .A1(n539), .A2(n397), .ZN(n441) );
  NOR2_X1 U507 ( .A1(n478), .A2(n441), .ZN(n442) );
  XOR2_X1 U508 ( .A(KEYINPUT25), .B(n442), .Z(n443) );
  NOR2_X1 U509 ( .A1(n444), .A2(n443), .ZN(n445) );
  NOR2_X1 U510 ( .A1(n445), .A2(n525), .ZN(n446) );
  NOR2_X1 U511 ( .A1(n447), .A2(n446), .ZN(n491) );
  NOR2_X1 U512 ( .A1(n589), .A2(n491), .ZN(n448) );
  NAND2_X1 U513 ( .A1(n557), .A2(n448), .ZN(n449) );
  XOR2_X1 U514 ( .A(KEYINPUT37), .B(n449), .Z(n455) );
  NOR2_X1 U515 ( .A1(n511), .A2(n455), .ZN(n450) );
  XNOR2_X1 U516 ( .A(n450), .B(KEYINPUT109), .ZN(n530) );
  NOR2_X1 U517 ( .A1(n539), .A2(n530), .ZN(n453) );
  XOR2_X1 U518 ( .A(KEYINPUT74), .B(n575), .Z(n562) );
  INV_X1 U519 ( .A(n562), .ZN(n470) );
  NOR2_X1 U520 ( .A1(n580), .A2(n470), .ZN(n454) );
  XOR2_X1 U521 ( .A(KEYINPUT78), .B(n454), .Z(n493) );
  NOR2_X1 U522 ( .A1(n493), .A2(n455), .ZN(n456) );
  NAND2_X1 U523 ( .A1(n517), .A2(n507), .ZN(n459) );
  XOR2_X1 U524 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n457) );
  XNOR2_X1 U525 ( .A(n459), .B(n458), .ZN(G1330GAT) );
  INV_X1 U526 ( .A(n560), .ZN(n565) );
  INV_X1 U527 ( .A(n557), .ZN(n584) );
  NOR2_X1 U528 ( .A1(n575), .A2(n460), .ZN(n461) );
  XNOR2_X1 U529 ( .A(n461), .B(KEYINPUT46), .ZN(n462) );
  NOR2_X1 U530 ( .A1(n584), .A2(n462), .ZN(n463) );
  XOR2_X1 U531 ( .A(KEYINPUT114), .B(n463), .Z(n464) );
  NOR2_X1 U532 ( .A1(n565), .A2(n464), .ZN(n467) );
  INV_X1 U533 ( .A(KEYINPUT115), .ZN(n465) );
  NOR2_X1 U534 ( .A1(n557), .A2(n589), .ZN(n468) );
  XOR2_X1 U535 ( .A(KEYINPUT45), .B(n468), .Z(n469) );
  NOR2_X1 U536 ( .A1(n580), .A2(n469), .ZN(n471) );
  NAND2_X1 U537 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U538 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U539 ( .A(n474), .B(KEYINPUT48), .Z(n535) );
  XOR2_X1 U540 ( .A(n397), .B(KEYINPUT119), .Z(n475) );
  NOR2_X1 U541 ( .A1(n535), .A2(n475), .ZN(n477) );
  NOR2_X1 U542 ( .A1(n478), .A2(n525), .ZN(n479) );
  AND2_X1 U543 ( .A1(n572), .A2(n479), .ZN(n482) );
  NOR2_X1 U544 ( .A1(n539), .A2(n483), .ZN(n566) );
  NAND2_X1 U545 ( .A1(n566), .A2(n543), .ZN(n487) );
  XOR2_X1 U546 ( .A(G176GAT), .B(KEYINPUT122), .Z(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n484) );
  NAND2_X1 U548 ( .A1(n584), .A2(n560), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT84), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT16), .ZN(n490) );
  NOR2_X1 U551 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT99), .B(n492), .ZN(n510) );
  NOR2_X1 U553 ( .A1(n493), .A2(n510), .ZN(n500) );
  NAND2_X1 U554 ( .A1(n525), .A2(n500), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(KEYINPUT34), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  INV_X1 U557 ( .A(n397), .ZN(n514) );
  NAND2_X1 U558 ( .A1(n500), .A2(n514), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT100), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G8GAT), .B(n497), .ZN(G1325GAT) );
  XOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U562 ( .A1(n500), .A2(n517), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  XOR2_X1 U564 ( .A(G22GAT), .B(KEYINPUT101), .Z(n502) );
  NAND2_X1 U565 ( .A1(n500), .A2(n520), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1327GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U568 ( .A1(n507), .A2(n525), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U571 ( .A1(n507), .A2(n514), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(KEYINPUT104), .ZN(n509) );
  NAND2_X1 U574 ( .A1(n520), .A2(n507), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  NOR2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n525), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n521), .A2(n514), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(KEYINPUT106), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  XOR2_X1 U583 ( .A(G71GAT), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U584 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  INV_X1 U590 ( .A(n525), .ZN(n571) );
  NOR2_X1 U591 ( .A1(n571), .A2(n530), .ZN(n527) );
  XNOR2_X1 U592 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n397), .ZN(n529) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n537), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n541) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(KEYINPUT116), .B(n536), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n537), .A2(n551), .ZN(n538) );
  NOR2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n548), .A2(n562), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U610 ( .A1(n548), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NAND2_X1 U612 ( .A1(n584), .A2(n548), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n565), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n559) );
  NOR2_X1 U619 ( .A1(n575), .A2(n559), .ZN(n553) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U621 ( .A1(n460), .A2(n559), .ZN(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n559), .ZN(n558) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n566), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n584), .A2(n566), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .Z(n577) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n583) );
  INV_X1 U641 ( .A(n583), .ZN(n588) );
  OR2_X1 U642 ( .A1(n588), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n587) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U655 ( .A(n591), .B(n590), .Z(G1355GAT) );
endmodule

