//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(KEYINPUT65), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(KEYINPUT65), .B2(new_n458), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n470), .A2(new_n473), .A3(new_n464), .A4(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT68), .Z(G160));
  INV_X1    g056(.A(new_n475), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(G112), .B2(new_n464), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n470), .A2(new_n473), .A3(G2105), .A4(new_n474), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n483), .B(new_n487), .C1(G124), .C2(new_n489), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n464), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n488), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n469), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(KEYINPUT70), .A3(new_n470), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n470), .A2(new_n473), .A3(new_n474), .A4(new_n499), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n500), .A2(KEYINPUT4), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n474), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n464), .A3(G138), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT71), .B1(new_n465), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n494), .B1(new_n504), .B2(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(new_n519), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n526), .A2(G62), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT73), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(new_n529), .A3(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND2_X1  g111(.A1(new_n528), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n524), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n540), .A2(new_n541), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(new_n528), .A2(G90), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n520), .A2(new_n521), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(G52), .A3(G543), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(new_n530), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n548), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n524), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n528), .A2(G81), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n550), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND4_X1  g140(.A1(new_n547), .A2(KEYINPUT75), .A3(G91), .A4(new_n526), .ZN(new_n566));
  OAI211_X1 g141(.A(G91), .B(new_n526), .C1(new_n520), .C2(new_n521), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n527), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n566), .A2(new_n569), .B1(G651), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  OAI211_X1 g149(.A(G53), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n573), .B2(new_n576), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G299));
  OAI21_X1  g155(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n528), .B2(G87), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n547), .A2(G49), .A3(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  AND2_X1   g160(.A1(KEYINPUT5), .A2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(KEYINPUT5), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G61), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n588), .A2(new_n589), .B1(G73), .B2(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n526), .A2(KEYINPUT77), .A3(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n550), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(G48), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n593));
  OAI211_X1 g168(.A(G86), .B(new_n526), .C1(new_n520), .C2(new_n521), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n550), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(G47), .A2(new_n524), .B1(new_n528), .B2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  OR3_X1    g183(.A1(G171), .A2(KEYINPUT80), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(G171), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n524), .A2(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(new_n516), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n547), .A2(new_n526), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n620), .ZN(G284));
  OAI211_X1 g196(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n620), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n608), .ZN(new_n623));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT81), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(G297));
  XOR2_X1   g201(.A(G297), .B(KEYINPUT82), .Z(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n620), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n559), .A2(new_n608), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n618), .A2(new_n619), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(new_n611), .A3(new_n613), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n630), .B1(new_n633), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n465), .A2(new_n478), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n488), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n482), .B2(G135), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n655), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n664), .A3(G14), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n667), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT86), .Z(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G5), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G171), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G1961), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(G21), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G168), .B2(new_n699), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G1966), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(G1961), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1341), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n560), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G16), .B2(G19), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n702), .B(new_n707), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G4), .A2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT89), .Z(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n632), .B2(new_n699), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1348), .ZN(new_n715));
  NOR2_X1   g290(.A1(G29), .A2(G35), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G162), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n711), .B(new_n715), .C1(G2090), .C2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n722));
  INV_X1    g297(.A(G140), .ZN(new_n723));
  INV_X1    g298(.A(G128), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n722), .B1(new_n475), .B2(new_n723), .C1(new_n724), .C2(new_n488), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT91), .Z(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G26), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  OAI22_X1  g308(.A1(new_n710), .A2(new_n708), .B1(G1966), .B2(new_n704), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n729), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT25), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(new_n464), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n737), .B(new_n739), .C1(G139), .C2(new_n482), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(new_n729), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(G2072), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n746), .A2(new_n745), .A3(G28), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n745), .B2(G28), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n729), .B1(new_n745), .B2(G28), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n744), .B(new_n749), .C1(new_n645), .C2(new_n729), .ZN(new_n750));
  NOR4_X1   g325(.A1(new_n734), .A2(new_n742), .A3(new_n743), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G160), .A2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(new_n753), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2084), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n729), .A2(G32), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT26), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(new_n478), .B2(G105), .ZN(new_n763));
  INV_X1    g338(.A(G129), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n488), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n482), .B2(G141), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n758), .B1(new_n768), .B2(new_n729), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT27), .B(G1996), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n769), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n729), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n729), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n751), .A2(new_n757), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n720), .A2(new_n733), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G299), .A2(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n699), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G1956), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G2090), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n784), .A2(KEYINPUT96), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n778), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n699), .A2(G23), .ZN(new_n791));
  INV_X1    g366(.A(G288), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n699), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n699), .A2(G22), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n699), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G6), .A2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n596), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n795), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n699), .A2(G24), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G290), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1986), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n795), .A2(new_n799), .A3(new_n809), .A4(new_n803), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n729), .A2(G25), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n482), .A2(G131), .ZN(new_n812));
  INV_X1    g387(.A(G119), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n464), .A2(G107), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n488), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n817), .B2(new_n729), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  NAND3_X1  g395(.A1(new_n808), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT87), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(KEYINPUT87), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n805), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(KEYINPUT88), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n821), .B(KEYINPUT87), .ZN(new_n829));
  INV_X1    g404(.A(new_n827), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n829), .A2(new_n805), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n790), .B1(new_n828), .B2(new_n831), .ZN(G311));
  INV_X1    g407(.A(new_n790), .ZN(new_n833));
  INV_X1    g408(.A(new_n831), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n830), .B1(new_n829), .B2(new_n805), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(G150));
  NOR2_X1   g411(.A1(new_n632), .A2(new_n628), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n528), .A2(G93), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n524), .A2(G55), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(new_n550), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n559), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n559), .A2(new_n843), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n838), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT97), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n767), .A2(new_n740), .ZN(new_n855));
  INV_X1    g430(.A(new_n766), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n740), .ZN(new_n857));
  INV_X1    g432(.A(new_n503), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT4), .B1(new_n501), .B2(new_n502), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n513), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n494), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n726), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n489), .A2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n464), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n482), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n637), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n817), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G160), .B(new_n645), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n864), .A2(new_n874), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n881), .B(new_n875), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n873), .A2(KEYINPUT98), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n879), .B(new_n880), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g462(.A(G288), .B1(new_n604), .B2(new_n606), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g465(.A1(G166), .A2(new_n596), .ZN(new_n891));
  NAND2_X1  g466(.A1(G305), .A2(G303), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n604), .A2(G288), .A3(new_n606), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n890), .A3(new_n892), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n893), .B1(new_n898), .B2(new_n888), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT42), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n578), .A2(new_n632), .A3(new_n579), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n573), .A2(new_n576), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT76), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n620), .B1(new_n904), .B2(new_n577), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT99), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n902), .B2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n846), .B(new_n633), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n902), .B2(new_n905), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n632), .B1(new_n578), .B2(new_n579), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n904), .A2(new_n577), .A3(new_n620), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(new_n911), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n901), .A2(new_n912), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n901), .B1(new_n912), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n843), .A2(new_n608), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(G331));
  XNOR2_X1  g500(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g502(.A1(G301), .A2(KEYINPUT102), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n546), .A2(new_n548), .A3(new_n929), .A4(new_n551), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(G168), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G168), .B1(new_n928), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n846), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G286), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n559), .B(new_n843), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n931), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(new_n906), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n944), .B2(new_n918), .ZN(new_n945));
  INV_X1    g520(.A(new_n900), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n934), .A2(KEYINPUT103), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT103), .B1(new_n934), .B2(new_n938), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n918), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n940), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n900), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n927), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n946), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n880), .ZN(new_n956));
  OAI211_X1 g531(.A(KEYINPUT104), .B(new_n913), .C1(new_n902), .C2(new_n905), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n939), .B(new_n957), .C1(new_n918), .C2(KEYINPUT104), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n942), .A2(new_n907), .A3(new_n909), .A4(new_n943), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n946), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n956), .A2(new_n960), .A3(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n926), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n947), .A2(new_n927), .A3(new_n953), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n956), .B2(new_n960), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(G397));
  AOI21_X1  g541(.A(G1384), .B1(new_n860), .B2(new_n861), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR4_X1   g546(.A1(new_n468), .A2(new_n477), .A3(new_n971), .A4(new_n479), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1996), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n768), .ZN(new_n977));
  INV_X1    g552(.A(G2067), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n726), .B(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT108), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n973), .B1(new_n980), .B2(new_n766), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n979), .B(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(G1996), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n973), .ZN(new_n985));
  INV_X1    g560(.A(new_n817), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n986), .A2(new_n819), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n819), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n991));
  NAND2_X1  g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(new_n985), .C1(new_n991), .C2(new_n992), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n977), .A2(new_n984), .A3(new_n989), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(G1976), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n590), .A2(new_n591), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n530), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n999), .A2(new_n1000), .B1(new_n592), .B2(new_n595), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  INV_X1    g577(.A(new_n595), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n530), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n997), .A4(G1981), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1001), .A2(KEYINPUT115), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n967), .B2(new_n972), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1000), .B1(new_n1004), .B2(KEYINPUT114), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n596), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1002), .B1(new_n1012), .B2(new_n1001), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n996), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n596), .A2(new_n1000), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(KEYINPUT116), .A3(new_n1015), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n1008), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n1021));
  AND3_X1   g596(.A1(G303), .A2(G8), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n1023));
  AOI22_X1  g598(.A1(G303), .A2(G8), .B1(new_n1023), .B2(KEYINPUT55), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n968), .B1(G164), .B2(G1384), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n507), .B1(new_n506), .B2(new_n509), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n465), .A2(KEYINPUT71), .A3(new_n511), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AND4_X1   g605(.A1(new_n470), .A2(new_n473), .A3(new_n474), .A4(new_n499), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n508), .B1(new_n1031), .B2(KEYINPUT70), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1032), .B2(new_n503), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT45), .B(new_n1027), .C1(new_n1033), .C2(new_n494), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1026), .A2(new_n972), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n798), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1027), .B1(new_n1033), .B2(new_n494), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1039));
  NAND2_X1  g614(.A1(new_n967), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .A4(new_n972), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1007), .B(new_n1025), .C1(new_n1036), .C2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n972), .B1(new_n967), .B2(new_n1039), .ZN(new_n1044));
  NOR3_X1   g619(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1046), .A2(new_n1041), .B1(new_n1035), .B2(new_n798), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1025), .B1(new_n1047), .B2(new_n1007), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G168), .A2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(G1966), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1027), .B(new_n969), .C1(new_n1033), .C2(new_n494), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n972), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G2084), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1038), .A2(new_n1040), .A3(new_n1055), .A4(new_n972), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT63), .B(new_n1049), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1043), .B1(new_n1048), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n862), .A2(new_n1027), .A3(new_n972), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n547), .A2(G87), .A3(new_n526), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n584), .A2(new_n1060), .A3(G1976), .A4(new_n581), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n583), .A2(KEYINPUT111), .A3(G1976), .A4(new_n584), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1059), .A2(G8), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT112), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1068), .A3(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1001), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT49), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n1008), .A3(new_n1006), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT113), .B(G1976), .Z(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1008), .A2(new_n1075), .A3(new_n1064), .A4(new_n1063), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1067), .A2(new_n1069), .A3(new_n1073), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1020), .B1(new_n1058), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1007), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1025), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(G8), .A3(G168), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1077), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1079), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1078), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n783), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n573), .A2(new_n1092), .A3(new_n576), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n573), .B2(new_n576), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1026), .A2(new_n1034), .A3(new_n972), .A4(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n1099));
  INV_X1    g674(.A(new_n972), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1039), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1037), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n967), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1956), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1097), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1099), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1091), .A2(KEYINPUT118), .A3(new_n1097), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1094), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n573), .A2(new_n1092), .A3(new_n576), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT119), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n1108), .A4(new_n1114), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1038), .A2(new_n972), .A3(new_n1040), .ZN(new_n1119));
  INV_X1    g694(.A(G1348), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n967), .A2(new_n978), .A3(new_n972), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n620), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1117), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT121), .B(G1996), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1026), .A2(new_n1034), .A3(new_n972), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1059), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n560), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1133), .A3(new_n560), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1091), .A2(new_n1136), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1095), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1098), .B1(new_n1138), .B2(KEYINPUT61), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n620), .B(KEYINPUT122), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1141), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n1122), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1123), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1123), .A2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n632), .A2(KEYINPUT122), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1142), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1098), .A2(new_n1125), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1054), .A2(G168), .A3(new_n1056), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT124), .B1(new_n1149), .B2(G8), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT51), .B1(new_n1150), .B2(KEYINPUT123), .ZN(new_n1151));
  NOR2_X1   g726(.A1(G286), .A2(KEYINPUT124), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1153));
  NOR2_X1   g728(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1154));
  OAI211_X1 g729(.A(G8), .B(new_n1149), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(G2078), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1026), .A2(new_n1034), .A3(new_n972), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1100), .B1(new_n1037), .B2(new_n968), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(KEYINPUT126), .A3(new_n1034), .A4(new_n1158), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT125), .B(G1961), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1119), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1026), .A2(new_n1034), .A3(new_n775), .A4(new_n972), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1157), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(G171), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1100), .B1(new_n967), .B2(new_n969), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1171), .B(new_n1158), .C1(KEYINPUT45), .C2(new_n967), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1166), .A2(new_n1172), .A3(new_n1168), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1170), .B(KEYINPUT54), .C1(G171), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1046), .A2(new_n1041), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1036), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1083), .B1(new_n1176), .B2(G8), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1177), .A2(new_n1077), .A3(new_n1043), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1179), .A2(G301), .A3(new_n1168), .A4(new_n1166), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1173), .A2(G171), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1156), .A2(new_n1174), .A3(new_n1178), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1090), .B1(new_n1148), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1156), .A2(KEYINPUT62), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1178), .A2(G171), .A3(new_n1173), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1189), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n995), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n990), .A2(new_n973), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT48), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n984), .A2(new_n977), .A3(new_n989), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n985), .B1(new_n983), .B2(new_n856), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n974), .B(KEYINPUT107), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT46), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT46), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1197), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1202), .A2(KEYINPUT47), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(KEYINPUT47), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n984), .A2(new_n977), .A3(new_n988), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n726), .A2(G2067), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n973), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1192), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n462), .A2(G227), .ZN(new_n1213));
  AND3_X1   g787(.A1(new_n665), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1212), .B1(new_n665), .B2(new_n1213), .ZN(new_n1215));
  NOR3_X1   g789(.A1(new_n1214), .A2(new_n1215), .A3(G229), .ZN(new_n1216));
  OAI211_X1 g790(.A(new_n886), .B(new_n1216), .C1(new_n954), .C2(new_n961), .ZN(G225));
  INV_X1    g791(.A(G225), .ZN(G308));
endmodule


