//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(new_n206), .A2(KEYINPUT0), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n212), .B1(KEYINPUT0), .B2(new_n206), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n214), .A2(new_n222), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(G226), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT67), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n228), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G20), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n208), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n244), .B1(new_n245), .B2(new_n246), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT72), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT72), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n253), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n207), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n252), .A2(new_n254), .A3(new_n207), .A4(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G68), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT11), .B1(new_n250), .B2(new_n255), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n258), .A2(G68), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT14), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G226), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G238), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G41), .A2(G45), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT70), .B1(new_n287), .B2(G1), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n289), .B(new_n257), .C1(G41), .C2(G45), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n288), .A2(G274), .A3(new_n283), .A4(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n281), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n281), .B2(new_n292), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n269), .B(G169), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n281), .A2(new_n292), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT13), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n281), .A2(new_n292), .A3(new_n293), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(G179), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n299), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n269), .B1(new_n302), .B2(G169), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n268), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n305), .B(new_n267), .C1(new_n306), .C2(new_n302), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n285), .A2(G226), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n310), .A2(new_n291), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT71), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n274), .A2(G222), .A3(new_n276), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n274), .A2(G1698), .ZN(new_n315));
  INV_X1    g0115(.A(G223), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n314), .B1(new_n246), .B2(new_n274), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n280), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n260), .A2(G50), .A3(new_n261), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  INV_X1    g0123(.A(G150), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n245), .B1(new_n324), .B2(new_n248), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G50), .A2(G58), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n208), .B1(new_n326), .B2(new_n243), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n255), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n322), .B(new_n328), .C1(G50), .C2(new_n258), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n312), .A2(new_n330), .A3(new_n313), .A4(new_n318), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n321), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n319), .A2(G200), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n329), .B(KEYINPUT9), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n312), .A2(G190), .A3(new_n313), .A4(new_n318), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT10), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT10), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .A4(new_n336), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n333), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n291), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  OAI211_X1 g0146(.A(G223), .B(new_n276), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(G226), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G87), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n280), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n344), .A2(new_n351), .A3(new_n306), .ZN(new_n352));
  AOI21_X1  g0152(.A(G200), .B1(new_n344), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT8), .B(G58), .Z(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n261), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n356), .A2(new_n259), .B1(new_n258), .B2(new_n355), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n345), .A2(new_n346), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n361), .B2(new_n208), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n273), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G58), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n243), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G58), .A2(G68), .ZN(new_n368));
  OAI21_X1  g0168(.A(G20), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n247), .A2(G159), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n360), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n272), .A2(new_n208), .A3(new_n273), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n243), .B1(new_n376), .B2(new_n363), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n255), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n358), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n342), .B1(new_n354), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n255), .ZN(new_n382));
  INV_X1    g0182(.A(new_n378), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n365), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n359), .B1(new_n377), .B2(new_n371), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n357), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n344), .A2(new_n351), .A3(new_n330), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n291), .A2(new_n343), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n280), .B2(new_n350), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n389), .B2(G169), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT18), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n344), .A2(new_n351), .A3(new_n330), .ZN(new_n392));
  AOI21_X1  g0192(.A(G169), .B1(new_n344), .B2(new_n351), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n380), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n344), .A2(new_n351), .A3(new_n306), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n389), .B2(G200), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n386), .A2(new_n398), .A3(KEYINPUT17), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n381), .A2(new_n391), .A3(new_n396), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n274), .A2(G232), .A3(new_n276), .ZN(new_n402));
  INV_X1    g0202(.A(G107), .ZN(new_n403));
  INV_X1    g0203(.A(G238), .ZN(new_n404));
  OAI221_X1 g0204(.A(new_n402), .B1(new_n403), .B2(new_n274), .C1(new_n315), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n280), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n285), .A2(G244), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(new_n291), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n320), .ZN(new_n410));
  INV_X1    g0210(.A(G87), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT15), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G87), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT74), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT74), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n245), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n355), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n208), .B2(new_n246), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n255), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n260), .A2(G77), .A3(new_n261), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(G77), .C2(new_n258), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n406), .A2(new_n330), .A3(new_n408), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n410), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n409), .A2(new_n306), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n406), .B2(new_n408), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n431), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n309), .A2(new_n341), .A3(new_n401), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT81), .ZN(new_n437));
  AOI21_X1  g0237(.A(G20), .B1(new_n271), .B2(G97), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G283), .ZN(new_n439));
  INV_X1    g0239(.A(G116), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n438), .A2(new_n439), .B1(G20), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n441), .A2(new_n255), .A3(KEYINPUT20), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT20), .B1(new_n441), .B2(new_n255), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n258), .A2(G116), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n251), .A2(KEYINPUT72), .B1(G1), .B2(G13), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n271), .A2(G1), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n447), .A2(new_n254), .A3(new_n258), .A4(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n446), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n437), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n441), .A2(new_n255), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(new_n255), .A3(KEYINPUT20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n451), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT81), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G264), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n461));
  OAI211_X1 g0261(.A(G257), .B(new_n276), .C1(new_n345), .C2(new_n346), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n272), .A2(G303), .A3(new_n273), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT80), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n461), .A2(new_n462), .A3(new_n466), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n280), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n280), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G270), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n472), .A2(new_n471), .ZN(new_n475));
  INV_X1    g0275(.A(G274), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n280), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n320), .B1(new_n469), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n460), .A2(new_n481), .A3(KEYINPUT21), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT21), .B1(new_n460), .B2(new_n481), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n283), .B1(new_n465), .B2(new_n467), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n474), .A2(G179), .A3(new_n478), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n460), .A2(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n483), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G200), .B1(new_n485), .B2(new_n479), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n452), .A3(new_n459), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(new_n493), .A3(new_n452), .A4(new_n459), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n469), .A2(G190), .A3(new_n480), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  AND2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT6), .A2(G97), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT76), .B1(new_n501), .B2(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT76), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(new_n403), .A3(KEYINPUT6), .A4(G97), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(G20), .B1(G77), .B2(new_n247), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT77), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n403), .B1(new_n376), .B2(new_n363), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G107), .B1(new_n362), .B2(new_n364), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(KEYINPUT77), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n255), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n258), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(new_n450), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(KEYINPUT4), .A2(G244), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n276), .B(new_n517), .C1(new_n345), .C2(new_n346), .ZN(new_n518));
  INV_X1    g0318(.A(G244), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n272), .B2(new_n273), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n518), .B(new_n439), .C1(new_n520), .C2(KEYINPUT4), .ZN(new_n521));
  OAI21_X1  g0321(.A(G250), .B1(new_n345), .B2(new_n346), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n276), .B1(new_n522), .B2(KEYINPUT4), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n280), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n473), .A2(G257), .B1(new_n475), .B2(new_n477), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n524), .A2(new_n330), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(G169), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n530));
  OAI211_X1 g0330(.A(G238), .B(new_n276), .C1(new_n345), .C2(new_n346), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n280), .ZN(new_n534));
  INV_X1    g0334(.A(G250), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n470), .B2(G1), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n257), .A2(new_n476), .A3(G45), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n283), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(G190), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n533), .B2(new_n280), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n432), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n544), .A2(KEYINPUT78), .A3(new_n208), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT78), .B1(new_n544), .B2(new_n208), .ZN(new_n546));
  NOR3_X1   g0346(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n208), .B(G68), .C1(new_n345), .C2(new_n346), .ZN(new_n549));
  INV_X1    g0349(.A(G97), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n245), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n549), .B1(KEYINPUT19), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n255), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n514), .A2(G87), .ZN(new_n554));
  INV_X1    g0354(.A(new_n258), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n419), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n534), .A2(G179), .A3(new_n539), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n320), .B2(new_n541), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT79), .ZN(new_n561));
  INV_X1    g0361(.A(new_n418), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n417), .B1(new_n412), .B2(new_n414), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n418), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n514), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n553), .A3(new_n556), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n543), .A2(new_n558), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n524), .A2(new_n525), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(G190), .ZN(new_n570));
  AOI21_X1  g0370(.A(G200), .B1(new_n524), .B2(new_n525), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n512), .B(new_n515), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n529), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n208), .B(G87), .C1(new_n345), .C2(new_n346), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT83), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n274), .A2(new_n577), .A3(new_n208), .A4(G87), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(KEYINPUT83), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n532), .A2(G20), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n208), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n403), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n574), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT22), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .A3(new_n581), .A4(new_n586), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n255), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n555), .A2(new_n403), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n592), .B2(new_n593), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n594), .A2(new_n596), .B1(new_n514), .B2(G107), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n598));
  OAI211_X1 g0398(.A(G250), .B(new_n276), .C1(new_n345), .C2(new_n346), .ZN(new_n599));
  INV_X1    g0399(.A(G294), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n271), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n280), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n473), .A2(G264), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n478), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G169), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n601), .A2(new_n280), .B1(new_n473), .B2(G264), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G179), .A3(new_n478), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n591), .A2(new_n597), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n591), .A2(new_n597), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n432), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n306), .A3(new_n478), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n489), .A2(new_n496), .A3(new_n573), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n436), .A2(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n436), .ZN(new_n617));
  INV_X1    g0417(.A(new_n567), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n541), .A2(new_n320), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n330), .B(new_n538), .C1(new_n533), .C2(new_n280), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT85), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n559), .B(new_n622), .C1(new_n320), .C2(new_n541), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n527), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n524), .A2(new_n330), .A3(new_n525), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n515), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n510), .A2(KEYINPUT77), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n508), .A2(new_n507), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n506), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n632), .B2(new_n255), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT86), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n557), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT86), .A4(new_n556), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n542), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n625), .A2(new_n634), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n560), .A2(new_n567), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n557), .B2(new_n542), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT26), .B1(new_n529), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n641), .A2(new_n625), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n460), .A2(new_n481), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n460), .A2(new_n487), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n605), .A2(new_n607), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n609), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(new_n482), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n624), .A2(new_n638), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n613), .A2(new_n591), .A3(new_n597), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n529), .A2(new_n572), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n645), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n617), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT87), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n338), .A2(new_n340), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n381), .A2(new_n399), .ZN(new_n663));
  INV_X1    g0463(.A(new_n304), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n307), .B(new_n663), .C1(new_n664), .C2(new_n430), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n391), .A2(new_n396), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n660), .B1(new_n668), .B2(new_n333), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n307), .A2(new_n663), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n304), .B2(new_n429), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n666), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT88), .B(new_n332), .C1(new_n672), .C2(new_n662), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n659), .A2(new_n674), .ZN(G369));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n257), .A2(new_n208), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n460), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n489), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n489), .A2(new_n496), .A3(new_n683), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n676), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT90), .ZN(new_n687));
  INV_X1    g0487(.A(new_n682), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n651), .B(new_n654), .C1(new_n610), .C2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT89), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n651), .B2(new_n688), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n608), .A2(KEYINPUT89), .A3(new_n682), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n686), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n687), .B1(new_n686), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n489), .A2(new_n682), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n698), .A2(new_n693), .B1(new_n608), .B2(new_n688), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(G399));
  AND2_X1   g0500(.A1(new_n547), .A2(new_n440), .ZN(new_n701));
  INV_X1    g0501(.A(G41), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n204), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n210), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n656), .A2(KEYINPUT93), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT93), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n652), .A2(new_n655), .A3(new_n709), .A4(new_n653), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n634), .A2(new_n640), .A3(new_n568), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n625), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n640), .B1(new_n653), .B2(new_n634), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n708), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n707), .B1(new_n715), .B2(new_n688), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n657), .A2(new_n688), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n573), .A2(new_n614), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n646), .A2(new_n647), .B1(new_n460), .B2(new_n487), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n496), .A2(new_n721), .A3(new_n482), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT31), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n541), .A2(G179), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n485), .B2(new_n479), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n569), .A2(new_n604), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n606), .A2(new_n524), .A3(new_n525), .A4(new_n541), .ZN(new_n729));
  INV_X1    g0529(.A(new_n486), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT91), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n469), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT91), .B1(new_n485), .B2(new_n486), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n728), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT92), .ZN(new_n736));
  INV_X1    g0536(.A(new_n729), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n731), .B1(new_n469), .B2(new_n730), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT91), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n734), .A2(KEYINPUT92), .A3(KEYINPUT30), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n724), .B(new_n735), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n682), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n723), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n741), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n735), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n719), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n706), .B1(new_n753), .B2(G1), .ZN(G364));
  NAND2_X1  g0554(.A1(new_n208), .A2(G13), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G45), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G1), .ZN(new_n758));
  INV_X1    g0558(.A(new_n703), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n274), .A2(new_n204), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n204), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n238), .A2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n361), .A2(new_n204), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n470), .B2(new_n211), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n207), .B1(G20), .B2(new_n320), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n760), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n330), .A2(new_n432), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n208), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n550), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n306), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n243), .B1(new_n785), .B2(new_n249), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n208), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n330), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n432), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G77), .A2(new_n790), .B1(new_n793), .B2(G107), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n208), .A2(new_n306), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n791), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n274), .C1(new_n411), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n788), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n786), .B(new_n797), .C1(G58), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n776), .A2(new_n787), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n806), .A2(KEYINPUT32), .A3(G159), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT32), .B1(new_n806), .B2(G159), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n780), .B(new_n801), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(G329), .ZN(new_n810));
  INV_X1    g0610(.A(new_n778), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G294), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n796), .B(KEYINPUT98), .Z(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT33), .B(G317), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n783), .B1(KEYINPUT99), .B2(new_n815), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n813), .A2(G303), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n361), .B1(new_n792), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G322), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n798), .A2(new_n821), .B1(new_n789), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(G326), .C2(new_n784), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n810), .A2(new_n812), .A3(new_n818), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n809), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n774), .B1(new_n771), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n684), .A2(new_n685), .ZN(new_n828));
  INV_X1    g0628(.A(new_n770), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n686), .ZN(new_n831));
  INV_X1    g0631(.A(new_n760), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n828), .A2(G330), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT100), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  AND2_X1   g0637(.A1(new_n427), .A2(new_n682), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n429), .B1(new_n434), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n430), .A2(new_n688), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n717), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n841), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n657), .A2(new_n688), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n760), .B1(new_n845), .B2(new_n751), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n751), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n771), .A2(new_n768), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n760), .B1(G77), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n806), .A2(G311), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n813), .A2(G107), .ZN(new_n852));
  INV_X1    g0652(.A(G303), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n783), .A2(new_n819), .B1(new_n785), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n361), .B1(new_n798), .B2(new_n600), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n789), .A2(new_n440), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n792), .A2(new_n411), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n851), .A2(new_n780), .A3(new_n852), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n790), .A2(G159), .B1(G137), .B2(new_n784), .ZN(new_n860));
  INV_X1    g0660(.A(G143), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n324), .B2(new_n783), .C1(new_n799), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT34), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n806), .A2(G132), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n811), .A2(G58), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n792), .A2(new_n243), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n361), .B(new_n867), .C1(new_n813), .C2(G50), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n862), .A2(new_n863), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n859), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n850), .B1(new_n871), .B2(new_n771), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n843), .B2(new_n769), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n847), .A2(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n209), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OAI211_X1 g0678(.A(new_n211), .B(G77), .C1(new_n366), .C2(new_n243), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n249), .A2(G68), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n257), .B(G13), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n394), .A2(new_n380), .ZN(new_n885));
  INV_X1    g0685(.A(new_n680), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n380), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n386), .A2(new_n398), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n885), .A2(new_n887), .A3(new_n888), .A4(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n887), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n400), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n884), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n897), .A4(new_n896), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(KEYINPUT102), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n897), .A3(new_n896), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT102), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n884), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n883), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n664), .A2(new_n688), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n890), .A2(KEYINPUT103), .A3(new_n893), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n896), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT103), .B1(new_n890), .B2(new_n893), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n884), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT39), .B1(new_n911), .B2(new_n901), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n267), .A2(new_n688), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n304), .A2(new_n307), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n304), .B2(new_n307), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n682), .B(new_n841), .C1(new_n645), .C2(new_n656), .ZN(new_n920));
  INV_X1    g0720(.A(new_n840), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n902), .A2(new_n905), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n922), .A2(new_n923), .B1(new_n667), .B2(new_n886), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n913), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n617), .B1(new_n716), .B2(new_n718), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n674), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n308), .A2(new_n914), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n304), .A2(new_n307), .A3(new_n915), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n841), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n615), .A2(KEYINPUT31), .B1(new_n744), .B2(new_n682), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n740), .A2(new_n741), .B1(new_n726), .B2(new_n727), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n747), .A2(KEYINPUT92), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n740), .A2(new_n736), .A3(new_n741), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n682), .A2(KEYINPUT31), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n932), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n929), .B1(new_n923), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n843), .B1(new_n916), .B2(new_n917), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n937), .A2(new_n938), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n746), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n929), .B1(new_n911), .B2(new_n901), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n436), .B1(new_n746), .B2(new_n943), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(G330), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n947), .B2(new_n949), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n928), .A2(new_n951), .B1(new_n257), .B2(new_n756), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n928), .A2(new_n951), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n882), .B1(new_n952), .B2(new_n953), .ZN(G367));
  NOR2_X1   g0754(.A1(new_n232), .A2(new_n765), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n772), .B1(new_n419), .B2(new_n204), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n760), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n813), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n361), .B1(new_n792), .B2(new_n550), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G283), .B2(new_n790), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n853), .C2(new_n799), .ZN(new_n961));
  INV_X1    g0761(.A(new_n796), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT46), .B1(new_n962), .B2(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT109), .B(G311), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n963), .B1(new_n784), .B2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(new_n600), .B2(new_n783), .C1(new_n778), .C2(new_n403), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n961), .B(new_n966), .C1(G317), .C2(new_n806), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n274), .B1(new_n798), .B2(new_n324), .C1(new_n861), .C2(new_n785), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G159), .B2(new_n782), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n796), .A2(new_n366), .B1(new_n789), .B2(new_n249), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n792), .A2(new_n246), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n969), .B(new_n972), .C1(new_n243), .C2(new_n778), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G137), .B2(new_n806), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  AOI21_X1  g0776(.A(new_n957), .B1(new_n976), .B2(new_n771), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n636), .A2(new_n637), .A3(new_n682), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n624), .ZN(new_n979));
  INV_X1    g0779(.A(new_n653), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n977), .B1(new_n829), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n758), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n529), .B(new_n572), .C1(new_n633), .C2(new_n688), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n529), .B2(new_n688), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n699), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT105), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n699), .A2(new_n986), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT106), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n995), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n697), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n989), .A2(new_n696), .A3(new_n996), .A4(new_n997), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n698), .A2(new_n693), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT107), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT107), .B1(new_n698), .B2(new_n693), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n752), .B1(new_n1001), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n703), .B(KEYINPUT41), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n984), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n696), .A2(new_n986), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n529), .B1(new_n985), .B2(new_n651), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT104), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n682), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n698), .A2(new_n693), .A3(new_n986), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1021), .A2(new_n1022), .B1(new_n1023), .B2(KEYINPUT42), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(KEYINPUT42), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n981), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT43), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1024), .A2(new_n1025), .A3(new_n1028), .A4(new_n1027), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1018), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1018), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n983), .B1(new_n1016), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(G387));
  OR2_X1    g0837(.A1(new_n693), .A2(new_n829), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n761), .A2(new_n701), .B1(G107), .B2(new_n204), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n228), .A2(new_n470), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n701), .B(new_n470), .C1(new_n243), .C2(new_n246), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1042));
  NOR3_X1   g0842(.A1(new_n1042), .A2(G50), .A3(new_n323), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(G50), .B2(new_n323), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n765), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n760), .B1(new_n1047), .B2(new_n773), .ZN(new_n1048));
  INV_X1    g0848(.A(G159), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n274), .B1(new_n792), .B2(new_n550), .C1(new_n785), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n962), .A2(G77), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n249), .B2(new_n798), .C1(new_n243), .C2(new_n789), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(new_n355), .C2(new_n782), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n564), .A2(new_n565), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n811), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(new_n324), .C2(new_n805), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n778), .A2(new_n819), .B1(new_n600), .B2(new_n796), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n790), .A2(G303), .B1(G322), .B2(new_n784), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n964), .A2(new_n782), .ZN(new_n1060));
  INV_X1    g0860(.A(G317), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1059), .B(new_n1060), .C1(new_n799), .C2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1057), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1058), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(KEYINPUT49), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n806), .A2(G326), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n274), .B1(new_n793), .B2(G116), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT49), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1048), .B1(new_n1070), .B2(new_n771), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1013), .A2(new_n758), .B1(new_n1038), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1012), .A2(new_n752), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n753), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n759), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1072), .A2(new_n1075), .ZN(G393));
  AOI21_X1  g0876(.A(new_n1001), .B1(new_n753), .B2(new_n1013), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1000), .B2(new_n999), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n703), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n798), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1080), .A2(G311), .B1(G317), .B2(new_n784), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n274), .B1(new_n793), .B2(G107), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n819), .B2(new_n796), .C1(new_n600), .C2(new_n789), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(G303), .C2(new_n782), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n811), .A2(G116), .B1(KEYINPUT52), .B2(new_n1081), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n821), .C2(new_n805), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n361), .B(new_n857), .C1(G68), .C2(new_n962), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n805), .B2(new_n861), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT112), .Z(new_n1090));
  NAND2_X1  g0890(.A1(new_n811), .A2(G77), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n790), .A2(new_n355), .B1(G50), .B2(new_n782), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n785), .A2(new_n324), .B1(new_n798), .B2(new_n1049), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1091), .B(new_n1092), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1087), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT113), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n771), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n986), .A2(new_n829), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT111), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n241), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n772), .B1(new_n550), .B2(new_n204), .C1(new_n1102), .C2(new_n765), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n760), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1001), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n984), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1079), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(G390));
  NOR2_X1   g0908(.A1(new_n933), .A2(new_n939), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1109), .A2(KEYINPUT114), .A3(new_n676), .A4(new_n436), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n948), .B2(G330), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n674), .B(new_n926), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n841), .A2(new_n676), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n919), .B(new_n1115), .C1(new_n933), .C2(new_n939), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n746), .B2(new_n749), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n919), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n844), .A2(new_n840), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n529), .A2(new_n624), .A3(new_n638), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n625), .B(new_n711), .C1(new_n1122), .C2(new_n640), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(KEYINPUT93), .B2(new_n656), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n682), .B1(new_n1124), .B2(new_n710), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n921), .B1(new_n1125), .B2(new_n839), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n918), .B1(new_n1109), .B2(new_n1117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1118), .A2(new_n919), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1114), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1116), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n901), .A2(KEYINPUT102), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1134), .A2(KEYINPUT101), .B1(new_n400), .B2(new_n895), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT38), .B1(new_n1135), .B2(new_n900), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n905), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT39), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n912), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1139), .A2(new_n1140), .B1(new_n922), .B2(new_n907), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n907), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n911), .B2(new_n901), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n715), .A2(new_n688), .A3(new_n839), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n840), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1144), .B1(new_n1146), .B2(new_n919), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1132), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1126), .B2(new_n918), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n918), .B1(new_n844), .B2(new_n840), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n906), .A2(new_n912), .B1(new_n1150), .B2(new_n1142), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1151), .A3(new_n1128), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1131), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1114), .A2(new_n1148), .A3(new_n1152), .A4(new_n1130), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n759), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1128), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1141), .A2(new_n1147), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1116), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n758), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n768), .B1(new_n906), .B2(new_n912), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n760), .B1(new_n355), .B2(new_n849), .ZN(new_n1163));
  INV_X1    g0963(.A(G137), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n783), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n962), .A2(G150), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT53), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G128), .C2(new_n784), .ZN(new_n1168));
  INV_X1    g0968(.A(G132), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n798), .A2(new_n1169), .B1(new_n792), .B2(new_n249), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n274), .B1(new_n789), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1168), .B(new_n1173), .C1(new_n1049), .C2(new_n778), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n806), .A2(G125), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n790), .A2(G97), .B1(G107), .B2(new_n782), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n819), .B2(new_n785), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT115), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n813), .A2(G87), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n274), .B(new_n867), .C1(G116), .C2(new_n1080), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1091), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n805), .A2(new_n600), .B1(KEYINPUT115), .B2(new_n1177), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1174), .A2(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1163), .B1(new_n1183), .B2(new_n771), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1162), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1156), .A2(new_n1161), .A3(new_n1185), .ZN(G378));
  AOI21_X1  g0986(.A(new_n676), .B1(new_n944), .B2(new_n945), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n329), .A2(new_n886), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT55), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n341), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n341), .A2(new_n1191), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1194), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n941), .A2(new_n1187), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n941), .B2(new_n1187), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n925), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n941), .A2(new_n1187), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1198), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1205), .A2(new_n1150), .B1(new_n666), .B2(new_n680), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1139), .A2(new_n1142), .A3(new_n1140), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n941), .A2(new_n1187), .A3(new_n1199), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1204), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1202), .A2(new_n1210), .A3(KEYINPUT120), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT120), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1204), .A2(new_n1208), .A3(new_n1212), .A4(new_n1209), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n758), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1199), .A2(new_n768), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n760), .B1(G50), .B2(new_n849), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n274), .A2(G41), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1051), .A2(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n366), .B2(new_n792), .C1(new_n805), .C2(new_n819), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT116), .Z(new_n1220));
  NOR2_X1   g1020(.A1(new_n798), .A2(new_n403), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT117), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n782), .A2(G97), .B1(new_n784), .B2(G116), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n778), .C2(new_n243), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1054), .B2(new_n790), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1220), .A2(KEYINPUT58), .A3(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G33), .A2(G41), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1217), .A2(G50), .A3(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT118), .B(G124), .Z(new_n1229));
  OAI221_X1 g1029(.A(new_n1227), .B1(new_n1049), .B2(new_n792), .C1(new_n805), .C2(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n796), .A2(new_n1171), .B1(new_n789), .B2(new_n1164), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G128), .B2(new_n1080), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n782), .A2(G132), .B1(new_n784), .B2(G125), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n778), .C2(new_n324), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1230), .B1(new_n1234), .B2(KEYINPUT59), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1228), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1226), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT58), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1216), .B1(new_n1240), .B2(new_n771), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1215), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1214), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1113), .B1(new_n1160), .B2(new_n1130), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1155), .A2(new_n1114), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1244), .B1(new_n1202), .B2(new_n1210), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n703), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1243), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(KEYINPUT121), .B(new_n1243), .C1(new_n1247), .C2(new_n1250), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n918), .A2(new_n768), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n760), .B1(G68), .B2(new_n849), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n806), .A2(G128), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n811), .A2(G50), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n274), .B1(new_n792), .B2(new_n366), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1169), .A2(new_n785), .B1(new_n783), .B2(new_n1171), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(G150), .C2(new_n790), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G137), .A2(new_n800), .B1(new_n813), .B2(G159), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1258), .A2(new_n1259), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n806), .A2(G303), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n813), .A2(G97), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n783), .A2(new_n440), .B1(new_n785), .B2(new_n600), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n798), .A2(new_n819), .B1(new_n789), .B2(new_n403), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n274), .A4(new_n971), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1055), .A3(new_n1266), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1257), .B1(new_n1271), .B2(new_n771), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT122), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1130), .A2(new_n758), .B1(new_n1256), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1015), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1131), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1114), .A2(new_n1130), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(G381));
  NAND3_X1  g1078(.A1(new_n1072), .A2(new_n1075), .A3(new_n836), .ZN(new_n1279));
  OR4_X1    g1079(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1279), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G387), .A2(new_n1280), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1081(.A(G378), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(G343), .C2(new_n1283), .ZN(G409));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n681), .A2(G213), .ZN(new_n1286));
  INV_X1    g1086(.A(G2897), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1130), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1113), .A2(new_n1290), .A3(new_n1121), .A4(new_n1129), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n703), .B1(new_n1114), .B2(new_n1130), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1294), .B2(new_n1274), .ZN(new_n1295));
  INV_X1    g1095(.A(G384), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1274), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1296), .B(new_n1297), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1288), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT124), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1286), .B1(new_n1302), .B2(new_n1287), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1302), .B2(new_n1287), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1299), .A2(new_n1300), .B1(new_n1301), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1301), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(KEYINPUT125), .A3(new_n1288), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1248), .A2(new_n1275), .A3(new_n1213), .A4(new_n1211), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n984), .B1(new_n1202), .B2(new_n1210), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1215), .B2(new_n1241), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G378), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(G378), .B2(new_n1251), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1286), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1305), .B(new_n1307), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G393), .A2(G396), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1315), .A2(new_n1279), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G387), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1279), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1036), .B2(KEYINPUT126), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1107), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1317), .A2(G390), .A3(new_n1319), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1251), .A2(G378), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1310), .A2(new_n1308), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1282), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1313), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1328));
  AND4_X1   g1128(.A1(new_n1285), .A2(new_n1314), .A3(new_n1323), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1301), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT123), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT123), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1327), .A2(new_n1332), .A3(new_n1301), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1329), .B1(KEYINPUT63), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1323), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT62), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(new_n1285), .A3(new_n1314), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1336), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1243), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT121), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1346));
  AOI21_X1  g1146(.A(G378), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1251), .A2(new_n1282), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1301), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1348), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1283), .A2(new_n1306), .A3(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1349), .A2(new_n1323), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1323), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1352), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  AOI211_X1 g1155(.A(KEYINPUT127), .B(new_n1323), .C1(new_n1349), .C2(new_n1351), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(G402));
endmodule


