//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  OR2_X1    g000(.A1(KEYINPUT2), .A2(G113), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT2), .A2(G113), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n187), .A2(new_n194), .A3(new_n196), .A4(new_n188), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT71), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n189), .A2(new_n191), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI22_X1  g020(.A1(KEYINPUT65), .A2(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(G131), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G134), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n206), .A2(KEYINPUT67), .A3(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT65), .B(new_n205), .C1(new_n206), .C2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n208), .A2(new_n210), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT69), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n212), .B2(G134), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n206), .B2(G137), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n218), .A2(new_n212), .A3(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(KEYINPUT1), .A3(G146), .ZN(new_n231));
  XNOR2_X1  g045(.A(G143), .B(G146), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(new_n231), .C1(G128), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT72), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n229), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n224), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n231), .A4(new_n230), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n202), .A2(KEYINPUT11), .B1(new_n212), .B2(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n216), .B1(new_n240), .B2(new_n203), .ZN(new_n241));
  INV_X1    g055(.A(new_n215), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n217), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n227), .B2(new_n229), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT64), .B1(new_n232), .B2(new_n247), .ZN(new_n250));
  AND4_X1   g064(.A1(KEYINPUT64), .A2(new_n227), .A3(new_n229), .A4(new_n247), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n223), .A2(new_n239), .B1(new_n244), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n244), .A2(new_n253), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n244), .A2(new_n258), .A3(new_n253), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n217), .A2(new_n222), .A3(new_n233), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n217), .A2(new_n222), .A3(new_n233), .A4(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n257), .A2(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n201), .B(new_n255), .C1(new_n264), .C2(KEYINPUT30), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT73), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n239), .A2(new_n223), .ZN(new_n267));
  INV_X1    g081(.A(new_n201), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n256), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT74), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n254), .A2(new_n271), .A3(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n263), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n244), .A2(new_n258), .A3(new_n253), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n258), .B1(new_n244), .B2(new_n253), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n201), .A4(new_n255), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n266), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G237), .A2(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G210), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n284), .B(KEYINPUT27), .Z(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT26), .ZN(new_n286));
  INV_X1    g100(.A(G101), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n277), .A2(new_n201), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n273), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n269), .A2(new_n292), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OR3_X1    g110(.A1(new_n294), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n254), .A2(new_n268), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n270), .B2(new_n272), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT29), .B(new_n295), .C1(new_n301), .C2(new_n292), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n302), .B2(new_n289), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n254), .A2(new_n268), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n271), .B1(new_n254), .B2(new_n268), .ZN(new_n305));
  AND4_X1   g119(.A1(new_n271), .A2(new_n267), .A3(new_n256), .A4(new_n268), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n307), .B2(KEYINPUT28), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT75), .A3(KEYINPUT29), .A4(new_n288), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n266), .A2(new_n288), .A3(new_n273), .A4(new_n281), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n315), .A2(KEYINPUT31), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n289), .B1(new_n294), .B2(new_n296), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n315), .B2(KEYINPUT31), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT32), .B(new_n314), .C1(new_n316), .C2(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n325), .A2(G952), .ZN(new_n326));
  NAND2_X1  g140(.A1(G234), .A2(G237), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT21), .B(G898), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(G902), .A3(G953), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT6), .ZN(new_n337));
  INV_X1    g151(.A(G104), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT3), .B1(new_n338), .B2(G107), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n340));
  INV_X1    g154(.A(G107), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(G107), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n344), .A2(new_n345), .A3(G101), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n199), .B2(new_n200), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(G101), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n339), .A2(new_n342), .A3(new_n287), .A4(new_n343), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  OAI211_X1 g166(.A(KEYINPUT4), .B(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT85), .B1(new_n341), .B2(G104), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n341), .A2(G104), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n341), .A2(KEYINPUT85), .A3(G104), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n287), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n339), .A2(new_n342), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n287), .A4(new_n343), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n349), .A2(new_n350), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n192), .A2(new_n198), .B1(new_n364), .B2(G113), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n347), .A2(new_n353), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(G110), .B(G122), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n337), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n347), .A2(new_n353), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(new_n365), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n367), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT91), .B(G224), .Z(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G953), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n233), .A2(G125), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n252), .A2(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n378), .A2(new_n379), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n383), .ZN(new_n385));
  INV_X1    g199(.A(new_n377), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n381), .A3(new_n380), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n372), .A2(new_n367), .A3(new_n337), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n374), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT92), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n374), .A2(new_n392), .A3(new_n388), .A4(new_n389), .ZN(new_n393));
  AOI21_X1  g207(.A(G902), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G210), .B1(G237), .B2(G902), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n382), .A2(new_n383), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n386), .A2(KEYINPUT7), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n362), .B(new_n365), .Z(new_n399));
  XNOR2_X1  g213(.A(new_n367), .B(KEYINPUT8), .ZN(new_n400));
  OAI221_X1 g214(.A(new_n398), .B1(new_n367), .B2(new_n372), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n395), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n395), .B1(new_n394), .B2(new_n401), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n324), .B(new_n335), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G116), .B(G122), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n341), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n195), .A2(G122), .ZN(new_n408));
  INV_X1    g222(.A(G122), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(G116), .ZN(new_n410));
  OAI21_X1  g224(.A(G107), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n226), .A2(G128), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n224), .A2(G143), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n206), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT13), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n224), .B2(G143), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n226), .A2(KEYINPUT13), .A3(G128), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G134), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n406), .B1(KEYINPUT14), .B2(new_n341), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n195), .B2(G122), .ZN(new_n423));
  OAI211_X1 g237(.A(G107), .B(new_n423), .C1(new_n408), .C2(new_n410), .ZN(new_n424));
  INV_X1    g238(.A(new_n415), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n206), .B1(new_n413), .B2(new_n414), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n422), .B(new_n424), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT9), .B(G234), .Z(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G217), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n429), .A2(new_n430), .A3(G953), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n421), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n421), .B2(new_n427), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n421), .A2(new_n427), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n437), .A2(new_n433), .A3(new_n431), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n436), .A2(new_n438), .A3(G902), .ZN(new_n439));
  INV_X1    g253(.A(G478), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT15), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n441), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT99), .ZN(new_n446));
  OR2_X1    g260(.A1(KEYINPUT93), .A2(G143), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(G214), .B2(new_n283), .ZN(new_n448));
  INV_X1    g262(.A(G237), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n325), .A3(G214), .ZN(new_n450));
  NOR2_X1   g264(.A1(KEYINPUT93), .A2(G143), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n209), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n451), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(G214), .A3(new_n283), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n210), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n453), .A2(new_n454), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n453), .A2(KEYINPUT95), .A3(new_n454), .A4(new_n457), .ZN(new_n462));
  INV_X1    g276(.A(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G125), .ZN(new_n464));
  INV_X1    g278(.A(G125), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G140), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT16), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n465), .A2(KEYINPUT16), .A3(G140), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n467), .A2(G146), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G146), .B1(new_n467), .B2(new_n468), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G113), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n338), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT18), .A2(G131), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n456), .A2(new_n455), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n456), .B2(new_n455), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT79), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n464), .A2(new_n466), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n464), .B2(new_n466), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n228), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n464), .A2(new_n466), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G146), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n472), .A2(new_n474), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n469), .B1(new_n453), .B2(new_n457), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT19), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n480), .B2(new_n481), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n483), .A2(KEYINPUT19), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n228), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  INV_X1    g308(.A(new_n474), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(KEYINPUT94), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n488), .A2(new_n492), .B1(new_n478), .B2(new_n485), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n474), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n502), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n487), .A2(new_n496), .A3(new_n499), .A4(KEYINPUT96), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n503), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  INV_X1    g323(.A(new_n487), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n474), .B1(new_n472), .B2(new_n486), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n311), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT97), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(new_n311), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(G475), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n444), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n446), .A2(new_n509), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n405), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n469), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n193), .B2(G128), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n193), .A2(G128), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G110), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT24), .B(G110), .Z(new_n528));
  NAND2_X1  g342(.A1(new_n224), .A2(G119), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n524), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT77), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n524), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n528), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n521), .B(new_n482), .C1(new_n527), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT22), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(G137), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT78), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n526), .A2(new_n539), .A3(G110), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n526), .B2(G110), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n540), .A2(new_n541), .B1(new_n469), .B2(new_n470), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n531), .A2(new_n533), .A3(new_n528), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n535), .B(new_n538), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT80), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n535), .B(new_n548), .C1(new_n543), .C2(new_n542), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n538), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT81), .B1(new_n552), .B2(new_n311), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT82), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT25), .ZN(new_n555));
  INV_X1    g369(.A(G234), .ZN(new_n556));
  OAI21_X1  g370(.A(G217), .B1(new_n556), .B2(G902), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT76), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n552), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n554), .B1(new_n561), .B2(G902), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(KEYINPUT25), .C1(new_n553), .C2(new_n554), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n558), .A2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n552), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n362), .A2(new_n233), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n362), .A2(new_n233), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n244), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT12), .B(new_n244), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n234), .B2(new_n238), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n362), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT87), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n582), .A3(new_n362), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n252), .A2(new_n346), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n353), .A2(new_n585), .A3(KEYINPUT84), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT84), .B1(new_n353), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n244), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT86), .B(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n570), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n584), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G140), .ZN(new_n593));
  INV_X1    g407(.A(G227), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G953), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n593), .B(new_n595), .Z(new_n596));
  AND3_X1   g410(.A1(new_n577), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n579), .A2(new_n582), .A3(new_n362), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n582), .B1(new_n579), .B2(new_n362), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n591), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n587), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n353), .A2(new_n585), .A3(KEYINPUT84), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n244), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n596), .B1(new_n604), .B2(new_n592), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n569), .B(new_n311), .C1(new_n597), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n569), .A2(new_n311), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n577), .A2(new_n592), .ZN(new_n609));
  INV_X1    g423(.A(new_n596), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n604), .A2(new_n592), .A3(new_n596), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(G469), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n606), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(G221), .B1(new_n429), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(KEYINPUT88), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n323), .A2(new_n520), .A3(new_n568), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  AND4_X1   g436(.A1(new_n280), .A2(new_n279), .A3(new_n201), .A4(new_n255), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n267), .A2(new_n256), .A3(KEYINPUT30), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n277), .B2(new_n278), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n280), .B1(new_n625), .B2(new_n201), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT31), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n288), .A4(new_n273), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n315), .A2(KEYINPUT31), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n317), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n311), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(G472), .B1(new_n314), .B2(new_n631), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n620), .A2(new_n633), .A3(new_n568), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n436), .B2(new_n438), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n432), .B1(new_n435), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n437), .A2(KEYINPUT101), .A3(new_n431), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT33), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n440), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n439), .A2(G478), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT102), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n439), .A2(G478), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n646), .B(new_n647), .C1(new_n440), .C2(new_n642), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n509), .A2(new_n516), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n391), .A2(new_n393), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n311), .A3(new_n401), .ZN(new_n653));
  INV_X1    g467(.A(new_n395), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n402), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n404), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n324), .A3(new_n335), .A4(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n634), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(new_n516), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n506), .A2(new_n507), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n502), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT20), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n508), .A2(new_n501), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n501), .B1(new_n664), .B2(new_n502), .ZN(new_n670));
  AOI211_X1 g484(.A(KEYINPUT20), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT103), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n663), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n446), .A2(new_n518), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n659), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n634), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT35), .B(G107), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NOR2_X1   g493(.A1(new_n551), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n550), .B(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n560), .A2(new_n563), .B1(new_n565), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n682), .A2(new_n519), .A3(new_n334), .ZN(new_n683));
  INV_X1    g497(.A(new_n324), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n655), .B2(new_n402), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n620), .A3(new_n633), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT37), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(G110), .Z(G12));
  AND3_X1   g503(.A1(new_n614), .A2(KEYINPUT88), .A3(new_n615), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT88), .B1(new_n614), .B2(new_n615), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n322), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT32), .B1(new_n631), .B2(new_n314), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n692), .B1(new_n695), .B2(new_n313), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n656), .A2(new_n324), .A3(new_n658), .ZN(new_n697));
  INV_X1    g511(.A(new_n682), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n669), .A2(new_n672), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n332), .A2(G900), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n328), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n516), .A2(new_n699), .A3(new_n674), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT105), .B1(new_n301), .B2(new_n288), .ZN(new_n706));
  OR3_X1    g520(.A1(new_n301), .A2(KEYINPUT105), .A3(new_n288), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n315), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n321), .A2(new_n322), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n698), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT40), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n701), .B(KEYINPUT39), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n620), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n655), .A2(new_n402), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT38), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n674), .A2(new_n650), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n620), .A2(new_n714), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n324), .B(new_n720), .C1(new_n721), .C2(new_n713), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n705), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n620), .A2(new_n714), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n684), .B(new_n719), .C1(new_n724), .C2(KEYINPUT40), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n715), .A2(new_n717), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(KEYINPUT106), .A3(new_n712), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n226), .ZN(G45));
  INV_X1    g543(.A(new_n701), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n682), .A2(new_n651), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n323), .A2(new_n697), .A3(new_n620), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT107), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n228), .ZN(G48));
  NOR2_X1   g548(.A1(new_n659), .A2(new_n651), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n311), .B1(new_n597), .B2(new_n605), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n737), .A2(new_n615), .A3(new_n606), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n735), .A2(new_n323), .A3(new_n568), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND3_X1  g555(.A1(new_n323), .A2(new_n568), .A3(new_n738), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n676), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n195), .ZN(G18));
  AND4_X1   g558(.A1(new_n324), .A2(new_n738), .A3(new_n656), .A4(new_n658), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n323), .A3(new_n683), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NAND3_X1  g561(.A1(new_n656), .A2(new_n324), .A3(new_n658), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n719), .ZN(new_n749));
  INV_X1    g563(.A(G472), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n631), .B2(new_n311), .ZN(new_n751));
  INV_X1    g565(.A(new_n314), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n308), .A2(new_n288), .ZN(new_n753));
  INV_X1    g567(.A(new_n315), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n753), .B1(new_n754), .B2(new_n628), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n752), .B1(new_n755), .B2(new_n630), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n751), .A2(new_n567), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n749), .A2(new_n757), .A3(new_n335), .A4(new_n738), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NOR3_X1   g573(.A1(new_n751), .A2(new_n756), .A3(new_n682), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n651), .A2(new_n730), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n745), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  NAND2_X1  g577(.A1(new_n606), .A2(new_n608), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n612), .A2(KEYINPUT109), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n612), .A2(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n611), .A2(KEYINPUT108), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n609), .A2(new_n768), .A3(new_n610), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n764), .B1(new_n770), .B2(G469), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n655), .A2(new_n324), .A3(new_n402), .ZN(new_n772));
  INV_X1    g586(.A(new_n615), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n323), .A2(new_n774), .A3(new_n568), .A4(new_n761), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(KEYINPUT110), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n777), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  NAND4_X1  g594(.A1(new_n323), .A2(new_n774), .A3(new_n568), .A4(new_n702), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  AOI21_X1  g596(.A(new_n650), .B1(new_n645), .B2(new_n648), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT43), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n650), .B2(KEYINPUT112), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n785), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n633), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n698), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n772), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n766), .A2(new_n765), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n767), .A2(new_n769), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT45), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n611), .A2(new_n612), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n802), .A3(G469), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n800), .A2(new_n802), .A3(KEYINPUT111), .A4(G469), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n607), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n606), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n773), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n793), .A4(new_n794), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n797), .A2(new_n811), .A3(new_n714), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G137), .ZN(G39));
  OAI21_X1  g628(.A(KEYINPUT47), .B1(new_n810), .B2(new_n773), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n323), .A2(new_n568), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n615), .C1(new_n808), .C2(new_n809), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n772), .A2(new_n651), .A3(new_n730), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n815), .A2(new_n816), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND2_X1  g635(.A1(new_n793), .A2(new_n738), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n711), .A2(new_n823), .A3(new_n329), .A4(new_n568), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n328), .B1(new_n786), .B2(new_n787), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n823), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n567), .B1(new_n695), .B2(new_n313), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI221_X1 g642(.A(new_n326), .B1(new_n651), .B2(new_n824), .C1(new_n828), .C2(KEYINPUT48), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(KEYINPUT48), .B2(new_n828), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n824), .A2(new_n650), .A3(new_n649), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n825), .A2(new_n757), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n738), .A2(new_n684), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n717), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n834), .A4(new_n836), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n831), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n826), .A2(new_n760), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n737), .A2(new_n606), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n615), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n815), .B2(new_n818), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n832), .A2(new_n793), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n841), .B(new_n842), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n830), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n852));
  XNOR2_X1  g666(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n852), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n323), .A2(new_n620), .A3(new_n698), .A4(new_n702), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n762), .B(new_n732), .C1(new_n858), .C2(new_n748), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n771), .A2(new_n773), .A3(new_n730), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n749), .A2(new_n682), .A3(new_n710), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n857), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n762), .A2(new_n732), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n703), .A3(new_n861), .A4(KEYINPUT52), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n645), .A2(new_n648), .B1(new_n509), .B2(new_n516), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n509), .A2(new_n516), .A3(new_n444), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n405), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n620), .A3(new_n633), .A4(new_n568), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n621), .A2(new_n686), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n743), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n760), .A2(new_n774), .A3(new_n761), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n323), .A2(new_n620), .A3(new_n698), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n699), .A2(new_n516), .A3(new_n445), .A4(new_n701), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT114), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n673), .A2(new_n878), .A3(new_n445), .A4(new_n701), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n793), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n781), .B(new_n874), .C1(new_n875), .C2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n739), .A2(new_n758), .A3(new_n746), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n779), .A2(new_n873), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n856), .B1(new_n866), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n659), .A2(new_n675), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n827), .A2(new_n886), .A3(new_n738), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n621), .A3(new_n686), .A4(new_n871), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n739), .A2(new_n758), .A3(new_n746), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n881), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n863), .A2(new_n865), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT53), .A4(new_n779), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n885), .A2(KEYINPUT115), .A3(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n779), .A2(new_n873), .A3(new_n882), .A4(new_n883), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n849), .A2(new_n852), .A3(new_n853), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n885), .A2(new_n899), .A3(new_n892), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n855), .A2(new_n897), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n832), .A2(new_n745), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n901), .A2(new_n902), .B1(G952), .B2(G953), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n568), .A2(new_n324), .A3(new_n615), .A4(new_n783), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n843), .B(KEYINPUT49), .ZN(new_n905));
  OR4_X1    g719(.A1(new_n710), .A2(new_n904), .A3(new_n717), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(G75));
  AOI21_X1  g721(.A(new_n311), .B1(new_n885), .B2(new_n892), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(G210), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n374), .A2(new_n389), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n388), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT55), .Z(new_n914));
  AND2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n911), .A2(new_n914), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n325), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  NOR3_X1   g732(.A1(new_n866), .A2(new_n884), .A3(new_n856), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n894), .B2(new_n891), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT54), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT120), .A3(new_n900), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n885), .A2(new_n892), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT54), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n607), .B(KEYINPUT57), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n605), .B2(new_n597), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n908), .A2(new_n805), .A3(new_n806), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n917), .B1(new_n928), .B2(new_n929), .ZN(G54));
  NAND2_X1  g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n908), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n664), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n917), .ZN(G60));
  NAND2_X1  g752(.A1(new_n897), .A2(new_n900), .ZN(new_n939));
  XNOR2_X1  g753(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n440), .A2(new_n311), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n636), .A2(new_n641), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  INV_X1    g762(.A(new_n917), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n942), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n922), .A2(new_n925), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n949), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n945), .B1(new_n939), .B2(new_n943), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT123), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(G63));
  OAI21_X1  g770(.A(KEYINPUT60), .B1(new_n430), .B2(new_n311), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n430), .A2(new_n311), .A3(KEYINPUT60), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n923), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n917), .B1(new_n959), .B2(new_n561), .ZN(new_n960));
  INV_X1    g774(.A(new_n681), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G66));
  OAI21_X1  g778(.A(G953), .B1(new_n376), .B2(new_n331), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n888), .A2(new_n889), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n912), .B1(G898), .B2(new_n325), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  INV_X1    g783(.A(new_n869), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n827), .A2(new_n793), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n721), .B1(KEYINPUT124), .B2(new_n970), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n859), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n723), .A2(new_n727), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n813), .A2(new_n820), .ZN(new_n981));
  AOI21_X1  g795(.A(G953), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n490), .A2(new_n491), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n625), .B(new_n983), .Z(new_n984));
  AOI21_X1  g798(.A(new_n325), .B1(G227), .B2(G900), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n594), .A2(G900), .A3(G953), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n779), .A2(new_n781), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT125), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n813), .A3(new_n820), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n811), .A2(new_n714), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n827), .A2(new_n749), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n975), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT126), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  INV_X1    g809(.A(new_n993), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n981), .A2(new_n995), .A3(new_n996), .A4(new_n989), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n987), .B1(new_n998), .B2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n986), .B1(new_n999), .B2(new_n984), .ZN(G72));
  AND3_X1   g814(.A1(new_n980), .A2(new_n966), .A3(new_n981), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n288), .B(new_n282), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n754), .A2(KEYINPUT127), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1004), .B1(new_n1006), .B2(new_n290), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n282), .A2(KEYINPUT127), .A3(new_n289), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n893), .A2(new_n896), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1005), .A2(new_n949), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n994), .A2(new_n997), .A3(new_n966), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n282), .B1(new_n1011), .B2(new_n1003), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1010), .B1(new_n289), .B2(new_n1012), .ZN(G57));
endmodule


