//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT25), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT22), .B(G137), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(G146), .B(new_n196), .C1(new_n200), .C2(new_n194), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT73), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n207), .C1(G119), .C2(new_n206), .ZN(new_n208));
  XNOR2_X1  g022(.A(G119), .B(G128), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT24), .B(G110), .Z(new_n210));
  OAI22_X1  g024(.A1(new_n208), .A2(G110), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G125), .B(G140), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G146), .A4(new_n196), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n202), .A2(new_n211), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n208), .A2(G110), .B1(new_n209), .B2(new_n210), .ZN(new_n219));
  INV_X1    g033(.A(new_n201), .ZN(new_n220));
  AOI21_X1  g034(.A(G146), .B1(new_n215), .B2(new_n196), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n193), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n222), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT74), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n222), .A3(KEYINPUT74), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n228), .B2(new_n193), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n188), .B1(new_n229), .B2(G902), .ZN(new_n230));
  INV_X1    g044(.A(G902), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n192), .B1(new_n226), .B2(new_n227), .ZN(new_n232));
  OAI221_X1 g046(.A(new_n231), .B1(new_n187), .B2(KEYINPUT25), .C1(new_n232), .C2(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(G234), .B2(new_n231), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(G902), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n232), .B2(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT9), .B(G234), .ZN(new_n242));
  OAI21_X1  g056(.A(G221), .B1(new_n242), .B2(G902), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(G110), .B(G140), .Z(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT76), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n190), .A2(G227), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n213), .A2(G143), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n213), .A2(KEYINPUT64), .A3(G143), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n256), .A2(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n251), .B2(G146), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(KEYINPUT65), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n256), .A3(new_n259), .A4(new_n252), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n255), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G104), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n267), .A2(KEYINPUT3), .A3(G107), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OR2_X1    g083(.A1(KEYINPUT77), .A2(G104), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT77), .A2(G104), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G107), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(G107), .B1(new_n270), .B2(new_n271), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n269), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G101), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n278));
  INV_X1    g092(.A(G101), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT4), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G107), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT77), .A2(G104), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT77), .A2(G104), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n268), .B1(new_n285), .B2(KEYINPUT3), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n279), .B1(new_n286), .B2(new_n272), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n266), .B(new_n277), .C1(new_n281), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n283), .A2(new_n284), .ZN(new_n289));
  AOI21_X1  g103(.A(G101), .B1(new_n289), .B2(G107), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n267), .A2(G107), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n286), .A2(new_n290), .B1(new_n292), .B2(G101), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n250), .A2(new_n252), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  OAI21_X1  g110(.A(G128), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT67), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n261), .A2(new_n256), .A3(new_n300), .A4(new_n252), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n293), .A2(new_n302), .A3(KEYINPUT10), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n261), .A2(new_n252), .A3(new_n256), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(G128), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n301), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n304), .B(KEYINPUT10), .C1(new_n293), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n286), .A2(new_n290), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n292), .A2(G101), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT10), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT78), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n288), .B(new_n303), .C1(new_n309), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n321), .A3(new_n324), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n249), .B1(new_n315), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT80), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n329), .B(new_n249), .C1(new_n315), .C2(new_n326), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n293), .B2(new_n302), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n310), .A2(new_n311), .ZN(new_n333));
  INV_X1    g147(.A(new_n301), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n295), .A2(new_n296), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n250), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(G128), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n337), .B2(new_n294), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n338), .A3(KEYINPUT79), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(new_n339), .A3(new_n312), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n326), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(KEYINPUT12), .A3(new_n326), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n328), .A2(new_n330), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n315), .A2(new_n326), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n315), .A2(new_n326), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n248), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G469), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n231), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n340), .A2(KEYINPUT12), .A3(new_n326), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT12), .B1(new_n340), .B2(new_n326), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n354), .A2(new_n355), .B1(new_n326), .B2(new_n315), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n288), .A2(new_n303), .ZN(new_n357));
  INV_X1    g171(.A(new_n309), .ZN(new_n358));
  INV_X1    g172(.A(new_n314), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n326), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n248), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n356), .A2(new_n248), .B1(new_n362), .B2(new_n347), .ZN(new_n363));
  OAI21_X1  g177(.A(G469), .B1(new_n363), .B2(G902), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n244), .B1(new_n353), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n266), .A2(new_n326), .ZN(new_n366));
  INV_X1    g180(.A(new_n319), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n317), .A2(G137), .ZN(new_n368));
  OAI21_X1  g182(.A(G131), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n369), .A2(new_n325), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n302), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT2), .B(G113), .Z(new_n372));
  XNOR2_X1  g186(.A(G116), .B(G119), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n366), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G237), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT69), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G237), .ZN(new_n380));
  AOI21_X1  g194(.A(G953), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G210), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT27), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n384), .A3(G210), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT26), .B(G101), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n386), .B1(new_n383), .B2(new_n385), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n376), .A2(KEYINPUT70), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT70), .B1(new_n376), .B2(new_n389), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT68), .ZN(new_n393));
  INV_X1    g207(.A(new_n371), .ZN(new_n394));
  INV_X1    g208(.A(new_n255), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n263), .A2(new_n264), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n263), .A2(new_n264), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n361), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n393), .B1(new_n402), .B2(KEYINPUT30), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n326), .B1(new_n266), .B2(KEYINPUT66), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n399), .B(new_n255), .C1(new_n262), .C2(new_n265), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n371), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(KEYINPUT68), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n366), .A2(new_n371), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n375), .B1(new_n410), .B2(KEYINPUT30), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n392), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n413));
  INV_X1    g227(.A(new_n389), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n376), .A2(KEYINPUT28), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n376), .A2(KEYINPUT28), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n406), .A2(new_n374), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT71), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n406), .A2(KEYINPUT68), .A3(new_n407), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT68), .B1(new_n406), .B2(new_n407), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n411), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n392), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n421), .B1(new_n426), .B2(KEYINPUT31), .ZN(new_n427));
  AOI211_X1 g241(.A(KEYINPUT71), .B(new_n413), .C1(new_n424), .C2(new_n425), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G472), .A2(G902), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT72), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT32), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n410), .A2(new_n375), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n415), .B2(new_n416), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT29), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n414), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n389), .B1(new_n424), .B2(new_n376), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n436), .B1(new_n419), .B2(new_n414), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G472), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n424), .A2(new_n413), .A3(new_n425), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n419), .A2(new_n414), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n374), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n403), .B2(new_n408), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT31), .B1(new_n448), .B2(new_n392), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT71), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n426), .A2(new_n421), .A3(KEYINPUT31), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n431), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n442), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n241), .B(new_n365), .C1(new_n433), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n379), .A2(G237), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n460));
  OAI211_X1 g274(.A(G214), .B(new_n190), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n251), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n381), .A2(G143), .A3(G214), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n464), .B2(G131), .ZN(new_n465));
  AOI211_X1 g279(.A(KEYINPUT87), .B(new_n324), .C1(new_n462), .C2(new_n463), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT17), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n196), .B1(new_n200), .B2(new_n194), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n213), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n201), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT89), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n378), .A2(new_n380), .ZN(new_n472));
  AND4_X1   g286(.A1(G143), .A2(new_n472), .A3(G214), .A4(new_n190), .ZN(new_n473));
  AOI21_X1  g287(.A(G143), .B1(new_n381), .B2(G214), .ZN(new_n474));
  OAI21_X1  g288(.A(G131), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT87), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n464), .A2(new_n458), .A3(G131), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n462), .A2(new_n324), .A3(new_n463), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n462), .A2(KEYINPUT86), .A3(new_n463), .A4(new_n324), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n476), .A2(new_n477), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n467), .B(new_n471), .C1(new_n482), .C2(KEYINPUT17), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT18), .A2(G131), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n462), .A2(new_n484), .A3(new_n463), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n200), .A2(G146), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n214), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT84), .B1(new_n473), .B2(new_n474), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n462), .A2(new_n492), .A3(new_n463), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n484), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT85), .B(new_n484), .C1(new_n491), .C2(new_n493), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n489), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G113), .B(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n267), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n483), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n483), .B2(new_n498), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n231), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT90), .B(new_n231), .C1(new_n501), .C2(new_n502), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(G475), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n202), .A2(new_n217), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n212), .B(KEYINPUT19), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n213), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n513), .A3(new_n213), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n482), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n500), .B1(new_n498), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n508), .B1(new_n501), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT20), .ZN(new_n519));
  INV_X1    g333(.A(new_n500), .ZN(new_n520));
  INV_X1    g334(.A(new_n493), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n492), .B1(new_n462), .B2(new_n463), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n495), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n494), .A2(new_n490), .A3(new_n495), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n488), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n482), .A2(new_n515), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n483), .A2(new_n498), .A3(new_n500), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n508), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n251), .A2(G128), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n251), .A2(G128), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n317), .ZN(new_n538));
  INV_X1    g352(.A(G116), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT14), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT91), .B(G122), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n539), .ZN(new_n543));
  OAI21_X1  g357(.A(G107), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n282), .B(new_n540), .C1(new_n542), .C2(new_n539), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n540), .ZN(new_n547));
  OAI21_X1  g361(.A(G107), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n545), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n537), .A2(new_n317), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n534), .B1(new_n536), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(KEYINPUT92), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(KEYINPUT92), .B1(KEYINPUT13), .B2(new_n535), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n317), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n546), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n242), .A2(new_n235), .A3(G953), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n546), .B(new_n558), .C1(new_n551), .C2(new_n556), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n231), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n231), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G952), .ZN(new_n573));
  AOI211_X1 g387(.A(G953), .B(new_n573), .C1(G234), .C2(G237), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT21), .B(G898), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT94), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n231), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n507), .A2(new_n533), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G210), .B1(G237), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n373), .A2(KEYINPUT5), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n539), .A2(KEYINPUT5), .A3(G119), .ZN(new_n585));
  INV_X1    g399(.A(G113), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n372), .A2(new_n373), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n310), .A2(new_n588), .A3(new_n311), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n281), .A2(new_n287), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n277), .A2(new_n374), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G122), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n594), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(KEYINPUT6), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT6), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n593), .A2(new_n599), .A3(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n338), .A2(new_n198), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n266), .B2(new_n198), .ZN(new_n602));
  INV_X1    g416(.A(G224), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G953), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT81), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n602), .B(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n598), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n588), .A2(new_n589), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n333), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n590), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n594), .B(KEYINPUT8), .Z(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT82), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT82), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n614), .B(new_n611), .C1(new_n609), .C2(new_n590), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT7), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n605), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n602), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n601), .B(new_n618), .C1(new_n198), .C2(new_n266), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n597), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n231), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n583), .B1(new_n607), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n611), .B1(new_n609), .B2(new_n590), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT82), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n620), .A2(new_n597), .A3(new_n621), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n598), .A2(new_n606), .A3(new_n600), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n582), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n624), .A2(KEYINPUT83), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(G214), .B1(G237), .B2(G902), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT83), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n633), .B(new_n583), .C1(new_n607), .C2(new_n623), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n581), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n457), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(new_n279), .ZN(G3));
  OAI21_X1  g453(.A(G472), .B1(new_n452), .B2(G902), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n429), .A2(new_n432), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n365), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n240), .ZN(new_n643));
  INV_X1    g457(.A(G475), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n483), .A2(new_n498), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n520), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n646), .B2(new_n529), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n647), .B2(KEYINPUT90), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n648), .A2(new_n505), .B1(new_n519), .B2(new_n532), .ZN(new_n649));
  INV_X1    g463(.A(new_n632), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n582), .B1(new_n628), .B2(new_n629), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n624), .A2(KEYINPUT95), .A3(new_n630), .ZN(new_n654));
  INV_X1    g468(.A(new_n579), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n557), .B2(new_n559), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n554), .A2(new_n555), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n550), .B(new_n549), .C1(new_n659), .C2(new_n317), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(KEYINPUT96), .A3(new_n546), .A4(new_n558), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n561), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT97), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n658), .A2(new_n663), .A3(new_n666), .A4(new_n661), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n562), .A2(new_n657), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n564), .A2(G902), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n665), .A2(new_n667), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n563), .A2(new_n564), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n649), .A2(new_n656), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n643), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT34), .B(G104), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  AND3_X1   g491(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT98), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n531), .B1(new_n530), .B2(new_n508), .ZN(new_n680));
  INV_X1    g494(.A(new_n508), .ZN(new_n681));
  AOI211_X1 g495(.A(KEYINPUT20), .B(new_n681), .C1(new_n528), .C2(new_n529), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n679), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n519), .A2(new_n532), .A3(KEYINPUT98), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n569), .A2(new_n571), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n648), .B2(new_n505), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n678), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n643), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT35), .B(G107), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  INV_X1    g505(.A(new_n635), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n193), .A2(KEYINPUT36), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n228), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n228), .A2(new_n693), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n694), .A2(new_n238), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n234), .B2(new_n236), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n692), .A2(new_n649), .A3(new_n580), .A4(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n642), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT37), .B(G110), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT99), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G12));
  AOI211_X1 g517(.A(new_n244), .B(new_n697), .C1(new_n353), .C2(new_n364), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n433), .B2(new_n456), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n653), .A2(new_n654), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT100), .B(G900), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n574), .B1(new_n578), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n685), .A3(new_n687), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT101), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  AOI211_X1 g525(.A(G469), .B(G902), .C1(new_n346), .C2(new_n350), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n356), .A2(new_n248), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n362), .A2(new_n347), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n352), .B1(new_n715), .B2(new_n231), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n243), .B(new_n698), .C1(new_n712), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(G472), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n415), .A2(new_n416), .B1(new_n374), .B2(new_n406), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT29), .B1(new_n719), .B2(new_n389), .ZN(new_n720));
  INV_X1    g534(.A(new_n376), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n409), .B2(new_n411), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n720), .B1(new_n722), .B2(new_n389), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n718), .B1(new_n723), .B2(new_n438), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n429), .B2(new_n454), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n453), .B1(new_n452), .B2(new_n431), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n717), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n706), .A2(new_n685), .A3(new_n687), .A4(new_n709), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n711), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G128), .ZN(G30));
  OAI21_X1  g546(.A(new_n414), .B1(new_n434), .B2(new_n721), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n426), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n718), .B1(new_n734), .B2(new_n231), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n429), .B2(new_n454), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n726), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT102), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n686), .B1(new_n507), .B2(new_n533), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n632), .A3(new_n697), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT103), .Z(new_n741));
  XOR2_X1   g555(.A(new_n708), .B(KEYINPUT39), .Z(new_n742));
  NAND2_X1  g556(.A1(new_n365), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT40), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n631), .A2(new_n634), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT38), .Z(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  OR4_X1    g561(.A1(new_n738), .A2(new_n741), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  AOI21_X1  g563(.A(new_n673), .B1(new_n507), .B2(new_n533), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n750), .A2(new_n706), .A3(new_n709), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n727), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  AOI21_X1  g567(.A(new_n240), .B1(new_n725), .B2(new_n726), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n353), .A2(new_n243), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n360), .A2(new_n361), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n249), .B1(new_n757), .B2(new_n347), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n327), .A2(KEYINPUT80), .B1(new_n344), .B2(new_n343), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n330), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n756), .B(G469), .C1(new_n760), .C2(G902), .ZN(new_n761));
  AOI21_X1  g575(.A(G902), .B1(new_n346), .B2(new_n350), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT104), .B1(new_n762), .B2(new_n352), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n755), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n754), .A2(new_n674), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT41), .B(G113), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G15));
  NAND3_X1  g581(.A1(new_n754), .A2(new_n688), .A3(new_n764), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G116), .ZN(G18));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n581), .A2(new_n697), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n433), .B2(new_n456), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n763), .A2(new_n761), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n712), .A2(new_n244), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n706), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n770), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n775), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n725), .A2(new_n726), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(KEYINPUT105), .A3(new_n778), .A4(new_n771), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  OR2_X1    g595(.A1(new_n435), .A2(new_n389), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n449), .A2(new_n443), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n432), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(KEYINPUT106), .A3(new_n432), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n640), .A2(new_n241), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n773), .A2(new_n678), .A3(new_n739), .A4(new_n774), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G122), .ZN(G24));
  NAND2_X1  g607(.A1(new_n750), .A2(new_n709), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n775), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n787), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n718), .B1(new_n429), .B2(new_n231), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n697), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G125), .ZN(G27));
  INV_X1    g614(.A(KEYINPUT42), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n650), .B1(new_n631), .B2(new_n634), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n750), .A2(new_n709), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n457), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n750), .A2(new_n709), .A3(new_n802), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n805), .A4(new_n365), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G131), .ZN(G33));
  AND4_X1   g622(.A1(new_n685), .A2(new_n802), .A3(new_n687), .A4(new_n709), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n778), .A3(new_n241), .A4(new_n365), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n352), .B1(new_n715), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n815), .B(new_n816), .C1(new_n812), .C2(new_n715), .ZN(new_n817));
  NAND2_X1  g631(.A1(G469), .A2(G902), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT46), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n712), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(KEYINPUT46), .A3(new_n818), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n244), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(new_n742), .ZN(new_n823));
  INV_X1    g637(.A(new_n802), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n649), .A2(new_n672), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT43), .Z(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n698), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n640), .A2(new_n641), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n829), .B2(KEYINPUT44), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n823), .B(new_n830), .C1(KEYINPUT44), .C2(new_n829), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  XOR2_X1   g646(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n833));
  OR2_X1    g647(.A1(new_n822), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n778), .A2(new_n803), .A3(new_n241), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  NAND2_X1  g653(.A1(new_n573), .A2(new_n190), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n834), .A2(new_n836), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n773), .A2(new_n353), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n243), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n845), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n826), .A2(new_n574), .A3(new_n789), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n802), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n650), .A3(new_n747), .A4(new_n764), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n764), .A2(new_n802), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n826), .A2(new_n574), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n798), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n574), .A2(new_n738), .A3(new_n241), .A4(new_n853), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n649), .A3(new_n673), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n852), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT50), .B1(new_n851), .B2(KEYINPUT115), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT51), .B1(new_n850), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n754), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT48), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n750), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n573), .B(G953), .C1(new_n849), .C2(new_n777), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n850), .A2(new_n860), .A3(KEYINPUT51), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(KEYINPUT116), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(KEYINPUT116), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n796), .A2(new_n797), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n805), .A3(new_n365), .A4(new_n698), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n686), .A2(new_n709), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n648), .B2(new_n505), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n685), .A2(new_n802), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT110), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n685), .A2(new_n802), .A3(new_n875), .A4(KEYINPUT110), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n727), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n880), .A3(new_n810), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n804), .B2(new_n806), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n792), .A2(new_n700), .A3(new_n765), .A4(new_n768), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n828), .A2(new_n241), .A3(new_n365), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n507), .A2(new_n533), .A3(new_n572), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(KEYINPUT109), .C1(new_n649), .C2(new_n673), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT109), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n649), .A2(new_n887), .A3(new_n572), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n635), .A2(new_n579), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n884), .A2(new_n890), .B1(new_n457), .B2(new_n637), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n882), .A2(new_n892), .A3(KEYINPUT111), .A4(new_n780), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n506), .A2(G475), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n646), .A2(new_n529), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT90), .B1(new_n896), .B2(new_n231), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n572), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n684), .B2(new_n683), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n678), .A3(new_n773), .A4(new_n774), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n241), .B1(new_n433), .B2(new_n456), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n900), .A2(new_n901), .B1(new_n788), .B2(new_n790), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n773), .A2(new_n678), .A3(new_n750), .A4(new_n774), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n901), .A2(new_n903), .B1(new_n642), .B2(new_n699), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n243), .B1(new_n712), .B2(new_n716), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n240), .B(new_n907), .C1(new_n725), .C2(new_n726), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n643), .A2(new_n906), .B1(new_n908), .B2(new_n636), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n909), .A3(new_n780), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n873), .A2(new_n880), .A3(new_n810), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n807), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n894), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n893), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT113), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n739), .A2(new_n706), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n697), .A2(new_n709), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n737), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n872), .A2(new_n698), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n764), .A2(new_n750), .A3(new_n706), .A4(new_n709), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n752), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT52), .B1(new_n923), .B2(new_n731), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n705), .A2(KEYINPUT101), .A3(new_n710), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT52), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n915), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n927), .B2(new_n922), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n795), .A2(new_n798), .B1(new_n727), .B2(new_n751), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n731), .A2(KEYINPUT52), .A3(new_n932), .A4(new_n919), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(KEYINPUT113), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT53), .B1(new_n914), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n893), .A2(new_n913), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT53), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT112), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n928), .C1(new_n927), .C2(new_n922), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n931), .A2(KEYINPUT112), .A3(new_n933), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n936), .A2(KEYINPUT54), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n914), .B2(new_n935), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n910), .A2(new_n912), .ZN(new_n946));
  AND4_X1   g760(.A1(KEYINPUT53), .A2(new_n941), .A3(new_n946), .A4(new_n940), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n841), .B1(new_n871), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n843), .B(KEYINPUT49), .Z(new_n952));
  NOR4_X1   g766(.A1(new_n825), .A2(new_n650), .A3(new_n240), .A4(new_n244), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n738), .A3(new_n747), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(G75));
  NOR2_X1   g769(.A1(new_n190), .A2(G952), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n905), .A2(new_n780), .A3(new_n909), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT111), .B1(new_n958), .B2(new_n882), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n910), .A2(new_n912), .A3(new_n894), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n930), .B(new_n934), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n947), .B1(new_n961), .B2(new_n938), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n231), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT56), .B1(new_n963), .B2(G210), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n598), .A2(new_n600), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n606), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n957), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n964), .B2(new_n968), .ZN(G51));
  XOR2_X1   g784(.A(new_n818), .B(KEYINPUT57), .Z(new_n971));
  AND3_X1   g785(.A1(new_n931), .A2(KEYINPUT113), .A3(new_n933), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT113), .B1(new_n931), .B2(new_n933), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT53), .B1(new_n974), .B2(new_n937), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT54), .B1(new_n975), .B2(new_n947), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n949), .B2(KEYINPUT118), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT118), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n962), .B2(new_n945), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n760), .B(KEYINPUT119), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(G902), .B1(new_n975), .B2(new_n947), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(new_n817), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n956), .B1(new_n982), .B2(new_n984), .ZN(G54));
  NAND4_X1  g799(.A1(new_n963), .A2(KEYINPUT58), .A3(G475), .A4(new_n530), .ZN(new_n986));
  NAND2_X1  g800(.A1(KEYINPUT58), .A2(G475), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n529), .B(new_n528), .C1(new_n983), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n988), .A3(new_n957), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT120), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n986), .A2(new_n988), .A3(KEYINPUT120), .A4(new_n957), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(G60));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n936), .A2(KEYINPUT54), .A3(new_n942), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n975), .A2(KEYINPUT54), .A3(new_n947), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT121), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n995), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n977), .B2(new_n979), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n995), .B1(new_n943), .B2(new_n949), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1001), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT121), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AND4_X1   g821(.A1(new_n957), .A2(new_n1002), .A3(new_n1004), .A4(new_n1007), .ZN(G63));
  INV_X1    g822(.A(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G217), .A2(G902), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT60), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT122), .B1(new_n962), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT122), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1011), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1013), .B(new_n1014), .C1(new_n975), .C2(new_n947), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1012), .A2(new_n229), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n957), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n694), .A2(new_n695), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1009), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n1018), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1023), .A2(KEYINPUT61), .A3(new_n957), .A4(new_n1016), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1021), .A2(new_n1024), .ZN(G66));
  OAI21_X1  g839(.A(G953), .B1(new_n577), .B2(new_n603), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n958), .B2(G953), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT123), .ZN(new_n1028));
  INV_X1    g842(.A(G898), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n965), .B1(new_n1029), .B2(G953), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1028), .B(new_n1030), .ZN(G69));
  NAND2_X1  g845(.A1(new_n409), .A2(new_n446), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(new_n510), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(G900), .B2(G953), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n838), .A2(new_n807), .A3(new_n810), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n731), .A2(new_n932), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n831), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n823), .A2(new_n754), .A3(new_n916), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1034), .B1(new_n1039), .B2(G953), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT125), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT62), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n748), .A2(new_n1043), .A3(new_n1036), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n743), .A2(new_n824), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n1045), .A2(new_n754), .A3(new_n886), .A4(new_n888), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n831), .A2(new_n838), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1043), .B1(new_n748), .B2(new_n1036), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1033), .B1(new_n1049), .B2(G953), .ZN(new_n1050));
  OAI211_X1 g864(.A(KEYINPUT125), .B(new_n1034), .C1(new_n1039), .C2(G953), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1042), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1053), .B(KEYINPUT124), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1040), .A2(new_n1050), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1054), .A2(new_n1056), .ZN(G72));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  OAI21_X1  g873(.A(new_n1059), .B1(new_n1039), .B2(new_n910), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n722), .A2(new_n414), .ZN(new_n1061));
  XOR2_X1   g875(.A(new_n1061), .B(KEYINPUT127), .Z(new_n1062));
  NAND2_X1  g876(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n936), .A2(new_n942), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1059), .B1(new_n439), .B2(new_n412), .ZN(new_n1065));
  OAI211_X1 g879(.A(new_n1063), .B(new_n957), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g880(.A(new_n1059), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1067), .B1(new_n1049), .B2(new_n958), .ZN(new_n1068));
  XOR2_X1   g882(.A(new_n1068), .B(KEYINPUT126), .Z(new_n1069));
  NOR2_X1   g883(.A1(new_n722), .A2(new_n414), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(G57));
endmodule


