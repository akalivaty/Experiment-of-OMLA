

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742;

  NAND2_X1 U376 ( .A1(n643), .A2(n644), .ZN(n646) );
  XNOR2_X1 U377 ( .A(n379), .B(G146), .ZN(n465) );
  NOR2_X1 U378 ( .A1(n735), .A2(n742), .ZN(n561) );
  XNOR2_X1 U379 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U380 ( .A(n482), .B(n481), .ZN(n493) );
  XNOR2_X1 U381 ( .A(n465), .B(n369), .ZN(n466) );
  XNOR2_X1 U382 ( .A(n370), .B(KEYINPUT17), .ZN(n369) );
  INV_X2 U383 ( .A(G128), .ZN(n386) );
  INV_X2 U384 ( .A(KEYINPUT64), .ZN(n391) );
  BUF_X1 U385 ( .A(n697), .Z(n354) );
  XNOR2_X1 U386 ( .A(n375), .B(n727), .ZN(n697) );
  XNOR2_X2 U387 ( .A(n509), .B(KEYINPUT32), .ZN(n738) );
  XNOR2_X1 U388 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X2 U389 ( .A(n463), .B(n385), .ZN(n482) );
  XNOR2_X1 U390 ( .A(n454), .B(n453), .ZN(n487) );
  XNOR2_X1 U391 ( .A(G119), .B(KEYINPUT3), .ZN(n453) );
  XOR2_X1 U392 ( .A(G146), .B(n483), .Z(n496) );
  NAND2_X1 U393 ( .A1(n439), .A2(G221), .ZN(n396) );
  NAND2_X1 U394 ( .A1(n706), .A2(n364), .ZN(n407) );
  XOR2_X1 U395 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n429) );
  XOR2_X1 U396 ( .A(G131), .B(G143), .Z(n427) );
  XNOR2_X1 U397 ( .A(n465), .B(n378), .ZN(n728) );
  INV_X1 U398 ( .A(KEYINPUT10), .ZN(n378) );
  XOR2_X1 U399 ( .A(KEYINPUT76), .B(G104), .Z(n498) );
  INV_X1 U400 ( .A(n644), .ZN(n411) );
  XNOR2_X1 U401 ( .A(n492), .B(n491), .ZN(n616) );
  XNOR2_X1 U402 ( .A(G110), .B(G107), .ZN(n719) );
  XOR2_X1 U403 ( .A(KEYINPUT23), .B(G119), .Z(n421) );
  XNOR2_X1 U404 ( .A(G110), .B(G128), .ZN(n420) );
  INV_X1 U405 ( .A(KEYINPUT84), .ZN(n399) );
  XNOR2_X1 U406 ( .A(n418), .B(n397), .ZN(n439) );
  INV_X1 U407 ( .A(KEYINPUT8), .ZN(n397) );
  XNOR2_X1 U408 ( .A(n551), .B(n550), .ZN(n683) );
  NOR2_X1 U409 ( .A1(n546), .A2(n566), .ZN(n547) );
  INV_X1 U410 ( .A(n555), .ZN(n652) );
  XNOR2_X1 U411 ( .A(n381), .B(n380), .ZN(n524) );
  XNOR2_X1 U412 ( .A(KEYINPUT13), .B(G475), .ZN(n380) );
  OR2_X1 U413 ( .A1(n703), .A2(G902), .ZN(n381) );
  INV_X1 U414 ( .A(KEYINPUT0), .ZN(n412) );
  XNOR2_X1 U415 ( .A(n479), .B(KEYINPUT25), .ZN(n371) );
  NOR2_X1 U416 ( .A1(n406), .A2(n711), .ZN(n405) );
  NOR2_X1 U417 ( .A1(n361), .A2(G472), .ZN(n406) );
  BUF_X1 U418 ( .A(n459), .Z(n372) );
  NAND2_X1 U419 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U420 ( .A(KEYINPUT18), .ZN(n370) );
  INV_X1 U421 ( .A(G125), .ZN(n379) );
  INV_X1 U422 ( .A(KEYINPUT4), .ZN(n385) );
  XNOR2_X1 U423 ( .A(G131), .B(G134), .ZN(n481) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n488) );
  XNOR2_X1 U425 ( .A(G137), .B(KEYINPUT97), .ZN(n484) );
  XNOR2_X1 U426 ( .A(G116), .B(G107), .ZN(n434) );
  XNOR2_X1 U427 ( .A(n455), .B(n357), .ZN(n414) );
  XOR2_X1 U428 ( .A(n581), .B(KEYINPUT38), .Z(n660) );
  XNOR2_X1 U429 ( .A(n433), .B(n356), .ZN(n703) );
  XNOR2_X1 U430 ( .A(G140), .B(G113), .ZN(n426) );
  INV_X1 U431 ( .A(G953), .ZN(n475) );
  XNOR2_X1 U432 ( .A(n501), .B(n496), .ZN(n375) );
  NOR2_X1 U433 ( .A1(n388), .A2(n553), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n543), .B(n389), .ZN(n388) );
  XNOR2_X1 U435 ( .A(n544), .B(KEYINPUT106), .ZN(n389) );
  BUF_X1 U436 ( .A(n535), .Z(n581) );
  OR2_X1 U437 ( .A1(n616), .A2(G902), .ZN(n390) );
  XNOR2_X1 U438 ( .A(n555), .B(n368), .ZN(n582) );
  INV_X1 U439 ( .A(KEYINPUT6), .ZN(n368) );
  XNOR2_X1 U440 ( .A(n367), .B(n360), .ZN(n520) );
  NOR2_X1 U441 ( .A1(n662), .A2(n411), .ZN(n410) );
  XNOR2_X1 U442 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U443 ( .A(n398), .B(n396), .ZN(n425) );
  NAND2_X1 U444 ( .A1(n683), .A2(n563), .ZN(n560) );
  NOR2_X1 U445 ( .A1(n408), .A2(n404), .ZN(n617) );
  NAND2_X1 U446 ( .A1(n407), .A2(n405), .ZN(n404) );
  INV_X1 U447 ( .A(KEYINPUT60), .ZN(n392) );
  AND2_X1 U448 ( .A1(n382), .A2(n601), .ZN(n355) );
  XOR2_X1 U449 ( .A(n427), .B(n426), .Z(n356) );
  XNOR2_X1 U450 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n357) );
  XOR2_X1 U451 ( .A(KEYINPUT70), .B(G472), .Z(n358) );
  OR2_X1 U452 ( .A1(n575), .A2(n532), .ZN(n359) );
  XOR2_X1 U453 ( .A(KEYINPUT71), .B(KEYINPUT22), .Z(n360) );
  XOR2_X1 U454 ( .A(n616), .B(n615), .Z(n361) );
  XOR2_X1 U455 ( .A(n705), .B(n704), .Z(n362) );
  XOR2_X1 U456 ( .A(KEYINPUT45), .B(KEYINPUT88), .Z(n363) );
  AND2_X1 U457 ( .A1(n361), .A2(G472), .ZN(n364) );
  NOR2_X1 U458 ( .A1(n372), .A2(G952), .ZN(n711) );
  INV_X1 U459 ( .A(n711), .ZN(n409) );
  XNOR2_X2 U460 ( .A(n480), .B(n371), .ZN(n643) );
  NOR2_X1 U461 ( .A1(n365), .A2(G953), .ZN(n690) );
  XNOR2_X1 U462 ( .A(n689), .B(n688), .ZN(n365) );
  XNOR2_X1 U463 ( .A(n383), .B(n592), .ZN(n382) );
  XNOR2_X1 U464 ( .A(n419), .B(n399), .ZN(n398) );
  NAND2_X1 U465 ( .A1(n545), .A2(n387), .ZN(n566) );
  XNOR2_X2 U466 ( .A(n494), .B(n495), .ZN(n727) );
  AND2_X2 U467 ( .A1(n736), .A2(n738), .ZN(n376) );
  XNOR2_X1 U468 ( .A(n414), .B(n487), .ZN(n457) );
  NAND2_X1 U469 ( .A1(n366), .A2(n458), .ZN(n417) );
  NAND2_X1 U470 ( .A1(n721), .A2(n499), .ZN(n366) );
  NAND2_X1 U471 ( .A1(n529), .A2(n410), .ZN(n367) );
  XNOR2_X2 U472 ( .A(n518), .B(KEYINPUT35), .ZN(n736) );
  NOR2_X2 U473 ( .A1(n697), .A2(G902), .ZN(n503) );
  XNOR2_X1 U474 ( .A(n471), .B(KEYINPUT19), .ZN(n562) );
  AND2_X2 U475 ( .A1(G224), .A2(n459), .ZN(n461) );
  XNOR2_X2 U476 ( .A(n390), .B(n358), .ZN(n555) );
  NOR2_X2 U477 ( .A1(n520), .A2(n643), .ZN(n508) );
  XOR2_X2 U478 ( .A(G122), .B(G104), .Z(n455) );
  INV_X1 U479 ( .A(n457), .ZN(n721) );
  XNOR2_X1 U480 ( .A(n416), .B(n464), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n415), .B(n417), .ZN(n691) );
  NAND2_X1 U482 ( .A1(n535), .A2(n659), .ZN(n471) );
  XNOR2_X2 U483 ( .A(n470), .B(n469), .ZN(n535) );
  XNOR2_X1 U484 ( .A(n403), .B(n402), .ZN(n401) );
  XNOR2_X1 U485 ( .A(n466), .B(n462), .ZN(n416) );
  NAND2_X1 U486 ( .A1(n562), .A2(n477), .ZN(n413) );
  XNOR2_X1 U487 ( .A(n373), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U488 ( .A1(n696), .A2(n711), .ZN(n373) );
  INV_X1 U489 ( .A(n587), .ZN(n510) );
  AND2_X2 U490 ( .A1(n374), .A2(n587), .ZN(n527) );
  XNOR2_X2 U491 ( .A(n559), .B(n504), .ZN(n587) );
  INV_X1 U492 ( .A(n646), .ZN(n374) );
  NAND2_X1 U493 ( .A1(n377), .A2(n376), .ZN(n403) );
  INV_X1 U494 ( .A(n737), .ZN(n377) );
  NAND2_X1 U495 ( .A1(n574), .A2(n384), .ZN(n383) );
  AND2_X1 U496 ( .A1(n591), .A2(n573), .ZN(n384) );
  XNOR2_X2 U497 ( .A(n386), .B(G143), .ZN(n463) );
  XNOR2_X2 U498 ( .A(n391), .B(G953), .ZN(n459) );
  XNOR2_X1 U499 ( .A(n393), .B(n392), .ZN(G60) );
  NAND2_X1 U500 ( .A1(n394), .A2(n409), .ZN(n393) );
  XNOR2_X1 U501 ( .A(n395), .B(n362), .ZN(n394) );
  NAND2_X1 U502 ( .A1(n706), .A2(G475), .ZN(n395) );
  AND2_X2 U503 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X2 U504 ( .A(n503), .B(n502), .ZN(n559) );
  NOR2_X2 U505 ( .A1(n715), .A2(n603), .ZN(n534) );
  XNOR2_X1 U506 ( .A(n515), .B(n514), .ZN(n517) );
  XNOR2_X1 U507 ( .A(n425), .B(n424), .ZN(n611) );
  XNOR2_X2 U508 ( .A(n400), .B(n363), .ZN(n715) );
  NAND2_X1 U509 ( .A1(n401), .A2(n533), .ZN(n400) );
  INV_X1 U510 ( .A(KEYINPUT44), .ZN(n402) );
  NOR2_X1 U511 ( .A1(n706), .A2(n361), .ZN(n408) );
  AND2_X4 U512 ( .A1(n609), .A2(n681), .ZN(n706) );
  XNOR2_X2 U513 ( .A(n413), .B(n412), .ZN(n529) );
  XNOR2_X1 U514 ( .A(n695), .B(n694), .ZN(n696) );
  INV_X1 U515 ( .A(n575), .ZN(n577) );
  NOR2_X1 U516 ( .A1(n633), .A2(n635), .ZN(n664) );
  INV_X1 U517 ( .A(n641), .ZN(n589) );
  INV_X1 U518 ( .A(n642), .ZN(n600) );
  XNOR2_X1 U519 ( .A(KEYINPUT48), .B(KEYINPUT89), .ZN(n592) );
  NOR2_X1 U520 ( .A1(n740), .A2(n600), .ZN(n601) );
  INV_X1 U521 ( .A(KEYINPUT41), .ZN(n550) );
  INV_X1 U522 ( .A(KEYINPUT123), .ZN(n613) );
  XOR2_X2 U523 ( .A(G137), .B(G140), .Z(n495) );
  XOR2_X1 U524 ( .A(n495), .B(KEYINPUT94), .Z(n419) );
  NAND2_X1 U525 ( .A1(n459), .A2(G234), .ZN(n418) );
  XNOR2_X1 U526 ( .A(n728), .B(KEYINPUT24), .ZN(n423) );
  XNOR2_X1 U527 ( .A(n421), .B(n420), .ZN(n422) );
  NAND2_X1 U528 ( .A1(n488), .A2(G214), .ZN(n428) );
  XNOR2_X1 U529 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U530 ( .A(n430), .B(KEYINPUT11), .Z(n432) );
  XNOR2_X1 U531 ( .A(n728), .B(n455), .ZN(n431) );
  XNOR2_X1 U532 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U533 ( .A(G134), .B(KEYINPUT9), .ZN(n443) );
  XNOR2_X1 U534 ( .A(n434), .B(n463), .ZN(n438) );
  XOR2_X1 U535 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n436) );
  XNOR2_X1 U536 ( .A(G122), .B(KEYINPUT7), .ZN(n435) );
  XNOR2_X1 U537 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U538 ( .A(n438), .B(n437), .Z(n441) );
  NAND2_X1 U539 ( .A1(G217), .A2(n439), .ZN(n440) );
  XNOR2_X1 U540 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n443), .B(n442), .ZN(n708) );
  NOR2_X1 U542 ( .A1(n708), .A2(G902), .ZN(n444) );
  XNOR2_X1 U543 ( .A(n444), .B(G478), .ZN(n522) );
  NAND2_X1 U544 ( .A1(n524), .A2(n522), .ZN(n662) );
  XOR2_X1 U545 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n448) );
  XOR2_X1 U546 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n446) );
  XOR2_X1 U547 ( .A(G902), .B(KEYINPUT15), .Z(n467) );
  INV_X1 U548 ( .A(n467), .ZN(n603) );
  NAND2_X1 U549 ( .A1(G234), .A2(n603), .ZN(n445) );
  XNOR2_X1 U550 ( .A(n446), .B(n445), .ZN(n478) );
  NAND2_X1 U551 ( .A1(n478), .A2(G221), .ZN(n447) );
  XNOR2_X1 U552 ( .A(n448), .B(n447), .ZN(n644) );
  OR2_X1 U553 ( .A1(G237), .A2(G902), .ZN(n468) );
  NAND2_X1 U554 ( .A1(G214), .A2(n468), .ZN(n659) );
  INV_X1 U555 ( .A(G116), .ZN(n449) );
  NAND2_X1 U556 ( .A1(G113), .A2(n449), .ZN(n452) );
  INV_X1 U557 ( .A(G113), .ZN(n450) );
  NAND2_X1 U558 ( .A1(n450), .A2(G116), .ZN(n451) );
  NAND2_X1 U559 ( .A1(n452), .A2(n451), .ZN(n454) );
  XNOR2_X1 U560 ( .A(KEYINPUT69), .B(n719), .ZN(n499) );
  INV_X1 U561 ( .A(n499), .ZN(n456) );
  NAND2_X1 U562 ( .A1(n457), .A2(n456), .ZN(n458) );
  INV_X1 U563 ( .A(KEYINPUT92), .ZN(n460) );
  XOR2_X1 U564 ( .A(KEYINPUT67), .B(G101), .Z(n483) );
  XNOR2_X1 U565 ( .A(n482), .B(n483), .ZN(n464) );
  NOR2_X2 U566 ( .A1(n691), .A2(n467), .ZN(n470) );
  NAND2_X1 U567 ( .A1(G210), .A2(n468), .ZN(n469) );
  NAND2_X1 U568 ( .A1(G237), .A2(G234), .ZN(n472) );
  XNOR2_X1 U569 ( .A(n472), .B(KEYINPUT14), .ZN(n473) );
  AND2_X1 U570 ( .A1(G952), .A2(n473), .ZN(n673) );
  NAND2_X1 U571 ( .A1(n673), .A2(n475), .ZN(n536) );
  NAND2_X1 U572 ( .A1(n473), .A2(G902), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n474), .B(KEYINPUT93), .ZN(n537) );
  NOR2_X1 U574 ( .A1(G898), .A2(n475), .ZN(n723) );
  NAND2_X1 U575 ( .A1(n537), .A2(n723), .ZN(n476) );
  NAND2_X1 U576 ( .A1(n536), .A2(n476), .ZN(n477) );
  NOR2_X1 U577 ( .A1(G902), .A2(n611), .ZN(n480) );
  NAND2_X1 U578 ( .A1(n478), .A2(G217), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n493), .B(n496), .ZN(n492) );
  XOR2_X1 U580 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n485) );
  XNOR2_X1 U581 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U582 ( .A(n487), .B(n486), .Z(n490) );
  NAND2_X1 U583 ( .A1(n488), .A2(G210), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U585 ( .A(n493), .ZN(n494) );
  NAND2_X1 U586 ( .A1(G227), .A2(n459), .ZN(n497) );
  XNOR2_X1 U587 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U588 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U589 ( .A(KEYINPUT68), .B(G469), .ZN(n502) );
  XNOR2_X1 U590 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n504) );
  NOR2_X1 U591 ( .A1(n652), .A2(n587), .ZN(n505) );
  NAND2_X1 U592 ( .A1(n508), .A2(n505), .ZN(n506) );
  XNOR2_X1 U593 ( .A(KEYINPUT103), .B(n506), .ZN(n737) );
  INV_X1 U594 ( .A(n582), .ZN(n511) );
  NOR2_X1 U595 ( .A1(n510), .A2(n511), .ZN(n507) );
  NAND2_X1 U596 ( .A1(n508), .A2(n507), .ZN(n509) );
  NAND2_X1 U597 ( .A1(n527), .A2(n511), .ZN(n513) );
  XNOR2_X1 U598 ( .A(KEYINPUT90), .B(KEYINPUT33), .ZN(n512) );
  XNOR2_X2 U599 ( .A(n513), .B(n512), .ZN(n658) );
  NAND2_X1 U600 ( .A1(n529), .A2(n658), .ZN(n515) );
  XNOR2_X1 U601 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n514) );
  OR2_X1 U602 ( .A1(n524), .A2(n522), .ZN(n565) );
  INV_X1 U603 ( .A(n565), .ZN(n516) );
  NAND2_X1 U604 ( .A1(n582), .A2(n643), .ZN(n519) );
  NOR2_X1 U605 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U606 ( .A1(n521), .A2(n510), .ZN(n618) );
  INV_X1 U607 ( .A(n522), .ZN(n523) );
  NOR2_X1 U608 ( .A1(n523), .A2(n524), .ZN(n633) );
  NAND2_X1 U609 ( .A1(n524), .A2(n523), .ZN(n626) );
  INV_X1 U610 ( .A(n626), .ZN(n635) );
  XOR2_X1 U611 ( .A(KEYINPUT83), .B(n664), .Z(n575) );
  INV_X1 U612 ( .A(n529), .ZN(n526) );
  NOR2_X1 U613 ( .A1(n559), .A2(n646), .ZN(n545) );
  NAND2_X1 U614 ( .A1(n555), .A2(n545), .ZN(n525) );
  NOR2_X1 U615 ( .A1(n526), .A2(n525), .ZN(n621) );
  XOR2_X1 U616 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n531) );
  AND2_X1 U617 ( .A1(n527), .A2(n652), .ZN(n528) );
  XNOR2_X1 U618 ( .A(KEYINPUT98), .B(n528), .ZN(n654) );
  NAND2_X1 U619 ( .A1(n654), .A2(n529), .ZN(n530) );
  XNOR2_X1 U620 ( .A(n531), .B(n530), .ZN(n636) );
  NOR2_X1 U621 ( .A1(n621), .A2(n636), .ZN(n532) );
  AND2_X1 U622 ( .A1(n618), .A2(n359), .ZN(n533) );
  XNOR2_X1 U623 ( .A(n534), .B(KEYINPUT86), .ZN(n602) );
  INV_X1 U624 ( .A(n660), .ZN(n546) );
  INV_X1 U625 ( .A(n536), .ZN(n541) );
  INV_X1 U626 ( .A(n372), .ZN(n538) );
  NAND2_X1 U627 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U628 ( .A1(G900), .A2(n539), .ZN(n540) );
  NOR2_X1 U629 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U630 ( .A(KEYINPUT78), .B(n542), .ZN(n553) );
  XOR2_X1 U631 ( .A(KEYINPUT30), .B(KEYINPUT107), .Z(n544) );
  NAND2_X1 U632 ( .A1(n652), .A2(n659), .ZN(n543) );
  XOR2_X1 U633 ( .A(KEYINPUT39), .B(n547), .Z(n599) );
  AND2_X1 U634 ( .A1(n633), .A2(n599), .ZN(n549) );
  XNOR2_X1 U635 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n548) );
  XNOR2_X1 U636 ( .A(n549), .B(n548), .ZN(n735) );
  NAND2_X1 U637 ( .A1(n660), .A2(n659), .ZN(n663) );
  NOR2_X1 U638 ( .A1(n663), .A2(n662), .ZN(n551) );
  XNOR2_X1 U639 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n552) );
  XNOR2_X1 U640 ( .A(n552), .B(KEYINPUT108), .ZN(n557) );
  NOR2_X1 U641 ( .A1(n643), .A2(n553), .ZN(n554) );
  NAND2_X1 U642 ( .A1(n644), .A2(n554), .ZN(n585) );
  NOR2_X1 U643 ( .A1(n555), .A2(n585), .ZN(n556) );
  XNOR2_X1 U644 ( .A(n557), .B(n556), .ZN(n558) );
  NOR2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n563) );
  XOR2_X1 U646 ( .A(KEYINPUT42), .B(n560), .Z(n742) );
  XNOR2_X1 U647 ( .A(n561), .B(KEYINPUT46), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n563), .A2(n562), .ZN(n630) );
  NAND2_X1 U649 ( .A1(KEYINPUT47), .A2(n630), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n564), .B(KEYINPUT82), .ZN(n571) );
  NAND2_X1 U651 ( .A1(KEYINPUT47), .A2(n664), .ZN(n568) );
  NOR2_X1 U652 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U653 ( .A1(n581), .A2(n567), .ZN(n629) );
  NAND2_X1 U654 ( .A1(n568), .A2(n629), .ZN(n569) );
  XNOR2_X1 U655 ( .A(KEYINPUT79), .B(n569), .ZN(n570) );
  NAND2_X1 U656 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n572), .B(KEYINPUT81), .ZN(n573) );
  INV_X1 U658 ( .A(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U659 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U660 ( .A(n578), .B(KEYINPUT74), .ZN(n579) );
  NOR2_X1 U661 ( .A1(n630), .A2(n579), .ZN(n580) );
  XOR2_X1 U662 ( .A(KEYINPUT73), .B(n580), .Z(n590) );
  INV_X1 U663 ( .A(n581), .ZN(n596) );
  INV_X1 U664 ( .A(n633), .ZN(n631) );
  NOR2_X1 U665 ( .A1(n582), .A2(n631), .ZN(n583) );
  NAND2_X1 U666 ( .A1(n583), .A2(n659), .ZN(n584) );
  OR2_X1 U667 ( .A1(n585), .A2(n584), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n596), .A2(n593), .ZN(n586) );
  XNOR2_X1 U669 ( .A(KEYINPUT36), .B(n586), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n641) );
  NOR2_X1 U671 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U672 ( .A(n593), .B(KEYINPUT104), .Z(n594) );
  NAND2_X1 U673 ( .A1(n594), .A2(n510), .ZN(n595) );
  XNOR2_X1 U674 ( .A(n595), .B(KEYINPUT43), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U676 ( .A(KEYINPUT105), .B(n598), .ZN(n740) );
  NAND2_X1 U677 ( .A1(n599), .A2(n635), .ZN(n642) );
  NAND2_X1 U678 ( .A1(n602), .A2(n355), .ZN(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT87), .B(n603), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n604), .A2(KEYINPUT2), .ZN(n605) );
  XNOR2_X1 U681 ( .A(KEYINPUT66), .B(n605), .ZN(n606) );
  INV_X1 U682 ( .A(KEYINPUT2), .ZN(n675) );
  NOR2_X1 U683 ( .A1(n715), .A2(n675), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n608), .A2(n355), .ZN(n681) );
  NAND2_X1 U685 ( .A1(n706), .A2(G217), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(n611), .ZN(n612) );
  NOR2_X2 U687 ( .A1(n612), .A2(n711), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(n613), .ZN(G66) );
  XOR2_X1 U689 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n615) );
  XOR2_X1 U690 ( .A(KEYINPUT63), .B(n617), .Z(G57) );
  XNOR2_X1 U691 ( .A(G101), .B(n618), .ZN(G3) );
  NAND2_X1 U692 ( .A1(n621), .A2(n633), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT112), .ZN(n620) );
  XNOR2_X1 U694 ( .A(G104), .B(n620), .ZN(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n623) );
  NAND2_X1 U696 ( .A1(n621), .A2(n635), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(n625) );
  XOR2_X1 U698 ( .A(G107), .B(KEYINPUT27), .Z(n624) );
  XNOR2_X1 U699 ( .A(n625), .B(n624), .ZN(G9) );
  NOR2_X1 U700 ( .A1(n630), .A2(n626), .ZN(n628) );
  XNOR2_X1 U701 ( .A(G128), .B(KEYINPUT29), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n628), .B(n627), .ZN(G30) );
  XNOR2_X1 U703 ( .A(G143), .B(n629), .ZN(G45) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U705 ( .A(G146), .B(n632), .Z(G48) );
  NAND2_X1 U706 ( .A1(n636), .A2(n633), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(G113), .ZN(G15) );
  XOR2_X1 U708 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n638) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U711 ( .A(G116), .B(n639), .ZN(G18) );
  XOR2_X1 U712 ( .A(G125), .B(KEYINPUT37), .Z(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n642), .ZN(G36) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(KEYINPUT49), .B(n645), .ZN(n650) );
  XOR2_X1 U717 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n648) );
  NAND2_X1 U718 ( .A1(n646), .A2(n510), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U723 ( .A(KEYINPUT51), .B(n655), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n656), .A2(n683), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT118), .B(n657), .Z(n670) );
  INV_X1 U726 ( .A(n658), .ZN(n668) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U733 ( .A(KEYINPUT52), .B(n671), .Z(n672) );
  NAND2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U735 ( .A(KEYINPUT119), .B(n674), .ZN(n687) );
  XOR2_X1 U736 ( .A(KEYINPUT80), .B(n675), .Z(n678) );
  INV_X1 U737 ( .A(n678), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n715), .A2(n676), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n677), .B(KEYINPUT85), .ZN(n680) );
  NOR2_X1 U740 ( .A1(n678), .A2(n355), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U743 ( .A1(n683), .A2(n658), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n689) );
  INV_X1 U746 ( .A(KEYINPUT120), .ZN(n688) );
  XNOR2_X1 U747 ( .A(KEYINPUT53), .B(n690), .ZN(G75) );
  NAND2_X1 U748 ( .A1(n706), .A2(G210), .ZN(n695) );
  BUF_X1 U749 ( .A(n691), .Z(n693) );
  XOR2_X1 U750 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n692) );
  XNOR2_X1 U751 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n354), .B(KEYINPUT57), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U754 ( .A1(n706), .A2(G469), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n711), .A2(n702), .ZN(G54) );
  INV_X1 U757 ( .A(n703), .ZN(n705) );
  XOR2_X1 U758 ( .A(KEYINPUT59), .B(KEYINPUT91), .Z(n704) );
  NAND2_X1 U759 ( .A1(n706), .A2(G478), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT122), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n711), .A2(n710), .ZN(G63) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n712) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n712), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n713), .A2(G898), .ZN(n714) );
  XOR2_X1 U766 ( .A(KEYINPUT124), .B(n714), .Z(n717) );
  NOR2_X1 U767 ( .A1(G953), .A2(n715), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n726) );
  XOR2_X1 U769 ( .A(G101), .B(KEYINPUT125), .Z(n718) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U771 ( .A(n721), .B(n720), .Z(n722) );
  NOR2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U773 ( .A(KEYINPUT126), .B(n724), .Z(n725) );
  XNOR2_X1 U774 ( .A(n726), .B(n725), .ZN(G69) );
  XOR2_X1 U775 ( .A(n728), .B(n727), .Z(n730) );
  XOR2_X1 U776 ( .A(n730), .B(n355), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n372), .ZN(n734) );
  XNOR2_X1 U778 ( .A(G227), .B(n730), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(G72) );
  XOR2_X1 U782 ( .A(n735), .B(G131), .Z(G33) );
  XNOR2_X1 U783 ( .A(G122), .B(n736), .ZN(G24) );
  XOR2_X1 U784 ( .A(n737), .B(G110), .Z(G12) );
  XOR2_X1 U785 ( .A(G119), .B(n738), .Z(n739) );
  XNOR2_X1 U786 ( .A(KEYINPUT127), .B(n739), .ZN(G21) );
  XOR2_X1 U787 ( .A(G140), .B(n740), .Z(n741) );
  XNOR2_X1 U788 ( .A(KEYINPUT116), .B(n741), .ZN(G42) );
  XOR2_X1 U789 ( .A(G137), .B(n742), .Z(G39) );
endmodule

