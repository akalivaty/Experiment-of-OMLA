//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G355));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n210), .B(new_n216), .C1(G58), .C2(G232), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G1), .B2(G20), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT66), .B(KEYINPUT1), .Z(new_n219));
  XNOR2_X1  g0019(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n203), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G1), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n225), .A2(new_n222), .A3(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NOR3_X1   g0028(.A1(new_n220), .A2(new_n224), .A3(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  INV_X1    g0032(.A(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n209), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n208), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n223), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(new_n225), .B2(G20), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G50), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n225), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  OR2_X1    g0054(.A1(KEYINPUT8), .A2(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT8), .A2(G58), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n257), .A2(KEYINPUT71), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n201), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n222), .B1(new_n261), .B2(new_n202), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT71), .B1(new_n257), .B2(new_n259), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n248), .A2(new_n223), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n251), .B1(G50), .B2(new_n252), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT67), .B(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n225), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(KEYINPUT70), .A3(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(G223), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(G222), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n283), .C1(new_n284), .C2(new_n279), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n272), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n223), .ZN(new_n291));
  NAND3_X1  g0091(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n294), .B2(new_n269), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n293), .A2(KEYINPUT69), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT69), .B1(new_n293), .B2(new_n296), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(KEYINPUT72), .B(new_n266), .C1(new_n302), .C2(G169), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT72), .ZN(new_n304));
  INV_X1    g0104(.A(new_n266), .ZN(new_n305));
  AOI21_X1  g0105(.A(G169), .B1(new_n287), .B2(new_n300), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n303), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n301), .A2(G200), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n252), .A2(G50), .ZN(new_n314));
  INV_X1    g0114(.A(new_n264), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n249), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(KEYINPUT9), .A3(new_n251), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n266), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n287), .A2(G190), .A3(new_n300), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n313), .A2(new_n317), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n301), .A2(G200), .B1(new_n266), .B2(new_n318), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(new_n317), .A4(new_n320), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT73), .A4(new_n309), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n312), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n297), .A2(new_n298), .A3(new_n213), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n272), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT69), .ZN(new_n335));
  AND3_X1   g0135(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT68), .B1(G33), .B2(G41), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n336), .A2(new_n337), .A3(new_n223), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n338), .B2(new_n295), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n293), .A2(new_n296), .A3(KEYINPUT69), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(G238), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n279), .A2(new_n282), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n344), .B1(new_n253), .B2(new_n214), .C1(new_n345), .C2(new_n233), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n286), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n331), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n346), .A2(new_n286), .ZN(new_n349));
  AOI211_X1 g0149(.A(KEYINPUT13), .B(new_n349), .C1(new_n334), .C2(new_n342), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n330), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n341), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT74), .B1(new_n341), .B2(new_n271), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT13), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n331), .B(new_n347), .C1(new_n353), .C2(new_n354), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(G179), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n330), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n352), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n254), .A2(G77), .B1(new_n258), .B2(G50), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n222), .B2(G68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n249), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT11), .ZN(new_n366));
  INV_X1    g0166(.A(new_n252), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n212), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT12), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n250), .A2(G68), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT75), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n255), .A2(new_n256), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n252), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n250), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n273), .A2(new_n275), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT77), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n279), .B2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT7), .A4(new_n222), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n242), .A2(new_n212), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n386), .B2(new_n202), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n258), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT16), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n381), .A2(new_n378), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT16), .B(new_n390), .C1(new_n392), .C2(new_n212), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n249), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n376), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n273), .A2(new_n275), .A3(G226), .A4(G1698), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n273), .A2(new_n275), .A3(G223), .A4(new_n282), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n286), .B1(new_n270), .B2(new_n225), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n293), .A2(new_n296), .A3(G232), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n400), .A2(G179), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n329), .B1(new_n400), .B2(new_n401), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n395), .A2(KEYINPUT18), .A3(new_n404), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n389), .B1(new_n384), .B2(G68), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n249), .B(new_n393), .C1(new_n409), .C2(KEYINPUT16), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n400), .A2(new_n411), .A3(new_n401), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n399), .A2(new_n286), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n413), .A2(new_n401), .A3(new_n271), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(G200), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n376), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT17), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n410), .A2(new_n418), .A3(new_n415), .A4(new_n376), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n407), .A2(new_n408), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n278), .A2(new_n280), .A3(G238), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n279), .A2(G232), .A3(new_n282), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n377), .A2(G107), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n286), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n299), .A2(G244), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n271), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n329), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n308), .A3(new_n426), .A4(new_n271), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n252), .A2(G77), .ZN(new_n430));
  INV_X1    g0230(.A(new_n374), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n432));
  XOR2_X1   g0232(.A(KEYINPUT15), .B(G87), .Z(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n254), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n430), .B1(new_n436), .B2(new_n249), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n250), .A2(G77), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n428), .A2(new_n429), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n427), .A2(G200), .ZN(new_n441));
  INV_X1    g0241(.A(new_n439), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n272), .B1(new_n424), .B2(new_n286), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G190), .A3(new_n426), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n420), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(G200), .B1(new_n348), .B2(new_n350), .ZN(new_n447));
  INV_X1    g0247(.A(new_n372), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n356), .A2(G190), .A3(new_n357), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n328), .A2(new_n373), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT24), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n279), .A2(KEYINPUT83), .A3(new_n222), .A4(G87), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT22), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n377), .A2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT84), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(KEYINPUT83), .A3(new_n458), .A4(G87), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT23), .B1(new_n464), .B2(G20), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(KEYINPUT23), .A3(G20), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n465), .A2(new_n467), .B1(new_n435), .B2(new_n208), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n452), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  AOI211_X1 g0270(.A(KEYINPUT24), .B(new_n468), .C1(new_n456), .C2(new_n462), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n249), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n367), .A2(KEYINPUT25), .A3(new_n464), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n367), .B2(new_n464), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n225), .A2(G33), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n265), .A2(new_n252), .A3(new_n476), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n464), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n269), .A2(G1), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n294), .A2(KEYINPUT5), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n481), .C1(new_n268), .C2(KEYINPUT5), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n482), .A2(new_n293), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G264), .ZN(new_n484));
  INV_X1    g0284(.A(G250), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n345), .A2(new_n485), .B1(new_n215), .B2(new_n276), .ZN(new_n486));
  INV_X1    g0286(.A(G294), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n253), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n286), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n480), .ZN(new_n490));
  XOR2_X1   g0290(.A(KEYINPUT67), .B(G41), .Z(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(G274), .A3(new_n293), .A4(new_n481), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n484), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G200), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G190), .B2(new_n495), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n472), .A2(new_n479), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n367), .A2(new_n214), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n477), .B2(new_n214), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n384), .A2(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT6), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n503), .A2(new_n214), .A3(G107), .ZN(new_n504));
  XNOR2_X1  g0304(.A(G97), .B(G107), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n258), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n506), .A2(new_n222), .B1(new_n284), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(KEYINPUT78), .A3(new_n249), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT78), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n384), .B2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n265), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n501), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(new_n282), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT79), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n286), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n482), .A2(G257), .A3(new_n293), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(G190), .A3(new_n494), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  INV_X1    g0330(.A(new_n526), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n482), .A2(new_n267), .A3(new_n338), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n494), .A2(KEYINPUT80), .A3(new_n526), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n515), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n501), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT78), .B1(new_n510), .B2(new_n249), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n513), .A2(new_n512), .A3(new_n265), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n533), .A2(new_n308), .A3(new_n525), .A4(new_n534), .ZN(new_n542));
  INV_X1    g0342(.A(new_n525), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n494), .A2(new_n526), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n329), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n273), .A2(new_n275), .A3(G238), .A4(new_n282), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  INV_X1    g0349(.A(G244), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n276), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n286), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n480), .A2(G274), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n293), .A2(G250), .A3(new_n490), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n254), .A2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  NAND3_X1  g0358(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n222), .ZN(new_n560));
  INV_X1    g0360(.A(G87), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n214), .A3(new_n464), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n557), .A2(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n279), .A2(new_n222), .A3(G68), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n265), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n433), .A2(new_n252), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n477), .A2(new_n561), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n552), .A2(G190), .A3(new_n553), .A4(new_n554), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n556), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n555), .A2(new_n329), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n563), .A2(new_n564), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n566), .B1(new_n572), .B2(new_n249), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT82), .B1(new_n477), .B2(new_n434), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n367), .A2(new_n249), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n433), .A4(new_n476), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n552), .A2(new_n308), .A3(new_n553), .A4(new_n554), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n571), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n570), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n499), .A2(new_n537), .A3(new_n547), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n495), .A2(G179), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n329), .B2(new_n495), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n469), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT24), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n463), .A2(new_n452), .A3(new_n469), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n265), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n585), .B1(new_n591), .B2(new_n478), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n483), .A2(G270), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n377), .A2(G303), .ZN(new_n594));
  INV_X1    g0394(.A(G264), .ZN(new_n595));
  OAI221_X1 g0395(.A(new_n594), .B1(new_n276), .B2(new_n595), .C1(new_n345), .C2(new_n215), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n286), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n597), .A3(new_n494), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n252), .A2(G116), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n575), .A2(G116), .A3(new_n476), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n265), .B1(G20), .B2(new_n208), .ZN(new_n602));
  AOI21_X1  g0402(.A(G20), .B1(new_n253), .B2(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n523), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n602), .A2(new_n604), .A3(KEYINPUT20), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n602), .B2(new_n604), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n600), .B(new_n601), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n598), .A2(new_n607), .A3(G169), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n598), .A2(new_n308), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n607), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n598), .A2(new_n607), .A3(KEYINPUT21), .A4(G169), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n607), .B1(new_n598), .B2(G200), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n411), .B2(new_n598), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n592), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n451), .A2(new_n583), .A3(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n407), .A2(new_n408), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n429), .A2(new_n439), .ZN(new_n621));
  AOI21_X1  g0421(.A(G169), .B1(new_n443), .B2(new_n426), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT85), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n428), .A2(new_n624), .A3(new_n429), .A4(new_n439), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n373), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n417), .A2(new_n419), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n450), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n620), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n326), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n312), .B(new_n327), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n451), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n537), .A2(new_n547), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n592), .A2(new_n614), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n570), .A2(new_n581), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n589), .A2(new_n590), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n478), .B1(new_n639), .B2(new_n249), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n640), .B2(new_n498), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n581), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n541), .A2(new_n582), .A3(new_n546), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n542), .A2(new_n545), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n511), .A2(new_n514), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n538), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(KEYINPUT26), .A3(new_n582), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n635), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n634), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G13), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G20), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n225), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n499), .B1(new_n640), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n592), .ZN(new_n665));
  INV_X1    g0465(.A(new_n592), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n663), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n607), .A2(new_n662), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n614), .B(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n616), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n672), .A3(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n665), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n614), .A2(new_n662), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n668), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n226), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n491), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n562), .A2(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n221), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n652), .A2(new_n663), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n662), .B1(new_n642), .B2(new_n651), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n583), .A2(new_n617), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT86), .B1(new_n691), .B2(new_n663), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT86), .ZN(new_n693));
  NOR4_X1   g0493(.A1(new_n583), .A2(new_n617), .A3(new_n693), .A4(new_n662), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n543), .A2(new_n555), .A3(new_n544), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n611), .A2(new_n695), .A3(new_n489), .A4(new_n484), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n598), .A2(new_n308), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n555), .A3(new_n495), .A4(new_n535), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n662), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n692), .A2(new_n694), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n690), .B1(G330), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n684), .B1(new_n707), .B2(G1), .ZN(G364));
  AOI21_X1  g0508(.A(new_n225), .B1(new_n656), .B2(G45), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n679), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n243), .A2(G45), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n678), .A2(new_n279), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n712), .B(new_n713), .C1(G45), .C2(new_n221), .ZN(new_n714));
  NAND3_X1  g0514(.A1(G355), .A2(new_n226), .A3(new_n279), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n714), .B(new_n715), .C1(G116), .C2(new_n226), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n223), .B1(G20), .B2(new_n329), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT88), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n222), .A2(new_n308), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n724), .A2(new_n411), .A3(G200), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  INV_X1    g0527(.A(G311), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(new_n411), .A3(new_n496), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n726), .A2(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n724), .A2(new_n496), .A3(G190), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT33), .B(G317), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n730), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(G20), .A2(G190), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n308), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G326), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G303), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n411), .A2(G179), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n222), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n222), .A2(G190), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n308), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(G283), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n743), .A2(new_n487), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n308), .A3(new_n496), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n279), .B(new_n747), .C1(G329), .C2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n736), .A2(new_n739), .A3(new_n741), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n738), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n279), .B1(new_n752), .B2(new_n240), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(G58), .B2(new_n725), .ZN(new_n754));
  INV_X1    g0554(.A(new_n740), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n754), .B1(new_n561), .B2(new_n755), .C1(new_n758), .C2(new_n214), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n734), .A2(G68), .ZN(new_n760));
  INV_X1    g0560(.A(new_n745), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  INV_X1    g0562(.A(G159), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT32), .B1(new_n748), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n748), .A2(KEYINPUT32), .A3(new_n763), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n729), .B(KEYINPUT89), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(G77), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n760), .A2(new_n762), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n751), .B1(new_n759), .B2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n716), .A2(new_n722), .B1(new_n769), .B2(new_n720), .ZN(new_n770));
  INV_X1    g0570(.A(new_n719), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n711), .B(new_n770), .C1(new_n672), .C2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT92), .Z(new_n773));
  AOI21_X1  g0573(.A(new_n711), .B1(new_n672), .B2(G330), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G330), .B2(new_n672), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT93), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n706), .A2(G330), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n439), .A2(new_n662), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n626), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT96), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n445), .A2(new_n440), .A3(new_n781), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n781), .B1(new_n623), .B2(new_n625), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n445), .A2(new_n440), .A3(new_n781), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT96), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n687), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n780), .B(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n711), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n766), .A2(G159), .B1(G137), .B2(new_n738), .ZN(new_n795));
  INV_X1    g0595(.A(G143), .ZN(new_n796));
  INV_X1    g0596(.A(new_n734), .ZN(new_n797));
  INV_X1    g0597(.A(G150), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(new_n796), .B2(new_n726), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT34), .Z(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n748), .A2(new_n801), .B1(new_n745), .B2(new_n212), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n279), .B1(new_n743), .B2(new_n242), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(G50), .C2(new_n740), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT95), .Z(new_n805));
  OAI21_X1  g0605(.A(new_n377), .B1(new_n755), .B2(new_n464), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n806), .A2(KEYINPUT94), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(KEYINPUT94), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n734), .C2(G283), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n766), .A2(G116), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(new_n561), .C2(new_n745), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n725), .A2(G294), .B1(G311), .B2(new_n749), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n813), .B2(new_n752), .C1(new_n758), .C2(new_n214), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n800), .A2(new_n805), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n720), .A2(new_n717), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(new_n720), .B1(new_n284), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n786), .A2(new_n789), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n817), .B(new_n711), .C1(new_n818), .C2(new_n718), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n794), .A2(new_n819), .ZN(G384));
  AND2_X1   g0620(.A1(new_n706), .A2(new_n818), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n372), .A2(new_n662), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT97), .ZN(new_n823));
  INV_X1    g0623(.A(new_n450), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n362), .C2(new_n372), .ZN(new_n825));
  INV_X1    g0625(.A(new_n823), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n373), .B2(new_n450), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT98), .ZN(new_n829));
  INV_X1    g0629(.A(new_n660), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n395), .B1(new_n404), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(new_n416), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n410), .A2(new_n376), .A3(new_n415), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n402), .A2(new_n403), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT16), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n212), .B1(new_n381), .B2(new_n378), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n389), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n393), .A2(new_n838), .A3(new_n249), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n835), .A2(new_n660), .B1(new_n376), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n376), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n830), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(KEYINPUT38), .C1(new_n420), .C2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n416), .A2(KEYINPUT17), .ZN(new_n846));
  INV_X1    g0646(.A(new_n419), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n395), .A2(KEYINPUT18), .A3(new_n404), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT18), .B1(new_n395), .B2(new_n404), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n846), .A2(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n660), .B1(new_n410), .B2(new_n376), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n410), .A2(new_n376), .B1(new_n835), .B2(new_n660), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n852), .B2(new_n834), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n850), .A2(new_n851), .B1(new_n833), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n829), .B(new_n845), .C1(new_n854), .C2(KEYINPUT38), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n844), .B1(new_n619), .B2(new_n629), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n833), .A2(new_n841), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(KEYINPUT98), .A3(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n821), .A2(new_n828), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n856), .B2(new_n857), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n845), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n706), .A2(new_n828), .A3(new_n818), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n861), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n706), .A2(new_n635), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n869), .B(new_n870), .Z(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(G330), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n440), .A2(new_n662), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n472), .A2(new_n479), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n585), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n583), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT26), .B1(new_n649), .B2(new_n582), .ZN(new_n879));
  NOR4_X1   g0679(.A1(new_n515), .A2(new_n638), .A3(new_n647), .A4(new_n645), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n581), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n663), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n874), .B1(new_n882), .B2(new_n790), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n828), .A2(new_n883), .A3(new_n866), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n865), .B2(new_n845), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n860), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n373), .A2(new_n662), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n884), .B1(new_n619), .B2(new_n830), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n872), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n687), .A2(new_n689), .ZN(new_n892));
  INV_X1    g0692(.A(new_n685), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n662), .B(new_n893), .C1(new_n642), .C2(new_n651), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n635), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT99), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT99), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n690), .A2(new_n897), .A3(new_n635), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n633), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n891), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n225), .B2(new_n656), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT35), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n222), .B(new_n223), .C1(new_n506), .C2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(G116), .C1(new_n902), .C2(new_n506), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n221), .A2(new_n284), .A3(new_n386), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n201), .A2(new_n212), .ZN(new_n907));
  OAI211_X1 g0707(.A(G1), .B(new_n655), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(G367));
  NOR2_X1   g0709(.A1(new_n758), .A2(new_n212), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n279), .B1(new_n752), .B2(new_n796), .C1(new_n242), .C2(new_n755), .ZN(new_n911));
  INV_X1    g0711(.A(G137), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n748), .A2(new_n912), .B1(new_n745), .B2(new_n284), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n734), .A2(G159), .B1(new_n201), .B2(new_n766), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT103), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n910), .B(new_n914), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n917), .B1(new_n916), .B2(new_n915), .C1(new_n798), .C2(new_n726), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n726), .A2(new_n813), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n745), .A2(new_n214), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n464), .B2(new_n743), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n279), .B(new_n922), .C1(G311), .C2(new_n738), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n740), .A2(G116), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT46), .Z(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(G317), .B2(new_n749), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n734), .A2(G294), .B1(G283), .B2(new_n766), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n918), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT47), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n793), .B1(new_n930), .B2(new_n720), .ZN(new_n931));
  INV_X1    g0731(.A(new_n713), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n721), .B1(new_n226), .B2(new_n434), .C1(new_n237), .C2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n663), .A2(new_n568), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n582), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n581), .B2(new_n934), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n931), .B(new_n933), .C1(new_n771), .C2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n537), .B(new_n547), .C1(new_n515), .C2(new_n663), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT100), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n649), .A2(new_n662), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT42), .ZN(new_n942));
  INV_X1    g0742(.A(new_n675), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n665), .A2(new_n668), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT101), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n941), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n669), .A2(new_n675), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT42), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n941), .A2(KEYINPUT101), .A3(new_n942), .A4(new_n944), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n547), .B1(new_n939), .B2(new_n592), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n663), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n956), .B1(new_n954), .B2(new_n957), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n948), .A2(new_n673), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n679), .B(KEYINPUT41), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n672), .A2(G330), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n943), .B1(new_n665), .B2(new_n668), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n949), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n949), .B2(new_n966), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n707), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n941), .B2(new_n676), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n941), .A2(new_n676), .A3(new_n972), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n941), .A2(KEYINPUT45), .A3(new_n676), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT45), .B1(new_n941), .B2(new_n676), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n974), .A2(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n673), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  INV_X1    g0781(.A(new_n975), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n973), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n983), .A3(new_n673), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n971), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n964), .B1(new_n985), .B2(new_n707), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n962), .B1(new_n986), .B2(new_n710), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n961), .B1(new_n958), .B2(new_n959), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT102), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(KEYINPUT102), .B(new_n961), .C1(new_n958), .C2(new_n959), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n937), .B1(new_n987), .B2(new_n992), .ZN(G387));
  AOI22_X1  g0793(.A1(new_n766), .A2(G303), .B1(G322), .B2(new_n738), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n797), .B2(new_n728), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G317), .B2(new_n725), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT48), .Z(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n746), .B2(new_n743), .C1(new_n487), .C2(new_n755), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT49), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n749), .A2(G326), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n999), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n279), .B1(new_n761), .B2(G116), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n279), .B1(new_n212), .B2(new_n729), .C1(new_n726), .C2(new_n240), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n431), .B2(new_n734), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n740), .A2(G77), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n738), .A2(KEYINPUT106), .A3(G159), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n921), .B(new_n1008), .C1(new_n798), .C2(new_n748), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT106), .B1(new_n738), .B2(G159), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n758), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n433), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1006), .A2(new_n1007), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1004), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n793), .B1(new_n1015), .B2(new_n720), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n722), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n431), .A2(new_n240), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n681), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n1018), .B2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(G68), .A2(G77), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n269), .A4(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n713), .B(new_n1023), .C1(new_n234), .C2(new_n269), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1020), .A2(new_n226), .A3(new_n279), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G107), .C2(new_n226), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT105), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1016), .B1(new_n669), .B2(new_n771), .C1(new_n1017), .C2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n969), .A2(new_n707), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n679), .A3(new_n970), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n710), .B1(new_n967), .B2(new_n968), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT104), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(G393));
  NAND3_X1  g0833(.A1(new_n980), .A2(new_n984), .A3(new_n710), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n720), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n377), .B1(new_n729), .B2(new_n487), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n762), .B1(new_n727), .B2(new_n748), .C1(new_n208), .C2(new_n743), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G303), .C2(new_n734), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n725), .A2(G311), .B1(new_n738), .B2(G317), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT52), .Z(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n746), .C2(new_n755), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT110), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n734), .A2(new_n201), .B1(new_n431), .B2(new_n766), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n725), .A2(G159), .B1(new_n738), .B2(G150), .ZN(new_n1044));
  XOR2_X1   g0844(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1012), .A2(G77), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n279), .B1(new_n748), .B2(new_n796), .C1(new_n212), .C2(new_n755), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G87), .B2(new_n761), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1035), .B1(new_n1042), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n948), .A2(new_n719), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n793), .B(new_n1051), .C1(new_n1052), .C2(KEYINPUT107), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n721), .B1(new_n214), .B2(new_n226), .C1(new_n246), .C2(new_n932), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT108), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(KEYINPUT107), .C2(new_n1052), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n971), .B1(new_n980), .B2(new_n984), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n679), .B1(new_n1057), .B2(KEYINPUT111), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n978), .A2(new_n979), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n673), .B1(new_n981), .B2(new_n983), .ZN(new_n1060));
  OAI211_X1 g0860(.A(KEYINPUT111), .B(new_n970), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n985), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1034), .B(new_n1056), .C1(new_n1058), .C2(new_n1062), .ZN(G390));
  AOI21_X1  g0863(.A(new_n360), .B1(new_n359), .B2(new_n330), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n330), .ZN(new_n1065));
  AOI211_X1 g0865(.A(KEYINPUT14), .B(new_n1065), .C1(new_n356), .C2(new_n357), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n448), .B1(new_n1067), .B2(new_n358), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n823), .B1(new_n1068), .B2(new_n824), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n373), .A2(new_n450), .A3(new_n826), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n873), .B1(new_n687), .B2(new_n818), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n860), .B(new_n889), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n888), .B1(new_n828), .B2(new_n883), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n887), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT112), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT112), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(new_n1074), .C2(new_n887), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n828), .A2(new_n706), .A3(new_n818), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(G330), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1075), .A2(new_n1079), .A3(KEYINPUT112), .A4(G330), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n828), .A2(new_n883), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n706), .A2(G330), .A3(new_n818), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n706), .A2(G330), .A3(new_n635), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n821), .A2(new_n1085), .A3(G330), .A4(new_n1084), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n899), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1081), .A2(new_n1091), .A3(new_n1082), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n679), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n887), .A2(new_n717), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT53), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n755), .B2(new_n798), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n740), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n734), .A2(G137), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n766), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1012), .A2(G159), .ZN(new_n1103));
  INV_X1    g0903(.A(G125), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n261), .A2(new_n745), .B1(new_n748), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n377), .B(new_n1105), .C1(G128), .C2(new_n738), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n726), .A2(new_n801), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n377), .B1(new_n752), .B2(new_n746), .C1(new_n561), .C2(new_n755), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n734), .B2(G107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n725), .A2(G116), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n766), .A2(G97), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1110), .A2(new_n1047), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n748), .A2(new_n487), .B1(new_n745), .B2(new_n212), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT113), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1107), .A2(new_n1108), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n720), .B1(new_n374), .B2(new_n816), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n711), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1083), .B2(new_n710), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1095), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G378));
  NAND2_X1  g0924(.A1(new_n326), .A2(new_n310), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n305), .A2(new_n660), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT55), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1129), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT55), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n1127), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT56), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1130), .A2(new_n1133), .A3(KEYINPUT56), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n869), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1138), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n863), .A3(new_n868), .A4(G330), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1140), .A2(new_n890), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n890), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n710), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1101), .A2(new_n740), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT116), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n726), .A2(new_n1149), .B1(new_n912), .B2(new_n729), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(new_n734), .C2(G132), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n1104), .B2(new_n752), .C1(new_n798), .C2(new_n758), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n749), .A2(G124), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G33), .B(G41), .C1(new_n761), .C2(G159), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n910), .B1(G116), .B2(new_n738), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT115), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n748), .A2(new_n746), .B1(new_n745), .B2(new_n242), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n491), .A2(new_n279), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n1007), .C1(new_n434), .C2(new_n729), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(new_n734), .C2(G97), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1159), .B(new_n1163), .C1(new_n464), .C2(new_n726), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT58), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1157), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n240), .B1(G33), .B2(G41), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1167), .B1(new_n1165), .B2(new_n1164), .C1(new_n1161), .C2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(new_n720), .B1(new_n261), .B2(new_n816), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n711), .B(new_n1170), .C1(new_n1138), .C2(new_n718), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1146), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT118), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n690), .A2(new_n897), .A3(new_n635), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n897), .B1(new_n690), .B2(new_n635), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n634), .B(new_n1089), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT117), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1093), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1091), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT117), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1177), .B(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT118), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1173), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT120), .B1(new_n1184), .B2(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1174), .B1(new_n1093), .B2(new_n1178), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1180), .A2(new_n1182), .A3(KEYINPUT118), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1145), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(KEYINPUT119), .B(new_n890), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1173), .B2(KEYINPUT119), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n679), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1172), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT121), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1185), .A2(new_n1191), .A3(new_n679), .A4(new_n1196), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT121), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n1172), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(G375));
  NAND2_X1  g1003(.A1(new_n1090), .A2(new_n1088), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1177), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n1091), .A3(new_n963), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1013), .B1(new_n746), .B2(new_n726), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  AOI21_X1  g1008(.A(new_n279), .B1(new_n740), .B2(G97), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n284), .B2(new_n745), .C1(new_n813), .C2(new_n748), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n797), .A2(new_n208), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G107), .C2(new_n766), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1208), .B(new_n1212), .C1(new_n487), .C2(new_n752), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n748), .A2(new_n1149), .B1(new_n745), .B2(new_n242), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n279), .B1(new_n729), .B2(new_n798), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n726), .A2(new_n912), .B1(new_n755), .B2(new_n763), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n734), .C2(new_n1101), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n240), .B2(new_n758), .C1(new_n801), .C2(new_n752), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1213), .A2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT123), .Z(new_n1221));
  OAI221_X1 g1021(.A(new_n711), .B1(new_n828), .B2(new_n718), .C1(new_n1035), .C2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n212), .B2(new_n816), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1204), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n710), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1225), .ZN(G381));
  AND3_X1   g1026(.A1(new_n1200), .A2(new_n1201), .A3(new_n1172), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1201), .B1(new_n1200), .B2(new_n1172), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1227), .A2(new_n1228), .A3(G378), .ZN(new_n1229));
  INV_X1    g1029(.A(G384), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1225), .A4(new_n1206), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n985), .A2(new_n707), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n709), .B1(new_n1232), .B2(new_n964), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1233), .A2(new_n962), .A3(new_n990), .A4(new_n991), .ZN(new_n1234));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n937), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n778), .A2(new_n1030), .A3(new_n1028), .A4(new_n1032), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1231), .A2(new_n1238), .ZN(G407));
  NAND3_X1  g1039(.A1(new_n1199), .A2(new_n1123), .A3(new_n1202), .ZN(new_n1240));
  OAI221_X1 g1040(.A(G213), .B1(G343), .B2(new_n1240), .C1(new_n1231), .C2(new_n1238), .ZN(G409));
  AND2_X1   g1041(.A1(G387), .A2(G390), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G396), .A2(G393), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n1237), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1245), .A2(new_n1244), .A3(new_n1237), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1242), .A2(new_n1243), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G387), .A2(G390), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1247), .A2(new_n1246), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1236), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1123), .B1(new_n1200), .B2(new_n1172), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1184), .A2(new_n963), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1194), .A2(new_n710), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1123), .A4(new_n1171), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n661), .A2(G213), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n680), .B1(new_n1205), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1091), .C1(new_n1260), .C2(new_n1205), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1225), .ZN(new_n1263));
  OR3_X1    g1063(.A1(new_n1263), .A2(KEYINPUT124), .A3(new_n1230), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1230), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT124), .B1(new_n1263), .B2(new_n1230), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n661), .A2(G213), .A3(G2897), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1267), .B(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1270), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1271), .A2(new_n1267), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1252), .B(new_n1269), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1273), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1259), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1259), .B2(new_n1268), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(new_n1253), .A2(KEYINPUT62), .A3(new_n1258), .A4(new_n1267), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1236), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1250), .B1(new_n1236), .B2(new_n1249), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1248), .A2(KEYINPUT126), .A3(new_n1251), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1276), .B1(new_n1283), .B2(new_n1289), .ZN(G405));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1253), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1240), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1240), .B2(new_n1292), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1267), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1289), .B1(new_n1229), .B2(new_n1253), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1240), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1268), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1295), .A2(new_n1298), .ZN(G402));
endmodule


