

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833;

  XNOR2_X1 U375 ( .A(n466), .B(n647), .ZN(n353) );
  XNOR2_X1 U376 ( .A(n629), .B(n393), .ZN(n680) );
  AND2_X1 U377 ( .A1(n504), .A2(n495), .ZN(n365) );
  XNOR2_X1 U378 ( .A(n396), .B(n806), .ZN(n480) );
  XNOR2_X1 U379 ( .A(G113), .B(G143), .ZN(n569) );
  BUF_X1 U380 ( .A(G107), .Z(n364) );
  XNOR2_X1 U381 ( .A(n552), .B(n394), .ZN(n608) );
  XNOR2_X1 U382 ( .A(n804), .B(KEYINPUT74), .ZN(n402) );
  XNOR2_X1 U383 ( .A(n574), .B(n573), .ZN(n610) );
  NAND2_X1 U384 ( .A1(n467), .A2(n353), .ZN(n671) );
  XNOR2_X2 U385 ( .A(n674), .B(KEYINPUT40), .ZN(n831) );
  NAND2_X1 U386 ( .A1(n550), .A2(n549), .ZN(n524) );
  NAND2_X1 U387 ( .A1(n547), .A2(G143), .ZN(n550) );
  NOR2_X2 U388 ( .A1(n671), .A2(n693), .ZN(n651) );
  XNOR2_X2 U389 ( .A(n651), .B(KEYINPUT110), .ZN(n471) );
  NAND2_X1 U390 ( .A1(n354), .A2(n522), .ZN(n523) );
  NAND2_X1 U391 ( .A1(n711), .A2(n712), .ZN(n354) );
  XNOR2_X2 U392 ( .A(n355), .B(KEYINPUT35), .ZN(n829) );
  NAND2_X1 U393 ( .A1(n430), .A2(n428), .ZN(n355) );
  XNOR2_X1 U394 ( .A(n608), .B(n553), .ZN(n806) );
  XNOR2_X2 U395 ( .A(n535), .B(n494), .ZN(n375) );
  NOR2_X2 U396 ( .A1(n730), .A2(n663), .ZN(n664) );
  XNOR2_X1 U397 ( .A(n427), .B(n526), .ZN(n702) );
  OR2_X2 U398 ( .A1(n567), .A2(n510), .ZN(n509) );
  NOR2_X1 U399 ( .A1(n828), .A2(n724), .ZN(n642) );
  XNOR2_X2 U400 ( .A(n660), .B(KEYINPUT1), .ZN(n747) );
  INV_X2 U401 ( .A(G113), .ZN(n395) );
  NOR2_X1 U402 ( .A1(n628), .A2(n629), .ZN(n721) );
  XNOR2_X1 U403 ( .A(n627), .B(KEYINPUT31), .ZN(n735) );
  NOR2_X1 U404 ( .A1(n735), .A2(n721), .ZN(n357) );
  NOR2_X1 U405 ( .A1(n638), .A2(n680), .ZN(n419) );
  AND2_X1 U406 ( .A1(n629), .A2(n624), .ZN(n625) );
  XNOR2_X1 U407 ( .A(n619), .B(n618), .ZN(n742) );
  XNOR2_X1 U408 ( .A(KEYINPUT71), .B(G131), .ZN(n379) );
  XNOR2_X1 U409 ( .A(n361), .B(n793), .ZN(n794) );
  NAND2_X1 U410 ( .A1(n413), .A2(n409), .ZN(n828) );
  AND2_X1 U411 ( .A1(n356), .A2(n653), .ZN(n387) );
  XNOR2_X1 U412 ( .A(n357), .B(KEYINPUT99), .ZN(n356) );
  NAND2_X1 U413 ( .A1(n412), .A2(n410), .ZN(n409) );
  AND2_X1 U414 ( .A1(n416), .A2(n414), .ZN(n413) );
  NAND2_X1 U415 ( .A1(n429), .A2(n433), .ZN(n428) );
  XNOR2_X1 U416 ( .A(n675), .B(n479), .ZN(n754) );
  AND2_X1 U417 ( .A1(n457), .A2(n476), .ZN(n676) );
  NOR2_X1 U418 ( .A1(n759), .A2(n762), .ZN(n675) );
  XNOR2_X1 U419 ( .A(n625), .B(KEYINPUT98), .ZN(n751) );
  OR2_X1 U420 ( .A1(n763), .A2(KEYINPUT47), .ZN(n663) );
  AND2_X1 U421 ( .A1(n541), .A2(n519), .ZN(n483) );
  AND2_X1 U422 ( .A1(n503), .A2(n502), .ZN(n501) );
  NAND2_X1 U423 ( .A1(n602), .A2(n601), .ZN(n427) );
  AND2_X1 U424 ( .A1(n506), .A2(n560), .ZN(n495) );
  XNOR2_X1 U425 ( .A(n610), .B(n423), .ZN(n817) );
  XNOR2_X1 U426 ( .A(n546), .B(n545), .ZN(n598) );
  INV_X1 U427 ( .A(n379), .ZN(n576) );
  XNOR2_X1 U428 ( .A(KEYINPUT97), .B(KEYINPUT24), .ZN(n366) );
  XOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n555) );
  XNOR2_X1 U430 ( .A(G119), .B(KEYINPUT3), .ZN(n552) );
  XNOR2_X1 U431 ( .A(G140), .B(KEYINPUT10), .ZN(n573) );
  XOR2_X1 U432 ( .A(G137), .B(KEYINPUT72), .Z(n611) );
  NAND2_X1 U433 ( .A1(n359), .A2(G210), .ZN(n711) );
  NAND2_X1 U434 ( .A1(n359), .A2(n358), .ZN(n522) );
  AND2_X1 U435 ( .A1(n710), .A2(G210), .ZN(n358) );
  XNOR2_X1 U436 ( .A(n449), .B(KEYINPUT65), .ZN(n359) );
  XNOR2_X1 U437 ( .A(n360), .B(G128), .ZN(n615) );
  XNOR2_X2 U438 ( .A(G110), .B(KEYINPUT23), .ZN(n360) );
  INV_X1 U439 ( .A(n366), .ZN(n613) );
  NAND2_X1 U440 ( .A1(n792), .A2(G475), .ZN(n361) );
  XNOR2_X2 U441 ( .A(n372), .B(KEYINPUT65), .ZN(n792) );
  NAND2_X1 U442 ( .A1(n474), .A2(n701), .ZN(n362) );
  NAND2_X1 U443 ( .A1(n474), .A2(n701), .ZN(n473) );
  BUF_X1 U444 ( .A(n702), .Z(n363) );
  XNOR2_X2 U445 ( .A(n640), .B(n491), .ZN(n659) );
  NAND2_X2 U446 ( .A1(n509), .A2(n508), .ZN(n626) );
  NAND2_X1 U447 ( .A1(n613), .A2(n612), .ZN(n368) );
  NAND2_X1 U448 ( .A1(n366), .A2(n367), .ZN(n369) );
  NAND2_X1 U449 ( .A1(n369), .A2(n368), .ZN(n614) );
  INV_X1 U450 ( .A(n612), .ZN(n367) );
  XNOR2_X1 U451 ( .A(n576), .B(n478), .ZN(n407) );
  NOR2_X1 U452 ( .A1(n387), .A2(n450), .ZN(n636) );
  BUF_X1 U453 ( .A(n735), .Z(n370) );
  NAND2_X1 U454 ( .A1(n549), .A2(n550), .ZN(n371) );
  NOR2_X1 U455 ( .A1(n747), .A2(n746), .ZN(n624) );
  NAND2_X1 U456 ( .A1(n362), .A2(n472), .ZN(n372) );
  NAND2_X1 U457 ( .A1(n362), .A2(n472), .ZN(n373) );
  BUF_X1 U458 ( .A(n801), .Z(n374) );
  NAND2_X1 U459 ( .A1(n473), .A2(n472), .ZN(n449) );
  NOR2_X2 U460 ( .A1(n801), .A2(G902), .ZN(n619) );
  NOR2_X2 U461 ( .A1(n785), .A2(G902), .ZN(n442) );
  XNOR2_X1 U462 ( .A(n371), .B(G134), .ZN(n376) );
  XNOR2_X1 U463 ( .A(n524), .B(G134), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n373), .B(KEYINPUT65), .ZN(n377) );
  BUF_X1 U465 ( .A(n437), .Z(n378) );
  AND2_X1 U466 ( .A1(n439), .A2(n469), .ZN(n438) );
  NAND2_X1 U467 ( .A1(n751), .A2(n626), .ZN(n627) );
  NAND2_X1 U468 ( .A1(n505), .A2(n504), .ZN(n669) );
  BUF_X1 U469 ( .A(n730), .Z(n380) );
  XNOR2_X1 U470 ( .A(n662), .B(KEYINPUT84), .ZN(n730) );
  INV_X1 U471 ( .A(n378), .ZN(n381) );
  BUF_X1 U472 ( .A(n659), .Z(n382) );
  NOR2_X1 U473 ( .A1(n383), .A2(n384), .ZN(n469) );
  AND2_X1 U474 ( .A1(KEYINPUT47), .A2(n763), .ZN(n383) );
  XNOR2_X1 U475 ( .A(G101), .B(KEYINPUT4), .ZN(n544) );
  XNOR2_X1 U476 ( .A(n669), .B(n399), .ZN(n757) );
  INV_X1 U477 ( .A(KEYINPUT38), .ZN(n399) );
  INV_X1 U478 ( .A(KEYINPUT106), .ZN(n491) );
  XNOR2_X1 U479 ( .A(n617), .B(KEYINPUT25), .ZN(n618) );
  AND2_X2 U480 ( .A1(n432), .A2(n652), .ZN(n431) );
  OR2_X2 U481 ( .A1(n626), .A2(n527), .ZN(n432) );
  OR2_X1 U482 ( .A1(G237), .A2(G902), .ZN(n557) );
  NOR2_X1 U483 ( .A1(n650), .A2(n452), .ZN(n655) );
  XNOR2_X1 U484 ( .A(n454), .B(n453), .ZN(n452) );
  INV_X1 U485 ( .A(KEYINPUT107), .ZN(n453) );
  NOR2_X1 U486 ( .A1(n648), .A2(n455), .ZN(n454) );
  NAND2_X1 U487 ( .A1(n500), .A2(n391), .ZN(n499) );
  INV_X1 U488 ( .A(G146), .ZN(n478) );
  INV_X1 U489 ( .A(KEYINPUT5), .ZN(n605) );
  XNOR2_X1 U490 ( .A(G137), .B(KEYINPUT79), .ZN(n606) );
  XNOR2_X1 U491 ( .A(n611), .B(n406), .ZN(n405) );
  XNOR2_X1 U492 ( .A(KEYINPUT96), .B(G140), .ZN(n406) );
  NAND2_X1 U493 ( .A1(n757), .A2(n756), .ZN(n762) );
  XNOR2_X1 U494 ( .A(KEYINPUT34), .B(KEYINPUT83), .ZN(n527) );
  AND2_X1 U495 ( .A1(n475), .A2(n464), .ZN(n463) );
  INV_X1 U496 ( .A(KEYINPUT8), .ZN(n585) );
  INV_X1 U497 ( .A(n611), .ZN(n423) );
  XOR2_X1 U498 ( .A(KEYINPUT7), .B(G122), .Z(n583) );
  XNOR2_X1 U499 ( .A(G116), .B(n364), .ZN(n582) );
  XOR2_X1 U500 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n588) );
  INV_X1 U501 ( .A(KEYINPUT80), .ZN(n520) );
  XOR2_X1 U502 ( .A(KEYINPUT11), .B(G122), .Z(n570) );
  NAND2_X1 U503 ( .A1(n624), .A2(n680), .ZN(n622) );
  INV_X1 U504 ( .A(KEYINPUT39), .ZN(n672) );
  NAND2_X1 U505 ( .A1(n768), .A2(n435), .ZN(n434) );
  AND2_X1 U506 ( .A1(n626), .A2(n527), .ZN(n435) );
  INV_X1 U507 ( .A(n527), .ZN(n433) );
  XNOR2_X1 U508 ( .A(n580), .B(n487), .ZN(n630) );
  XNOR2_X1 U509 ( .A(n581), .B(n488), .ZN(n487) );
  INV_X1 U510 ( .A(G475), .ZN(n488) );
  XNOR2_X1 U511 ( .A(n459), .B(n458), .ZN(n457) );
  INV_X1 U512 ( .A(KEYINPUT28), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n421), .B(G478), .ZN(n634) );
  OR2_X1 U514 ( .A1(n797), .A2(G902), .ZN(n421) );
  XNOR2_X1 U515 ( .A(n595), .B(KEYINPUT22), .ZN(n596) );
  NOR2_X1 U516 ( .A1(n481), .A2(G952), .ZN(n803) );
  NAND2_X1 U517 ( .A1(n437), .A2(n468), .ZN(n436) );
  INV_X1 U518 ( .A(KEYINPUT86), .ZN(n468) );
  INV_X1 U519 ( .A(KEYINPUT85), .ZN(n489) );
  INV_X1 U520 ( .A(KEYINPUT93), .ZN(n558) );
  NAND2_X1 U521 ( .A1(n746), .A2(KEYINPUT108), .ZN(n541) );
  NAND2_X1 U522 ( .A1(n649), .A2(n456), .ZN(n455) );
  INV_X1 U523 ( .A(G900), .ZN(n456) );
  INV_X1 U524 ( .A(G128), .ZN(n547) );
  INV_X1 U525 ( .A(KEYINPUT44), .ZN(n641) );
  NAND2_X1 U526 ( .A1(n525), .A2(n745), .ZN(n750) );
  NOR2_X1 U527 ( .A1(n746), .A2(KEYINPUT108), .ZN(n539) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n494) );
  XNOR2_X1 U529 ( .A(n461), .B(n460), .ZN(n562) );
  XNOR2_X1 U530 ( .A(KEYINPUT78), .B(KEYINPUT94), .ZN(n460) );
  XNOR2_X1 U531 ( .A(n561), .B(KEYINPUT14), .ZN(n461) );
  NAND2_X1 U532 ( .A1(G234), .A2(G237), .ZN(n561) );
  XNOR2_X1 U533 ( .A(n639), .B(KEYINPUT32), .ZN(n516) );
  NOR2_X1 U534 ( .A1(n658), .A2(n485), .ZN(n681) );
  NAND2_X1 U535 ( .A1(n501), .A2(n497), .ZN(n654) );
  AND2_X1 U536 ( .A1(n499), .A2(n498), .ZN(n497) );
  NAND2_X1 U537 ( .A1(KEYINPUT68), .A2(KEYINPUT0), .ZN(n514) );
  NAND2_X1 U538 ( .A1(n515), .A2(n568), .ZN(n513) );
  AND2_X1 U539 ( .A1(n512), .A2(n511), .ZN(n510) );
  NAND2_X1 U540 ( .A1(n515), .A2(KEYINPUT0), .ZN(n511) );
  NAND2_X1 U541 ( .A1(KEYINPUT68), .A2(n568), .ZN(n512) );
  XNOR2_X1 U542 ( .A(n609), .B(n604), .ZN(n526) );
  XOR2_X1 U543 ( .A(KEYINPUT67), .B(n700), .Z(n701) );
  INV_X1 U544 ( .A(n554), .ZN(n401) );
  XNOR2_X1 U545 ( .A(n600), .B(n404), .ZN(n403) );
  XNOR2_X1 U546 ( .A(n551), .B(n405), .ZN(n404) );
  XNOR2_X1 U547 ( .A(n529), .B(KEYINPUT45), .ZN(n528) );
  INV_X1 U548 ( .A(KEYINPUT88), .ZN(n529) );
  INV_X1 U549 ( .A(KEYINPUT41), .ZN(n479) );
  INV_X1 U550 ( .A(n669), .ZN(n693) );
  INV_X1 U551 ( .A(n486), .ZN(n476) );
  XNOR2_X1 U552 ( .A(G122), .B(KEYINPUT16), .ZN(n553) );
  XNOR2_X1 U553 ( .A(n424), .B(n817), .ZN(n801) );
  XNOR2_X1 U554 ( .A(n589), .B(n422), .ZN(n797) );
  XNOR2_X1 U555 ( .A(n578), .B(n390), .ZN(n791) );
  AND2_X2 U556 ( .A1(n431), .A2(n434), .ZN(n430) );
  NOR2_X1 U557 ( .A1(n691), .A2(n382), .ZN(n418) );
  INV_X1 U558 ( .A(KEYINPUT56), .ZN(n530) );
  INV_X1 U559 ( .A(n803), .ZN(n532) );
  NOR2_X1 U560 ( .A1(n652), .A2(KEYINPUT86), .ZN(n384) );
  INV_X1 U561 ( .A(KEYINPUT68), .ZN(n515) );
  XOR2_X1 U562 ( .A(n559), .B(n558), .Z(n385) );
  OR2_X1 U563 ( .A1(n385), .A2(n697), .ZN(n386) );
  AND2_X1 U564 ( .A1(n514), .A2(n513), .ZN(n388) );
  AND2_X1 U565 ( .A1(n476), .A2(n538), .ZN(n389) );
  XOR2_X1 U566 ( .A(n577), .B(n579), .Z(n390) );
  AND2_X1 U567 ( .A1(n756), .A2(KEYINPUT19), .ZN(n391) );
  NOR2_X1 U568 ( .A1(n696), .A2(n740), .ZN(n392) );
  INV_X1 U569 ( .A(n485), .ZN(n417) );
  BUF_X1 U570 ( .A(n742), .Z(n485) );
  XOR2_X1 U571 ( .A(KEYINPUT104), .B(KEYINPUT6), .Z(n393) );
  INV_X1 U572 ( .A(KEYINPUT81), .ZN(n464) );
  XNOR2_X2 U573 ( .A(n395), .B(G116), .ZN(n394) );
  XNOR2_X2 U574 ( .A(n556), .B(n397), .ZN(n396) );
  XNOR2_X2 U575 ( .A(n398), .B(n555), .ZN(n397) );
  NAND2_X1 U576 ( .A1(n584), .A2(G224), .ZN(n398) );
  XNOR2_X1 U577 ( .A(n400), .B(n379), .ZN(n443) );
  XNOR2_X1 U578 ( .A(n590), .B(n376), .ZN(n422) );
  XNOR2_X1 U579 ( .A(n407), .B(n376), .ZN(n600) );
  XNOR2_X2 U580 ( .A(n403), .B(n401), .ZN(n785) );
  XNOR2_X2 U581 ( .A(n402), .B(n598), .ZN(n554) );
  NAND2_X1 U582 ( .A1(n408), .A2(G217), .ZN(n587) );
  NAND2_X1 U583 ( .A1(n408), .A2(G221), .ZN(n517) );
  XNOR2_X2 U584 ( .A(n586), .B(n585), .ZN(n408) );
  AND2_X1 U585 ( .A1(n419), .A2(n411), .ZN(n410) );
  NOR2_X1 U586 ( .A1(n485), .A2(n516), .ZN(n411) );
  INV_X1 U587 ( .A(n637), .ZN(n412) );
  NAND2_X1 U588 ( .A1(n415), .A2(n516), .ZN(n414) );
  NAND2_X1 U589 ( .A1(n419), .A2(n417), .ZN(n415) );
  NAND2_X1 U590 ( .A1(n637), .A2(n516), .ZN(n416) );
  NOR2_X1 U591 ( .A1(n637), .A2(n485), .ZN(n420) );
  AND2_X1 U592 ( .A1(n420), .A2(n418), .ZN(n724) );
  XNOR2_X1 U593 ( .A(n517), .B(n425), .ZN(n424) );
  XNOR2_X1 U594 ( .A(n614), .B(n484), .ZN(n425) );
  XNOR2_X2 U595 ( .A(n426), .B(G472), .ZN(n640) );
  NOR2_X2 U596 ( .A1(n702), .A2(G902), .ZN(n426) );
  INV_X1 U597 ( .A(n768), .ZN(n429) );
  XNOR2_X2 U598 ( .A(n622), .B(KEYINPUT33), .ZN(n768) );
  NAND2_X1 U599 ( .A1(n438), .A2(n436), .ZN(n490) );
  INV_X1 U600 ( .A(n471), .ZN(n437) );
  NAND2_X1 U601 ( .A1(n471), .A2(n470), .ZN(n439) );
  NAND2_X1 U602 ( .A1(n659), .A2(n756), .ZN(n466) );
  BUF_X1 U603 ( .A(n443), .Z(n440) );
  NAND2_X1 U604 ( .A1(n661), .A2(n441), .ZN(n508) );
  NOR2_X1 U605 ( .A1(n566), .A2(n388), .ZN(n441) );
  XNOR2_X2 U606 ( .A(n442), .B(G469), .ZN(n660) );
  AND2_X2 U607 ( .A1(n483), .A2(n542), .ZN(n444) );
  NOR2_X1 U608 ( .A1(n809), .A2(n446), .ZN(n445) );
  NOR2_X1 U609 ( .A1(n809), .A2(n446), .ZN(n778) );
  NAND2_X1 U610 ( .A1(n375), .A2(n392), .ZN(n446) );
  NAND2_X1 U611 ( .A1(n375), .A2(n392), .ZN(n821) );
  NOR2_X1 U612 ( .A1(n668), .A2(n667), .ZN(n537) );
  NAND2_X1 U613 ( .A1(n448), .A2(n447), .ZN(n467) );
  NAND2_X1 U614 ( .A1(n463), .A2(n444), .ZN(n447) );
  NAND2_X1 U615 ( .A1(n462), .A2(KEYINPUT81), .ZN(n448) );
  NAND2_X1 U616 ( .A1(n635), .A2(n451), .ZN(n450) );
  INV_X1 U617 ( .A(n714), .ZN(n451) );
  NAND2_X1 U618 ( .A1(n681), .A2(n659), .ZN(n459) );
  NAND2_X1 U619 ( .A1(n444), .A2(n475), .ZN(n462) );
  NAND2_X1 U620 ( .A1(n381), .A2(n652), .ZN(n728) );
  AND2_X1 U621 ( .A1(n652), .A2(KEYINPUT86), .ZN(n470) );
  XNOR2_X1 U622 ( .A(n443), .B(n478), .ZN(n477) );
  XNOR2_X1 U623 ( .A(n440), .B(KEYINPUT4), .ZN(n818) );
  NAND2_X1 U624 ( .A1(n778), .A2(KEYINPUT2), .ZN(n472) );
  NAND2_X1 U625 ( .A1(n493), .A2(n492), .ZN(n474) );
  NAND2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n475) );
  INV_X1 U627 ( .A(n660), .ZN(n540) );
  NAND2_X1 U628 ( .A1(n477), .A2(n598), .ZN(n602) );
  XNOR2_X1 U629 ( .A(n679), .B(n678), .ZN(n688) );
  NAND2_X1 U630 ( .A1(n754), .A2(n676), .ZN(n677) );
  XNOR2_X2 U631 ( .A(n480), .B(n554), .ZN(n713) );
  INV_X1 U632 ( .A(n615), .ZN(n484) );
  BUF_X2 U633 ( .A(n584), .Z(n481) );
  XNOR2_X2 U634 ( .A(n482), .B(n528), .ZN(n809) );
  NAND2_X1 U635 ( .A1(n646), .A2(n645), .ZN(n482) );
  XNOR2_X1 U636 ( .A(n490), .B(n489), .ZN(n668) );
  BUF_X1 U637 ( .A(n660), .Z(n486) );
  NOR2_X2 U638 ( .A1(n705), .A2(n803), .ZN(n709) );
  NAND2_X1 U639 ( .A1(n729), .A2(n725), .ZN(n653) );
  NAND2_X1 U640 ( .A1(n633), .A2(n634), .ZN(n725) );
  NOR2_X2 U641 ( .A1(n794), .A2(n803), .ZN(n795) );
  XNOR2_X1 U642 ( .A(n821), .B(n520), .ZN(n493) );
  NOR2_X1 U643 ( .A1(n809), .A2(n698), .ZN(n492) );
  NAND2_X1 U644 ( .A1(n365), .A2(n507), .ZN(n503) );
  OR2_X2 U645 ( .A1(n713), .A2(n386), .ZN(n504) );
  INV_X1 U646 ( .A(n496), .ZN(n505) );
  NAND2_X1 U647 ( .A1(n507), .A2(n506), .ZN(n496) );
  NAND2_X1 U648 ( .A1(n496), .A2(n391), .ZN(n502) );
  OR2_X1 U649 ( .A1(n756), .A2(KEYINPUT19), .ZN(n498) );
  INV_X1 U650 ( .A(n504), .ZN(n500) );
  NAND2_X1 U651 ( .A1(n385), .A2(n697), .ZN(n506) );
  NAND2_X1 U652 ( .A1(n713), .A2(n385), .ZN(n507) );
  NAND2_X1 U653 ( .A1(n594), .A2(n626), .ZN(n597) );
  INV_X4 U654 ( .A(KEYINPUT64), .ZN(n518) );
  XNOR2_X2 U655 ( .A(n518), .B(G953), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n584), .A2(G234), .ZN(n586) );
  INV_X1 U657 ( .A(n655), .ZN(n519) );
  XOR2_X2 U658 ( .A(G146), .B(G125), .Z(n574) );
  XNOR2_X1 U659 ( .A(n523), .B(n534), .ZN(n533) );
  XNOR2_X1 U660 ( .A(n371), .B(n574), .ZN(n556) );
  INV_X1 U661 ( .A(n629), .ZN(n525) );
  XNOR2_X1 U662 ( .A(n531), .B(n530), .ZN(G51) );
  NAND2_X1 U663 ( .A1(n533), .A2(n532), .ZN(n531) );
  INV_X1 U664 ( .A(n713), .ZN(n534) );
  NAND2_X1 U665 ( .A1(n536), .A2(n689), .ZN(n535) );
  XNOR2_X1 U666 ( .A(n537), .B(KEYINPUT76), .ZN(n536) );
  NAND2_X2 U667 ( .A1(n742), .A2(n743), .ZN(n746) );
  INV_X1 U668 ( .A(n746), .ZN(n538) );
  NAND2_X1 U669 ( .A1(n660), .A2(KEYINPUT108), .ZN(n542) );
  XNOR2_X2 U670 ( .A(n543), .B(G110), .ZN(n804) );
  XNOR2_X2 U671 ( .A(G104), .B(G107), .ZN(n543) );
  NOR2_X1 U672 ( .A1(n654), .A2(n566), .ZN(n567) );
  XNOR2_X1 U673 ( .A(n606), .B(n605), .ZN(n607) );
  INV_X1 U674 ( .A(KEYINPUT19), .ZN(n560) );
  XNOR2_X1 U675 ( .A(n608), .B(n607), .ZN(n609) );
  INV_X1 U676 ( .A(KEYINPUT66), .ZN(n639) );
  XNOR2_X1 U677 ( .A(n707), .B(n706), .ZN(n708) );
  INV_X1 U678 ( .A(n544), .ZN(n546) );
  XNOR2_X1 U679 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n545) );
  INV_X2 U680 ( .A(G143), .ZN(n548) );
  NAND2_X1 U681 ( .A1(n548), .A2(G128), .ZN(n549) );
  AND2_X1 U682 ( .A1(G227), .A2(n481), .ZN(n551) );
  INV_X1 U683 ( .A(n747), .ZN(n691) );
  NAND2_X1 U684 ( .A1(G214), .A2(n557), .ZN(n756) );
  XOR2_X1 U685 ( .A(G902), .B(KEYINPUT15), .Z(n697) );
  NAND2_X1 U686 ( .A1(G210), .A2(n557), .ZN(n559) );
  NAND2_X1 U687 ( .A1(G952), .A2(n562), .ZN(n773) );
  NOR2_X1 U688 ( .A1(G953), .A2(n773), .ZN(n650) );
  NAND2_X1 U689 ( .A1(G902), .A2(n562), .ZN(n648) );
  INV_X1 U690 ( .A(n648), .ZN(n563) );
  INV_X1 U691 ( .A(G953), .ZN(n782) );
  NOR2_X1 U692 ( .A1(G898), .A2(n782), .ZN(n808) );
  NAND2_X1 U693 ( .A1(n563), .A2(n808), .ZN(n564) );
  XNOR2_X1 U694 ( .A(KEYINPUT95), .B(n564), .ZN(n565) );
  NOR2_X1 U695 ( .A1(n650), .A2(n565), .ZN(n566) );
  INV_X1 U696 ( .A(KEYINPUT0), .ZN(n568) );
  XNOR2_X1 U697 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n581) );
  XNOR2_X1 U698 ( .A(n570), .B(n569), .ZN(n579) );
  XOR2_X1 U699 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n572) );
  NOR2_X1 U700 ( .A1(G953), .A2(G237), .ZN(n603) );
  NAND2_X1 U701 ( .A1(G214), .A2(n603), .ZN(n571) );
  XNOR2_X1 U702 ( .A(n572), .B(n571), .ZN(n575) );
  XOR2_X1 U703 ( .A(n575), .B(n610), .Z(n578) );
  XNOR2_X1 U704 ( .A(n576), .B(G104), .ZN(n577) );
  NOR2_X1 U705 ( .A1(G902), .A2(n791), .ZN(n580) );
  XNOR2_X1 U706 ( .A(n583), .B(n582), .ZN(n590) );
  XNOR2_X1 U707 ( .A(n588), .B(n587), .ZN(n589) );
  NOR2_X1 U708 ( .A1(n630), .A2(n634), .ZN(n591) );
  XNOR2_X1 U709 ( .A(n591), .B(KEYINPUT105), .ZN(n759) );
  INV_X1 U710 ( .A(n697), .ZN(n698) );
  NAND2_X1 U711 ( .A1(G234), .A2(n698), .ZN(n592) );
  XNOR2_X1 U712 ( .A(KEYINPUT20), .B(n592), .ZN(n616) );
  NAND2_X1 U713 ( .A1(n616), .A2(G221), .ZN(n593) );
  XNOR2_X1 U714 ( .A(n593), .B(KEYINPUT21), .ZN(n656) );
  NOR2_X1 U715 ( .A1(n759), .A2(n656), .ZN(n594) );
  INV_X1 U716 ( .A(KEYINPUT75), .ZN(n595) );
  XNOR2_X2 U717 ( .A(n597), .B(n596), .ZN(n637) );
  INV_X1 U718 ( .A(n598), .ZN(n599) );
  NAND2_X1 U719 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U720 ( .A1(n603), .A2(G210), .ZN(n604) );
  INV_X1 U721 ( .A(n640), .ZN(n629) );
  NOR2_X1 U722 ( .A1(n637), .A2(n680), .ZN(n620) );
  XNOR2_X1 U723 ( .A(G119), .B(KEYINPUT82), .ZN(n612) );
  NAND2_X1 U724 ( .A1(n616), .A2(G217), .ZN(n617) );
  NAND2_X1 U725 ( .A1(n620), .A2(n485), .ZN(n621) );
  NOR2_X1 U726 ( .A1(n691), .A2(n621), .ZN(n714) );
  INV_X1 U727 ( .A(n656), .ZN(n743) );
  AND2_X1 U728 ( .A1(n634), .A2(n630), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n829), .A2(KEYINPUT44), .ZN(n635) );
  NAND2_X1 U730 ( .A1(n389), .A2(n626), .ZN(n628) );
  INV_X1 U731 ( .A(n634), .ZN(n632) );
  XOR2_X1 U732 ( .A(n630), .B(KEYINPUT102), .Z(n633) );
  INV_X1 U733 ( .A(n633), .ZN(n631) );
  NAND2_X1 U734 ( .A1(n632), .A2(n631), .ZN(n729) );
  XNOR2_X1 U735 ( .A(n636), .B(KEYINPUT90), .ZN(n646) );
  XOR2_X1 U736 ( .A(n747), .B(KEYINPUT92), .Z(n685) );
  INV_X1 U737 ( .A(n685), .ZN(n638) );
  XNOR2_X1 U738 ( .A(n642), .B(n641), .ZN(n644) );
  NAND2_X1 U739 ( .A1(n642), .A2(n829), .ZN(n643) );
  NAND2_X1 U740 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U741 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n647) );
  INV_X1 U742 ( .A(n481), .ZN(n649) );
  INV_X1 U743 ( .A(n653), .ZN(n763) );
  INV_X1 U744 ( .A(n654), .ZN(n661) );
  NOR2_X1 U745 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U746 ( .A(KEYINPUT73), .B(n657), .ZN(n658) );
  NAND2_X1 U747 ( .A1(n661), .A2(n676), .ZN(n662) );
  XNOR2_X1 U748 ( .A(n664), .B(KEYINPUT77), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n380), .A2(KEYINPUT47), .ZN(n665) );
  NAND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n667) );
  INV_X1 U751 ( .A(n757), .ZN(n670) );
  NOR2_X1 U752 ( .A1(n671), .A2(n670), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n673), .B(n672), .ZN(n695) );
  INV_X1 U754 ( .A(n729), .ZN(n732) );
  NAND2_X1 U755 ( .A1(n695), .A2(n732), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n677), .B(KEYINPUT42), .ZN(n833) );
  NAND2_X1 U757 ( .A1(n831), .A2(n833), .ZN(n679) );
  XOR2_X1 U758 ( .A(KEYINPUT46), .B(KEYINPUT89), .Z(n678) );
  NAND2_X1 U759 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U760 ( .A1(n729), .A2(n682), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n683), .A2(n756), .ZN(n690) );
  NOR2_X1 U762 ( .A1(n693), .A2(n690), .ZN(n684) );
  XNOR2_X1 U763 ( .A(KEYINPUT36), .B(n684), .ZN(n686) );
  NAND2_X1 U764 ( .A1(n686), .A2(n685), .ZN(n738) );
  INV_X1 U765 ( .A(n738), .ZN(n687) );
  NOR2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n689) );
  OR2_X1 U767 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U768 ( .A(n692), .B(KEYINPUT43), .ZN(n694) );
  NAND2_X1 U769 ( .A1(n694), .A2(n693), .ZN(n741) );
  INV_X1 U770 ( .A(n741), .ZN(n696) );
  INV_X1 U771 ( .A(n725), .ZN(n734) );
  AND2_X1 U772 ( .A1(n695), .A2(n734), .ZN(n740) );
  XNOR2_X1 U773 ( .A(KEYINPUT87), .B(n698), .ZN(n699) );
  NAND2_X1 U774 ( .A1(n699), .A2(KEYINPUT2), .ZN(n700) );
  NAND2_X1 U775 ( .A1(n792), .A2(G472), .ZN(n704) );
  XNOR2_X1 U776 ( .A(n363), .B(KEYINPUT62), .ZN(n703) );
  XNOR2_X1 U777 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U778 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n707) );
  INV_X1 U779 ( .A(KEYINPUT91), .ZN(n706) );
  XNOR2_X1 U780 ( .A(n709), .B(n708), .ZN(G57) );
  XOR2_X1 U781 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n712) );
  INV_X1 U782 ( .A(n712), .ZN(n710) );
  XOR2_X1 U783 ( .A(G101), .B(n714), .Z(n715) );
  XNOR2_X1 U784 ( .A(KEYINPUT112), .B(n715), .ZN(G3) );
  XOR2_X1 U785 ( .A(G104), .B(KEYINPUT113), .Z(n717) );
  NAND2_X1 U786 ( .A1(n721), .A2(n732), .ZN(n716) );
  XNOR2_X1 U787 ( .A(n717), .B(n716), .ZN(G6) );
  XOR2_X1 U788 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n719) );
  XNOR2_X1 U789 ( .A(n364), .B(KEYINPUT26), .ZN(n718) );
  XNOR2_X1 U790 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U791 ( .A(KEYINPUT114), .B(n720), .Z(n723) );
  NAND2_X1 U792 ( .A1(n721), .A2(n734), .ZN(n722) );
  XNOR2_X1 U793 ( .A(n723), .B(n722), .ZN(G9) );
  XOR2_X1 U794 ( .A(G110), .B(n724), .Z(G12) );
  NOR2_X1 U795 ( .A1(n380), .A2(n725), .ZN(n727) );
  XNOR2_X1 U796 ( .A(G128), .B(KEYINPUT29), .ZN(n726) );
  XNOR2_X1 U797 ( .A(n727), .B(n726), .ZN(G30) );
  XNOR2_X1 U798 ( .A(n728), .B(G143), .ZN(G45) );
  NOR2_X1 U799 ( .A1(n380), .A2(n729), .ZN(n731) );
  XOR2_X1 U800 ( .A(G146), .B(n731), .Z(G48) );
  NAND2_X1 U801 ( .A1(n370), .A2(n732), .ZN(n733) );
  XNOR2_X1 U802 ( .A(n733), .B(G113), .ZN(G15) );
  NAND2_X1 U803 ( .A1(n370), .A2(n734), .ZN(n736) );
  XNOR2_X1 U804 ( .A(n736), .B(G116), .ZN(G18) );
  XOR2_X1 U805 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n737) );
  XNOR2_X1 U806 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U807 ( .A(G125), .B(n739), .ZN(G27) );
  XOR2_X1 U808 ( .A(G134), .B(n740), .Z(G36) );
  XNOR2_X1 U809 ( .A(G140), .B(n741), .ZN(G42) );
  AND2_X1 U810 ( .A1(n754), .A2(n768), .ZN(n776) );
  XNOR2_X1 U811 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n772) );
  NOR2_X1 U812 ( .A1(n743), .A2(n485), .ZN(n744) );
  XNOR2_X1 U813 ( .A(n744), .B(KEYINPUT49), .ZN(n745) );
  NAND2_X1 U814 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U815 ( .A(KEYINPUT50), .B(n748), .Z(n749) );
  NOR2_X1 U816 ( .A1(n750), .A2(n749), .ZN(n752) );
  NOR2_X1 U817 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U818 ( .A(n753), .B(KEYINPUT51), .ZN(n755) );
  NAND2_X1 U819 ( .A1(n755), .A2(n754), .ZN(n770) );
  NOR2_X1 U820 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U821 ( .A(KEYINPUT117), .B(n758), .ZN(n761) );
  INV_X1 U822 ( .A(n759), .ZN(n760) );
  NAND2_X1 U823 ( .A1(n761), .A2(n760), .ZN(n766) );
  NOR2_X1 U824 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U825 ( .A(KEYINPUT118), .B(n764), .Z(n765) );
  NAND2_X1 U826 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U827 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U828 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U829 ( .A(n772), .B(n771), .ZN(n774) );
  NOR2_X1 U830 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U831 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U832 ( .A(KEYINPUT120), .B(n777), .Z(n780) );
  XOR2_X1 U833 ( .A(n445), .B(KEYINPUT2), .Z(n779) );
  NOR2_X1 U834 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U835 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U836 ( .A(n783), .B(KEYINPUT53), .ZN(n784) );
  XNOR2_X1 U837 ( .A(KEYINPUT121), .B(n784), .ZN(G75) );
  XOR2_X1 U838 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n787) );
  XNOR2_X1 U839 ( .A(n785), .B(KEYINPUT122), .ZN(n786) );
  XNOR2_X1 U840 ( .A(n787), .B(n786), .ZN(n789) );
  NAND2_X1 U841 ( .A1(n792), .A2(G469), .ZN(n788) );
  XNOR2_X1 U842 ( .A(n789), .B(n788), .ZN(n790) );
  NOR2_X1 U843 ( .A1(n803), .A2(n790), .ZN(G54) );
  XOR2_X1 U844 ( .A(n791), .B(KEYINPUT59), .Z(n793) );
  XNOR2_X1 U845 ( .A(n795), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U846 ( .A1(n377), .A2(G478), .ZN(n796) );
  XNOR2_X1 U847 ( .A(n796), .B(KEYINPUT123), .ZN(n798) );
  XOR2_X1 U848 ( .A(n798), .B(n797), .Z(n799) );
  NOR2_X1 U849 ( .A1(n803), .A2(n799), .ZN(G63) );
  NAND2_X1 U850 ( .A1(G217), .A2(n792), .ZN(n800) );
  XNOR2_X1 U851 ( .A(n374), .B(n800), .ZN(n802) );
  NOR2_X1 U852 ( .A1(n803), .A2(n802), .ZN(G66) );
  XOR2_X1 U853 ( .A(n804), .B(G101), .Z(n805) );
  XNOR2_X1 U854 ( .A(n806), .B(n805), .ZN(n807) );
  NOR2_X1 U855 ( .A1(n808), .A2(n807), .ZN(n816) );
  NOR2_X1 U856 ( .A1(G953), .A2(n809), .ZN(n810) );
  XOR2_X1 U857 ( .A(KEYINPUT124), .B(n810), .Z(n814) );
  NAND2_X1 U858 ( .A1(G953), .A2(G224), .ZN(n811) );
  XNOR2_X1 U859 ( .A(KEYINPUT61), .B(n811), .ZN(n812) );
  NAND2_X1 U860 ( .A1(n812), .A2(G898), .ZN(n813) );
  NAND2_X1 U861 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U862 ( .A(n816), .B(n815), .ZN(G69) );
  XNOR2_X1 U863 ( .A(KEYINPUT96), .B(n817), .ZN(n819) );
  XNOR2_X1 U864 ( .A(n819), .B(n818), .ZN(n823) );
  XOR2_X1 U865 ( .A(n823), .B(KEYINPUT125), .Z(n820) );
  XNOR2_X1 U866 ( .A(n446), .B(n820), .ZN(n822) );
  NAND2_X1 U867 ( .A1(n822), .A2(n481), .ZN(n827) );
  XNOR2_X1 U868 ( .A(G227), .B(n823), .ZN(n824) );
  NAND2_X1 U869 ( .A1(n824), .A2(G900), .ZN(n825) );
  NAND2_X1 U870 ( .A1(n825), .A2(G953), .ZN(n826) );
  NAND2_X1 U871 ( .A1(n827), .A2(n826), .ZN(G72) );
  XOR2_X1 U872 ( .A(G119), .B(n828), .Z(G21) );
  XOR2_X1 U873 ( .A(n829), .B(G122), .Z(n830) );
  XNOR2_X1 U874 ( .A(KEYINPUT126), .B(n830), .ZN(G24) );
  XOR2_X1 U875 ( .A(G131), .B(n831), .Z(n832) );
  XNOR2_X1 U876 ( .A(KEYINPUT127), .B(n832), .ZN(G33) );
  XNOR2_X1 U877 ( .A(G137), .B(n833), .ZN(G39) );
endmodule

