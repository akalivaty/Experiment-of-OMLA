//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT66), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n215), .B(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT67), .Z(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n202), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n203), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n229));
  INV_X1    g0029(.A(G97), .ZN(new_n230));
  INV_X1    g0030(.A(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G107), .ZN(new_n232));
  INV_X1    g0032(.A(G264), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT68), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n226), .B(new_n228), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(G116), .ZN(new_n237));
  INV_X1    g0037(.A(G270), .ZN(new_n238));
  OAI221_X1 g0038(.A(new_n236), .B1(new_n235), .B2(new_n234), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(new_n212), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT1), .Z(new_n241));
  NAND2_X1  g0041(.A1(new_n222), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(KEYINPUT69), .Z(G361));
  XNOR2_X1  g0043(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G226), .B(G232), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G250), .B(G257), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G264), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n238), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G358));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G87), .B(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(G107), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(G116), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n255), .B(new_n258), .ZN(G351));
  INV_X1    g0059(.A(G58), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n224), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(new_n201), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n262), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT81), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n210), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n265), .B1(new_n274), .B2(G68), .ZN(new_n275));
  AOI211_X1 g0075(.A(KEYINPUT81), .B(new_n224), .C1(new_n272), .C2(new_n273), .ZN(new_n276));
  OAI211_X1 g0076(.A(KEYINPUT16), .B(new_n264), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT82), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT7), .B1(new_n281), .B2(new_n210), .ZN(new_n282));
  INV_X1    g0082(.A(new_n273), .ZN(new_n283));
  OAI21_X1  g0083(.A(G68), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT81), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n274), .A2(new_n265), .A3(G68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT82), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT16), .A4(new_n264), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n278), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n279), .B2(new_n280), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n268), .A2(KEYINPUT71), .A3(new_n269), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(new_n210), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n283), .B1(new_n294), .B2(new_n271), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n264), .B1(new_n295), .B2(new_n224), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT16), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G1), .A2(G13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n290), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT8), .B(G58), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT74), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n301), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G1), .B2(new_n210), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n307), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n304), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n316));
  INV_X1    g0116(.A(G274), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n268), .A2(new_n269), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G223), .B2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G226), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G41), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n218), .B(KEYINPUT73), .C1(new_n267), .C2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT73), .ZN(new_n327));
  AND2_X1   g0127(.A1(G33), .A2(G41), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n300), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n318), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(G1), .B(G13), .C1(new_n267), .C2(new_n325), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n316), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G232), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n331), .A2(G179), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n331), .B2(new_n335), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT18), .B1(new_n315), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n313), .B1(new_n290), .B2(new_n303), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n342), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT83), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT83), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G190), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n331), .A2(new_n351), .A3(new_n335), .ZN(new_n352));
  AOI21_X1  g0152(.A(G200), .B1(new_n331), .B2(new_n335), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n345), .B1(new_n342), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n302), .B1(new_n289), .B2(new_n278), .ZN(new_n357));
  NOR4_X1   g0157(.A1(new_n357), .A2(KEYINPUT17), .A3(new_n313), .A4(new_n354), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n341), .A2(new_n344), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n267), .A2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G77), .B1(new_n263), .B2(G50), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n210), .B2(G68), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT11), .A3(new_n301), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n224), .B2(new_n309), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n312), .A2(G68), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT12), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT11), .B1(new_n362), .B2(new_n301), .ZN(new_n367));
  OR3_X1    g0167(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT79), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n333), .A2(new_n225), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n318), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n322), .A2(G232), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n292), .B2(new_n293), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n223), .A2(new_n322), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n330), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n372), .B(new_n374), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT13), .ZN(new_n383));
  INV_X1    g0183(.A(new_n377), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n279), .A2(new_n280), .A3(new_n291), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT71), .B1(new_n268), .B2(new_n269), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n379), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n375), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n330), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n372), .A4(new_n374), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n370), .B1(new_n392), .B2(G169), .ZN(new_n393));
  AOI211_X1 g0193(.A(KEYINPUT14), .B(new_n337), .C1(new_n383), .C2(new_n391), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n383), .A2(new_n391), .A3(G179), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n369), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n371), .B1(new_n388), .B2(new_n330), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n390), .B1(new_n398), .B2(new_n374), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n381), .B1(new_n387), .B2(new_n375), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n318), .B(KEYINPUT78), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n400), .A2(KEYINPUT13), .A3(new_n401), .A4(new_n371), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n392), .A2(new_n370), .A3(G169), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n404), .A2(new_n396), .A3(new_n369), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n368), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n368), .B1(new_n392), .B2(G200), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n383), .A2(new_n391), .A3(G190), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(KEYINPUT80), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT80), .ZN(new_n413));
  INV_X1    g0213(.A(new_n368), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n404), .A2(new_n396), .A3(new_n405), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT79), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n406), .ZN(new_n417));
  INV_X1    g0217(.A(new_n411), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n359), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n309), .A2(G50), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n312), .A2(new_n202), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n263), .ZN(new_n426));
  INV_X1    g0226(.A(G150), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n210), .B1(new_n201), .B2(new_n202), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n428), .B(new_n429), .C1(new_n307), .C2(new_n360), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n425), .B(KEYINPUT9), .C1(new_n308), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n292), .A2(new_n293), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G222), .A3(new_n322), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G77), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n432), .A2(KEYINPUT72), .A3(G222), .A4(new_n322), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(G223), .A3(G1698), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n435), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n318), .B1(new_n440), .B2(new_n330), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n334), .A2(G226), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(G190), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT9), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n423), .B(KEYINPUT75), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n430), .A2(new_n308), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n431), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n441), .A2(new_n442), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G200), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n450), .C1(KEYINPUT77), .C2(KEYINPUT10), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT10), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n431), .A2(new_n443), .A3(new_n447), .A4(KEYINPUT77), .ZN(new_n453));
  INV_X1    g0253(.A(new_n450), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n431), .A2(new_n443), .A3(new_n447), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n449), .ZN(new_n457));
  INV_X1    g0257(.A(G179), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n425), .B1(new_n308), .B2(new_n430), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n460), .C1(G169), .C2(new_n457), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n451), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n432), .A2(G238), .A3(G1698), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n432), .A2(G232), .A3(new_n322), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n464), .C1(new_n232), .C2(new_n432), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n330), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n333), .A2(new_n227), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n318), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n470), .A2(new_n337), .ZN(new_n471));
  XOR2_X1   g0271(.A(KEYINPUT15), .B(G87), .Z(new_n472));
  AND2_X1   g0272(.A1(new_n472), .A2(new_n360), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n305), .A2(new_n426), .B1(new_n210), .B2(new_n203), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n301), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n310), .A2(G77), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n476), .C1(G77), .C2(new_n312), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n470), .B2(G179), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n470), .A2(G200), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT76), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n481), .B(new_n483), .C1(new_n346), .C2(new_n470), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n477), .A2(new_n482), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n462), .A2(new_n480), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n420), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n210), .B(G87), .C1(new_n385), .C2(new_n386), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT22), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  AOI21_X1  g0294(.A(G20), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n210), .A2(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT23), .ZN(new_n498));
  AND4_X1   g0298(.A1(new_n489), .A2(new_n492), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n490), .B2(new_n491), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n489), .B1(new_n500), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n301), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n231), .A2(G1698), .ZN(new_n503));
  OAI221_X1 g0303(.A(new_n503), .B1(G250), .B2(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n504));
  INV_X1    g0304(.A(G294), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n267), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n330), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G41), .ZN(new_n510));
  INV_X1    g0310(.A(G45), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G1), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n325), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n317), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(G264), .A3(new_n332), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT89), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n514), .A2(KEYINPUT89), .A3(G264), .A4(new_n332), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n507), .A2(new_n516), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G200), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n507), .A2(new_n346), .A3(new_n516), .A4(new_n517), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n312), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n267), .A2(G1), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n526), .A2(new_n301), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(new_n232), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT25), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n502), .A2(new_n525), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n263), .A2(G77), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n232), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n230), .A2(new_n232), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n206), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n534), .B(new_n539), .C1(new_n295), .C2(new_n232), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n301), .B1(new_n230), .B2(new_n526), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n528), .A2(G97), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n322), .A2(KEYINPUT4), .A3(G244), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G250), .A2(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n432), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(new_n322), .C1(new_n279), .C2(new_n280), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n547), .A2(new_n548), .B1(G33), .B2(G283), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n381), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n514), .A2(G257), .A3(new_n332), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n550), .A2(new_n515), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n547), .A2(new_n548), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n292), .A2(new_n293), .B1(new_n543), .B2(new_n544), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n330), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n516), .A3(new_n551), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G190), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n541), .B(new_n542), .C1(new_n554), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n540), .A2(new_n301), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n526), .A2(new_n230), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n542), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n559), .A2(G179), .A3(new_n516), .A4(new_n551), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n553), .B2(new_n337), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n533), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n514), .A2(G270), .A3(new_n332), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n292), .A2(new_n293), .A3(G303), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n233), .A2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n320), .B(new_n572), .C1(G257), .C2(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n574), .B2(new_n330), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n516), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n526), .A2(new_n237), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n528), .A2(G116), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n556), .B(new_n210), .C1(G33), .C2(new_n230), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n301), .C1(new_n210), .C2(G116), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT20), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n577), .B(new_n578), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n584), .A3(G169), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n571), .A2(new_n573), .B1(new_n329), .B2(new_n326), .ZN(new_n589));
  NOR4_X1   g0389(.A1(new_n589), .A2(new_n458), .A3(new_n515), .A4(new_n570), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n337), .B1(new_n575), .B2(new_n516), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(KEYINPUT21), .ZN(new_n592));
  INV_X1    g0392(.A(new_n584), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT88), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT88), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n589), .A2(new_n515), .A3(new_n570), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n596), .A2(new_n586), .A3(new_n337), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n584), .C1(new_n597), .C2(new_n590), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n588), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT85), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n511), .B2(G1), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n209), .A2(KEYINPUT85), .A3(G45), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n332), .A2(G250), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G250), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n209), .A2(G45), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(KEYINPUT86), .A3(new_n332), .A4(new_n602), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n512), .A2(G274), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n225), .A2(new_n322), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n227), .A2(G1698), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n279), .C2(new_n280), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n494), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n330), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n210), .B1(new_n375), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G87), .B2(new_n207), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n375), .B2(G20), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n210), .B(G68), .C1(new_n279), .C2(new_n280), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n472), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n624), .A2(new_n301), .B1(new_n526), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n528), .A2(G87), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n605), .A2(new_n609), .B1(new_n330), .B2(new_n615), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(G190), .A3(new_n611), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n618), .A2(new_n626), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(G179), .A2(new_n610), .A3(new_n611), .A4(new_n616), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n337), .B1(new_n628), .B2(new_n611), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n301), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n625), .A2(new_n526), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n528), .A2(new_n472), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT87), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n626), .A2(new_n639), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n630), .B1(new_n633), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n502), .A2(new_n529), .A3(new_n532), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n507), .A2(new_n516), .A3(new_n517), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n644), .A2(new_n337), .B1(new_n521), .B2(new_n458), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n596), .A2(new_n350), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n593), .C1(new_n522), .C2(new_n596), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n569), .A2(new_n599), .A3(new_n646), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n488), .A2(new_n649), .ZN(G372));
  INV_X1    g0450(.A(new_n461), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n418), .A2(new_n479), .ZN(new_n652));
  OAI22_X1  g0452(.A1(new_n417), .A2(new_n652), .B1(new_n356), .B2(new_n358), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n343), .B1(new_n342), .B2(new_n339), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT18), .B(new_n340), .C1(new_n357), .C2(new_n313), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n451), .A2(new_n456), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n651), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n617), .A2(G169), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n628), .A2(G179), .A3(new_n611), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n637), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n638), .A3(new_n640), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(new_n565), .A3(new_n567), .A4(new_n630), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n618), .A2(new_n629), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n626), .A2(KEYINPUT90), .A3(new_n627), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT90), .B1(new_n626), .B2(new_n627), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n668), .A2(new_n671), .B1(new_n662), .B2(new_n637), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n565), .A2(new_n567), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n565), .B2(new_n567), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n667), .B(new_n672), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n643), .B2(new_n645), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n672), .A2(new_n533), .A3(new_n562), .A4(new_n568), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n666), .B(new_n676), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n659), .B1(new_n488), .B2(new_n681), .ZN(G369));
  INV_X1    g0482(.A(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G20), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n209), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n599), .B(new_n648), .C1(new_n593), .C2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n677), .A2(new_n584), .A3(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n643), .A2(new_n645), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n533), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n643), .A2(new_n690), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n698), .B2(new_n691), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n599), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n533), .B(new_n691), .C1(new_n703), .C2(new_n697), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n213), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n706), .A2(KEYINPUT92), .A3(G41), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT92), .B1(new_n706), .B2(G41), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n220), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n663), .B1(new_n714), .B2(KEYINPUT26), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n703), .A2(new_n697), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n715), .B1(KEYINPUT26), .B2(new_n665), .C1(new_n716), .C2(new_n679), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n680), .A2(new_n691), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n507), .A2(new_n519), .A3(new_n520), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n617), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT93), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n722), .B2(new_n617), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n724), .A2(new_n590), .A3(new_n553), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n560), .B1(new_n723), .B2(KEYINPUT93), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n590), .A4(new_n726), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n617), .B(KEYINPUT94), .Z(new_n732));
  NOR2_X1   g0532(.A1(new_n553), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n576), .A3(new_n521), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n690), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT31), .B(new_n736), .C1(new_n649), .C2(new_n690), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(KEYINPUT31), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n718), .A2(new_n721), .B1(new_n739), .B2(G330), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n713), .B1(new_n740), .B2(G1), .ZN(G364));
  AOI21_X1  g0541(.A(new_n209), .B1(new_n684), .B2(G45), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n709), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT96), .Z(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n694), .A2(G330), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n696), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n255), .A2(G45), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n706), .A2(new_n320), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n748), .B(new_n749), .C1(G45), .C2(new_n220), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n432), .A2(new_n213), .A3(G355), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n750), .B(new_n751), .C1(G116), .C2(new_n213), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n300), .B1(G20), .B2(new_n337), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n755), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n694), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n756), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n210), .A2(new_n458), .A3(new_n522), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n350), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT98), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n346), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n210), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(G326), .B1(G294), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT99), .Z(new_n770));
  NAND2_X1  g0570(.A1(new_n762), .A2(new_n346), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G317), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT33), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n773), .A2(KEYINPUT33), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n210), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(new_n346), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n210), .A2(new_n458), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n776), .B1(new_n777), .B2(new_n779), .C1(new_n780), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n778), .A2(new_n782), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n432), .B1(G329), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G303), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n350), .A2(new_n522), .A3(new_n781), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n770), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n767), .A2(new_n230), .ZN(new_n795));
  INV_X1    g0595(.A(new_n789), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(G87), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n260), .B2(new_n793), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n436), .B(new_n798), .C1(G68), .C2(new_n772), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n800));
  INV_X1    g0600(.A(G159), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n785), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n779), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G107), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n785), .B2(new_n801), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n783), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n802), .B(new_n806), .C1(G77), .C2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n799), .B(new_n808), .C1(new_n202), .C2(new_n763), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n761), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n744), .B1(new_n760), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n747), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT100), .Z(G396));
  NAND2_X1  g0613(.A1(new_n739), .A2(G330), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n471), .A2(new_n478), .A3(new_n690), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n477), .A2(new_n690), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n484), .B2(new_n485), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n817), .B2(new_n479), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n719), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n814), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n745), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n436), .B1(new_n780), .B2(new_n785), .ZN(new_n822));
  INV_X1    g0622(.A(G87), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n779), .A2(new_n823), .B1(new_n789), .B2(new_n232), .ZN(new_n824));
  INV_X1    g0624(.A(new_n793), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(G294), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n237), .B2(new_n783), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n822), .B(new_n827), .C1(G97), .C2(new_n768), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n772), .A2(KEYINPUT101), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n772), .A2(KEYINPUT101), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n828), .B1(new_n777), .B2(new_n831), .C1(new_n788), .C2(new_n763), .ZN(new_n832));
  INV_X1    g0632(.A(new_n763), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G137), .B1(G159), .B2(new_n807), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT102), .B(G143), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n427), .B2(new_n771), .C1(new_n793), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n779), .A2(new_n224), .B1(new_n789), .B2(new_n202), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n281), .B(new_n839), .C1(G58), .C2(new_n768), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n838), .B(new_n840), .C1(new_n841), .C2(new_n785), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n745), .B1(new_n843), .B2(new_n756), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n756), .A2(new_n753), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(G77), .B2(new_n846), .C1(new_n754), .C2(new_n818), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n821), .A2(new_n847), .ZN(G384));
  INV_X1    g0648(.A(new_n688), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n359), .A2(new_n315), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n342), .B1(new_n339), .B2(new_n688), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n304), .A2(new_n314), .A3(new_n355), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n315), .B1(new_n340), .B2(new_n849), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n852), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n850), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT107), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(KEYINPUT17), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n342), .A2(new_n345), .A3(new_n355), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n861), .A2(new_n862), .B1(new_n654), .B2(new_n655), .ZN(new_n863));
  INV_X1    g0663(.A(new_n264), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n285), .B2(new_n286), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n301), .B1(new_n865), .B2(KEYINPUT16), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT106), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n301), .C1(new_n865), .C2(KEYINPUT16), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n290), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n688), .B1(new_n870), .B2(new_n314), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n860), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n359), .A2(KEYINPUT107), .A3(new_n871), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n870), .A2(new_n314), .B1(new_n339), .B2(new_n688), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n875), .B2(new_n853), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n873), .A2(new_n874), .B1(new_n857), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n859), .B1(new_n877), .B2(KEYINPUT38), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n737), .A2(new_n738), .A3(new_n818), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n411), .B1(new_n414), .B2(new_n691), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n408), .A2(KEYINPUT105), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n417), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n408), .A2(new_n691), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT40), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n737), .A2(new_n738), .A3(new_n818), .ZN(new_n889));
  INV_X1    g0689(.A(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n416), .A2(new_n406), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n882), .B1(new_n891), .B2(new_n368), .ZN(new_n892));
  AOI211_X1 g0692(.A(KEYINPUT105), .B(new_n414), .C1(new_n416), .C2(new_n406), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n885), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n876), .A2(new_n857), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n897), .B(new_n898), .C1(new_n873), .C2(new_n874), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n873), .A2(new_n874), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n876), .A2(new_n857), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n888), .B(new_n896), .C1(new_n899), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n420), .A2(new_n487), .A3(new_n739), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n904), .B(new_n905), .Z(new_n906));
  INV_X1    g0706(.A(G330), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n881), .A2(new_n883), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(new_n690), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n900), .A2(new_n901), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n897), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n863), .A2(new_n860), .A3(new_n872), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT107), .B1(new_n359), .B2(new_n871), .ZN(new_n915));
  OAI211_X1 g0715(.A(KEYINPUT38), .B(new_n901), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n911), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n850), .A2(new_n858), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n897), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(KEYINPUT39), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n910), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n656), .A2(new_n849), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n885), .B1(new_n909), .B2(new_n890), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n680), .A2(new_n691), .A3(new_n818), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  INV_X1    g0728(.A(new_n815), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n926), .B1(new_n930), .B2(new_n931), .C1(new_n899), .C2(new_n902), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n922), .A2(new_n924), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n718), .A2(new_n420), .A3(new_n487), .A4(new_n721), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n659), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n908), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n209), .B2(new_n684), .ZN(new_n938));
  OAI211_X1 g0738(.A(G20), .B(new_n218), .C1(new_n538), .C2(KEYINPUT35), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n237), .B(new_n939), .C1(KEYINPUT35), .C2(new_n538), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT36), .Z(new_n941));
  NOR3_X1   g0741(.A1(new_n261), .A2(new_n220), .A3(new_n203), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT103), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n224), .A2(G50), .ZN(new_n944));
  OAI211_X1 g0744(.A(G1), .B(new_n683), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n941), .A3(new_n945), .ZN(G367));
  OAI22_X1  g0746(.A1(new_n260), .A2(new_n789), .B1(new_n783), .B2(new_n202), .ZN(new_n947));
  INV_X1    g0747(.A(G137), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n432), .B1(new_n948), .B2(new_n785), .C1(new_n793), .C2(new_n427), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n947), .B(new_n949), .C1(G68), .C2(new_n768), .ZN(new_n950));
  INV_X1    g0750(.A(new_n831), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n951), .A2(G159), .B1(new_n765), .B2(new_n835), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n803), .A2(G77), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT112), .Z(new_n955));
  NOR2_X1   g0755(.A1(new_n783), .A2(new_n777), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n951), .A2(G294), .B1(G311), .B2(new_n765), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n281), .B1(new_n785), .B2(new_n773), .C1(new_n230), .C2(new_n779), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT111), .Z(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT46), .B1(new_n796), .B2(G116), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT110), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n796), .A2(KEYINPUT46), .A3(G116), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n232), .B2(new_n767), .C1(new_n793), .C2(new_n788), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n955), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n745), .B1(new_n967), .B2(new_n756), .ZN(new_n968));
  INV_X1    g0768(.A(new_n749), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n757), .B1(new_n213), .B2(new_n625), .C1(new_n251), .C2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n671), .A2(new_n691), .ZN(new_n971));
  MUX2_X1   g0771(.A(new_n672), .B(new_n663), .S(new_n971), .Z(new_n972));
  OAI211_X1 g0772(.A(new_n968), .B(new_n970), .C1(new_n759), .C2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n742), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n568), .A2(new_n691), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n565), .A2(new_n690), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n562), .A2(new_n568), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n704), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT45), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(new_n704), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT44), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n702), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n703), .A2(new_n691), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(new_n699), .ZN(new_n987));
  INV_X1    g0787(.A(new_n986), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n701), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n696), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n985), .A2(new_n740), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n740), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n709), .B(KEYINPUT41), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n974), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n979), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT42), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n568), .B1(new_n995), .B2(new_n698), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n691), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n997), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT109), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1000), .B(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n702), .A2(new_n995), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n973), .B1(new_n994), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT113), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(G387));
  NOR2_X1   g0808(.A1(new_n305), .A2(G50), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT50), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n710), .B1(new_n224), .B2(new_n203), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g0811(.A(G45), .B(new_n1011), .C1(new_n1010), .C2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n749), .B1(new_n248), .B2(new_n511), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n436), .A2(new_n706), .A3(new_n710), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n213), .A2(G107), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n757), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n744), .B(new_n1017), .C1(new_n701), .C2(new_n759), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n765), .A2(G322), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n780), .B2(new_n831), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n788), .B2(new_n783), .C1(new_n773), .C2(new_n793), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n768), .A2(G283), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n796), .A2(G294), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n786), .A2(G326), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n320), .B1(new_n803), .B2(G116), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n625), .A2(new_n767), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n793), .A2(new_n202), .B1(new_n763), .B2(new_n801), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G97), .C2(new_n803), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G77), .A2(new_n796), .B1(new_n807), .B2(G68), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n427), .B2(new_n785), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n307), .B2(new_n772), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(new_n1038), .A3(new_n320), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1018), .B1(new_n1040), .B2(new_n756), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT115), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n974), .B2(new_n990), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n990), .A2(new_n740), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n709), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n990), .A2(new_n740), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1043), .A2(new_n1047), .ZN(G393));
  XNOR2_X1  g0848(.A(new_n985), .B(new_n1046), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n1045), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n985), .A2(new_n974), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n995), .A2(new_n755), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT116), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n436), .B1(new_n792), .B2(new_n785), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n804), .B1(new_n777), .B2(new_n789), .C1(new_n505), .C2(new_n783), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n951), .C2(G303), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n793), .A2(new_n780), .B1(new_n763), .B2(new_n773), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n237), .C2(new_n767), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n320), .B1(new_n779), .B2(new_n823), .C1(new_n836), .C2(new_n785), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n224), .A2(new_n789), .B1(new_n783), .B2(new_n305), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n951), .C2(G50), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n768), .A2(G77), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n793), .A2(new_n801), .B1(new_n763), .B2(new_n427), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n761), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n258), .A2(new_n749), .B1(G97), .B2(new_n706), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n745), .B(new_n1067), .C1(new_n757), .C2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT117), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n1053), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1050), .A2(new_n1051), .A3(new_n1071), .ZN(G390));
  OAI21_X1  g0872(.A(KEYINPUT39), .B1(new_n899), .B2(new_n902), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n910), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n930), .A2(new_n931), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n925), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n878), .A2(new_n911), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n817), .A2(new_n479), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n717), .A2(new_n691), .A3(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1080), .A2(new_n929), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1074), .B(new_n920), .C1(new_n1081), .C2(new_n925), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n879), .B(G330), .C1(new_n884), .C2(new_n885), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1078), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n737), .A2(new_n738), .A3(G330), .A4(new_n818), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n894), .A2(new_n1089), .A3(new_n895), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1081), .A2(new_n1084), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n896), .A2(G330), .B1(new_n925), .B2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n1075), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n420), .A2(G330), .A3(new_n487), .A4(new_n739), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT118), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n934), .A2(new_n1094), .A3(new_n1095), .A4(new_n659), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n934), .A2(new_n1094), .A3(new_n659), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT118), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1093), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1088), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT119), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT119), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1088), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1102), .A2(new_n1104), .A3(new_n1045), .A4(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1088), .A2(new_n742), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n917), .A2(new_n921), .A3(new_n754), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n307), .A2(new_n846), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n436), .B1(new_n224), .B2(new_n779), .C1(new_n505), .C2(new_n785), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n951), .B2(G107), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1063), .B1(new_n230), .B2(new_n783), .C1(new_n763), .C2(new_n777), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G116), .B2(new_n825), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n823), .C2(new_n789), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  AOI22_X1  g0915(.A1(new_n833), .A2(G128), .B1(new_n807), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n841), .B2(new_n793), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n432), .B1(new_n1118), .B2(new_n785), .C1(new_n801), .C2(new_n767), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n202), .B2(new_n779), .C1(new_n948), .C2(new_n831), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n796), .A2(G150), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1114), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1124), .A2(new_n756), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1108), .A2(new_n745), .A3(new_n1109), .A4(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1107), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1106), .A2(new_n1127), .ZN(G378));
  OAI211_X1 g0928(.A(new_n879), .B(new_n888), .C1(new_n884), .C2(new_n885), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n916), .B2(new_n913), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n888), .B1(new_n920), .B2(new_n896), .ZN(new_n1131));
  OAI21_X1  g0931(.A(G330), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT56), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n460), .A2(new_n849), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n462), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT55), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n451), .A2(new_n456), .A3(new_n461), .A4(new_n1134), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT55), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(KEYINPUT56), .A3(new_n1139), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1132), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n904), .A2(G330), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(KEYINPUT122), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1074), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n925), .B(new_n1075), .C1(new_n916), .C2(new_n913), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n923), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1147), .A2(new_n933), .A3(KEYINPUT122), .A4(new_n1149), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1098), .A2(new_n1096), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1105), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(KEYINPUT123), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT123), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1154), .A2(new_n1155), .B1(new_n1157), .B2(new_n1105), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(KEYINPUT57), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1148), .B1(new_n904), .B2(G330), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n907), .B(new_n1146), .C1(new_n887), .C2(new_n903), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1153), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1147), .A2(new_n933), .A3(new_n1149), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1157), .A2(new_n1105), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n709), .B1(new_n1169), .B2(KEYINPUT57), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1161), .A2(new_n1164), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1148), .A2(new_n753), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n845), .A2(new_n202), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n325), .B(new_n281), .C1(new_n785), .C2(new_n777), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n771), .A2(new_n230), .B1(new_n203), .B2(new_n789), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G68), .C2(new_n768), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n803), .A2(G58), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n237), .B2(new_n763), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n472), .B2(new_n807), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(new_n232), .C2(new_n793), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n202), .B1(new_n279), .B2(G41), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n763), .A2(new_n1118), .B1(new_n771), .B2(new_n841), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G137), .B2(new_n807), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n796), .A2(new_n1115), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n825), .A2(G128), .B1(G150), .B2(new_n768), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT59), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G33), .B1(new_n786), .B2(G124), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n325), .C1(new_n801), .C2(new_n779), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT121), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1182), .B(new_n1183), .C1(new_n1189), .C2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n745), .B1(new_n1193), .B2(new_n756), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1172), .A2(new_n1173), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1156), .B2(new_n974), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1171), .A2(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1093), .A2(new_n974), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n951), .A2(new_n1115), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n796), .A2(G159), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n768), .A2(G50), .B1(new_n807), .B2(G150), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1200), .A2(new_n1177), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n793), .A2(new_n948), .B1(new_n763), .B2(new_n841), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n786), .A2(G128), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n320), .A3(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n825), .A2(G283), .B1(G97), .B2(new_n796), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n807), .A2(G107), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n833), .A2(G294), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n953), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n432), .B(new_n1033), .C1(G303), .C2(new_n786), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n237), .B2(new_n831), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1203), .A2(new_n1207), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n745), .B1(new_n1214), .B2(new_n756), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(G68), .B2(new_n846), .C1(new_n926), .C2(new_n754), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1199), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1100), .A2(new_n993), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1157), .A2(new_n1093), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(G381));
  NOR2_X1   g1021(.A1(G375), .A2(G378), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(G396), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1043), .A2(new_n1224), .A3(new_n1047), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(G390), .ZN(new_n1226));
  OR2_X1    g1026(.A1(G381), .A2(G384), .ZN(new_n1227));
  OR4_X1    g1027(.A1(G387), .A2(new_n1223), .A3(new_n1226), .A4(new_n1227), .ZN(G407));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1045), .B(new_n1100), .C1(new_n1220), .C2(KEYINPUT60), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1157), .A2(new_n1093), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1220), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1232), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n821), .B(new_n847), .C1(new_n1238), .C2(new_n1217), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1237), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT125), .B1(new_n1220), .B2(KEYINPUT60), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G384), .B(new_n1218), .C1(new_n1242), .C2(new_n1232), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1171), .A2(G378), .A3(new_n1197), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n933), .B1(new_n1246), .B2(KEYINPUT122), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1155), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n993), .B(new_n1158), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT124), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n974), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1156), .A2(new_n1253), .A3(new_n993), .A4(new_n1158), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1195), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G378), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1231), .B(new_n1244), .C1(new_n1245), .C2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT63), .B1(new_n1258), .B2(KEYINPUT126), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G393), .A2(G396), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT113), .B1(new_n1260), .B2(new_n1225), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(G390), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1225), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(G390), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1006), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1006), .C1(G390), .C2(new_n1261), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1245), .A2(new_n1257), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1231), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1231), .A2(G2897), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1244), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1239), .A2(new_n1243), .A3(new_n1272), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1269), .A2(new_n1270), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1259), .A2(new_n1268), .A3(new_n1277), .A4(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1231), .B1(new_n1245), .B2(new_n1257), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1286), .B2(new_n1278), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1284), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1283), .B1(new_n1291), .B2(new_n1268), .ZN(G405));
  NAND3_X1  g1092(.A1(new_n1278), .A2(G375), .A3(new_n1256), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1278), .B1(new_n1256), .B2(G375), .ZN(new_n1295));
  OAI211_X1 g1095(.A(KEYINPUT127), .B(new_n1245), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1256), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1244), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1245), .A2(KEYINPUT127), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1293), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1268), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1296), .A2(new_n1268), .A3(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(G402));
endmodule


