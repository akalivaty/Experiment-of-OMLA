//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G127gat), .ZN(new_n209));
  INV_X1    g008(.A(G127gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G134gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n206), .A2(new_n207), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n211), .ZN(new_n213));
  XNOR2_X1  g012(.A(G113gat), .B(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n217), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n238), .A3(new_n231), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n230), .B2(new_n231), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n229), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n229), .B(KEYINPUT67), .C1(new_n240), .C2(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT23), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n221), .A2(KEYINPUT25), .A3(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n236), .A2(new_n237), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n217), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n219), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n230), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(G183gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT68), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n262), .B2(KEYINPUT27), .ZN(new_n265));
  INV_X1    g064(.A(G190gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n259), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT69), .B(new_n259), .C1(new_n264), .C2(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT27), .B(G183gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT28), .A3(new_n266), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n258), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n216), .B1(new_n251), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n266), .B(new_n265), .C1(new_n273), .C2(KEYINPUT68), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT69), .B1(new_n277), .B2(new_n259), .ZN(new_n278));
  INV_X1    g077(.A(new_n271), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n258), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n216), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n235), .A2(new_n233), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n217), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n234), .B1(new_n287), .B2(new_n221), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n237), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n245), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n239), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT67), .B1(new_n292), .B2(new_n229), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n250), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n282), .A2(new_n283), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT34), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n305), .A3(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n299), .B2(new_n300), .ZN(new_n308));
  AOI211_X1 g107(.A(KEYINPUT73), .B(KEYINPUT34), .C1(new_n298), .C2(KEYINPUT72), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n297), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n251), .A2(new_n275), .A3(new_n216), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n283), .B1(new_n282), .B2(new_n295), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT33), .ZN(new_n316));
  XNOR2_X1  g115(.A(G15gat), .B(G43gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n315), .B(KEYINPUT32), .C1(new_n316), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n315), .B2(KEYINPUT32), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(new_n316), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n319), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n297), .B1(new_n276), .B2(new_n296), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n276), .A2(new_n296), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT33), .B1(new_n329), .B2(new_n312), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n328), .A2(KEYINPUT71), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n320), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G228gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  AND2_X1   g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n340), .B1(new_n343), .B2(KEYINPUT75), .ZN(new_n344));
  XNOR2_X1  g143(.A(G141gat), .B(G148gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n340), .B2(new_n338), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n345), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n338), .A2(new_n340), .ZN(new_n352));
  NAND2_X1  g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n343), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  INV_X1    g158(.A(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G218gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n358), .A3(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n357), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  INV_X1    g170(.A(new_n367), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n364), .B1(new_n362), .B2(new_n358), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n356), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n348), .A2(new_n357), .A3(new_n351), .A4(new_n355), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n371), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n372), .A2(new_n373), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n336), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n336), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n356), .B2(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n356), .A2(new_n368), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n379), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n377), .B2(new_n371), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(G22gat), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n351), .A2(new_n355), .ZN(new_n390));
  INV_X1    g189(.A(new_n339), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT2), .B1(new_n345), .B2(new_n346), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n343), .A2(KEYINPUT75), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n374), .B2(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n368), .A2(new_n369), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n382), .B1(new_n398), .B2(new_n387), .ZN(new_n399));
  INV_X1    g198(.A(G22gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n384), .A3(new_n383), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G78gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n389), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n389), .B2(new_n402), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  INV_X1    g206(.A(G106gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n389), .A2(new_n402), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G78gat), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n413), .B2(new_n404), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT71), .B1(new_n328), .B2(new_n330), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n315), .A2(KEYINPUT32), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n417), .A2(new_n323), .A3(new_n321), .A4(new_n325), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n419), .A2(new_n307), .A3(new_n310), .A4(new_n320), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n333), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n283), .B1(new_n356), .B2(KEYINPUT3), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n377), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n351), .A2(new_n355), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n283), .A3(new_n348), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n395), .A2(new_n429), .A3(new_n283), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n283), .B1(new_n426), .B2(new_n348), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n390), .A2(new_n394), .A3(new_n216), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n423), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT77), .B1(new_n435), .B2(KEYINPUT5), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n216), .B1(new_n390), .B2(new_n394), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n422), .B1(new_n427), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT77), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n430), .A3(KEYINPUT78), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n444), .A3(KEYINPUT4), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n377), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n443), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT0), .ZN(new_n451));
  XNOR2_X1  g250(.A(G57gat), .B(G85gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n442), .A2(new_n453), .A3(new_n448), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT79), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n442), .A2(new_n459), .A3(new_n453), .A4(new_n448), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n435), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(new_n463), .B1(new_n431), .B2(new_n425), .ZN(new_n464));
  INV_X1    g263(.A(new_n448), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n454), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n468), .A3(new_n454), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n455), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G64gat), .B(G92gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n472), .B(new_n473), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT74), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n282), .A2(new_n295), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(new_n371), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n280), .A2(new_n281), .B1(new_n289), .B2(new_n294), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(new_n477), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n480), .A2(new_n482), .A3(new_n379), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n477), .B1(new_n481), .B2(KEYINPUT29), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n478), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n386), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n475), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n379), .B1(new_n480), .B2(new_n482), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n386), .A3(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n474), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n488), .A2(new_n489), .A3(new_n492), .A4(new_n474), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n471), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT35), .B1(new_n421), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n457), .A2(new_n458), .A3(new_n466), .A4(new_n460), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n455), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT35), .B1(new_n491), .B2(new_n493), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n500), .A2(new_n415), .A3(new_n420), .A4(new_n333), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n415), .B1(new_n471), .B2(new_n494), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504));
  AND4_X1   g303(.A1(new_n320), .A2(new_n419), .A3(new_n307), .A4(new_n310), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n320), .A2(new_n419), .B1(new_n307), .B2(new_n310), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n333), .A2(KEYINPUT36), .A3(new_n420), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n489), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT37), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT37), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n489), .A3(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n512), .A2(new_n513), .A3(new_n475), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n490), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n498), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n490), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n515), .A2(new_n513), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n474), .B1(new_n511), .B2(KEYINPUT37), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(KEYINPUT84), .A3(new_n455), .A4(new_n497), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n515), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n518), .A2(new_n523), .B1(new_n526), .B2(KEYINPUT38), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n446), .A2(new_n445), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n422), .B1(new_n529), .B2(new_n443), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n427), .A2(new_n437), .A3(new_n422), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT39), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n454), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT40), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n528), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT83), .A4(KEYINPUT40), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n494), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n537), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n466), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n415), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n509), .A2(KEYINPUT82), .B1(new_n527), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n546));
  AOI211_X1 g345(.A(new_n546), .B(new_n503), .C1(new_n508), .C2(new_n507), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n502), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT16), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(G1gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G1gat), .B2(new_n550), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(G8gat), .Z(new_n554));
  XOR2_X1   g353(.A(G43gat), .B(G50gat), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G29gat), .ZN(new_n558));
  INV_X1    g357(.A(G36gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(G29gat), .A2(G36gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT14), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n555), .A2(new_n556), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n564), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n561), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n557), .B1(new_n560), .B2(new_n563), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n554), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT89), .ZN(new_n575));
  INV_X1    g374(.A(new_n554), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(new_n570), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT90), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT18), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n554), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n575), .B(KEYINPUT13), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G169gat), .B(G197gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n582), .A2(new_n584), .A3(new_n590), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT92), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n581), .A2(KEYINPUT18), .B1(new_n587), .B2(new_n589), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n584), .A4(new_n596), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n584), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n596), .B(KEYINPUT87), .Z(new_n605));
  AND3_X1   g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n610));
  INV_X1    g409(.A(new_n572), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G99gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT8), .B1(new_n614), .B2(new_n408), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT93), .B(G92gat), .Z(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n625), .A3(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT95), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(new_n585), .ZN(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n610), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  AOI211_X1 g438(.A(KEYINPUT97), .B(new_n639), .C1(new_n632), .C2(new_n635), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n632), .A2(new_n635), .A3(new_n639), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n643), .B(KEYINPUT96), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n650), .B2(new_n641), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n637), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT97), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n610), .A3(new_n637), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT98), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n649), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G57gat), .B(G64gat), .Z(new_n658));
  INV_X1    g457(.A(G71gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n403), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(KEYINPUT9), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G71gat), .B(G78gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g462(.A(KEYINPUT21), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G127gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n554), .B1(new_n664), .B2(new_n663), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n671));
  INV_X1    g470(.A(G155gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(G183gat), .B(G211gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n670), .B(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n657), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n663), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n624), .A2(new_n681), .A3(new_n626), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n624), .B2(new_n626), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(KEYINPUT100), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n624), .A2(new_n681), .A3(new_n626), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT10), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n683), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT10), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n689), .A2(new_n679), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n684), .A2(KEYINPUT100), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n685), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n685), .A2(new_n692), .A3(new_n697), .A4(new_n693), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR4_X1   g500(.A1(new_n549), .A2(new_n609), .A3(new_n678), .A4(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n471), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  AND3_X1   g505(.A1(new_n702), .A2(new_n541), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G8gat), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n702), .B2(new_n541), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT42), .B2(new_n707), .ZN(G1325gat));
  INV_X1    g510(.A(G15gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n505), .A2(new_n506), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n702), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n507), .A2(new_n508), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n702), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(new_n712), .ZN(G1326gat));
  INV_X1    g517(.A(new_n415), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT43), .B(G22gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  NOR2_X1   g521(.A1(new_n655), .A2(KEYINPUT98), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n650), .A2(new_n641), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n646), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n642), .B1(new_n641), .B2(new_n648), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n677), .A2(new_n701), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n548), .A2(new_n608), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(G29gat), .A3(new_n471), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT45), .Z(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n657), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n548), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n728), .A2(new_n608), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT101), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n502), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n496), .A2(new_n501), .A3(KEYINPUT102), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n518), .A2(new_n523), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n526), .A2(KEYINPUT38), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n415), .A3(new_n543), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n509), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n657), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n734), .B(new_n736), .C1(new_n746), .C2(KEYINPUT44), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n738), .A2(new_n739), .B1(new_n744), .B2(new_n509), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n732), .B1(new_n750), .B2(new_n657), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n751), .A2(KEYINPUT103), .A3(new_n734), .A4(new_n736), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n749), .A2(new_n703), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n731), .B1(new_n558), .B2(new_n753), .ZN(G1328gat));
  NOR3_X1   g553(.A1(new_n729), .A2(G36gat), .A3(new_n494), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT46), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n749), .A2(new_n541), .A3(new_n752), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(new_n559), .ZN(G1329gat));
  INV_X1    g557(.A(new_n713), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n729), .A2(G43gat), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G43gat), .B1(new_n747), .B2(new_n715), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n716), .A3(new_n752), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n760), .B1(new_n765), .B2(G43gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n764), .B(KEYINPUT105), .C1(new_n766), .C2(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1330gat));
  NOR3_X1   g571(.A1(new_n729), .A2(G50gat), .A3(new_n415), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n749), .A2(new_n719), .A3(new_n752), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G50gat), .ZN(new_n775));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n747), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n719), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n775), .A2(KEYINPUT48), .B1(new_n778), .B2(new_n780), .ZN(G1331gat));
  INV_X1    g580(.A(new_n701), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n750), .A2(new_n608), .A3(new_n678), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n703), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT106), .B(G57gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1332gat));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n541), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT49), .B(G64gat), .Z(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(G1333gat));
  AOI21_X1  g589(.A(new_n659), .B1(new_n783), .B2(new_n716), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n759), .A2(G71gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n783), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n783), .A2(new_n719), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g595(.A1(new_n751), .A2(new_n734), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n677), .A2(new_n608), .A3(new_n782), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n471), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n740), .A2(new_n745), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n677), .A2(new_n608), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n727), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n802), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(KEYINPUT107), .A3(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n782), .A2(G85gat), .A3(new_n471), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n800), .B1(new_n810), .B2(new_n811), .ZN(G1336gat));
  NAND3_X1  g611(.A1(new_n805), .A2(KEYINPUT108), .A3(new_n807), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n782), .A2(G92gat), .A3(new_n494), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n803), .A2(new_n815), .A3(new_n804), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n751), .A2(new_n541), .A3(new_n734), .A4(new_n798), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n616), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n808), .A2(new_n809), .A3(new_n814), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n797), .A2(KEYINPUT109), .A3(new_n541), .A4(new_n798), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n818), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n616), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n821), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n821), .A2(new_n828), .A3(new_n823), .A4(new_n822), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n820), .B1(new_n829), .B2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n799), .B2(new_n715), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n713), .A2(new_n614), .A3(new_n701), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n810), .B2(new_n833), .ZN(G1338gat));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n782), .A2(G106gat), .A3(new_n415), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n808), .A2(new_n809), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n751), .A2(new_n719), .A3(new_n734), .A4(new_n798), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n838), .B2(G106gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n813), .A2(new_n816), .A3(new_n836), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(G106gat), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n835), .B(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n840), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT111), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(G1339gat));
  NAND4_X1  g648(.A1(new_n657), .A2(new_n609), .A3(new_n677), .A4(new_n782), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n573), .A2(new_n578), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n852), .A2(new_n575), .B1(new_n587), .B2(new_n589), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n595), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n602), .ZN(new_n857));
  INV_X1    g656(.A(new_n700), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n691), .A2(new_n690), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n680), .A3(new_n688), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n697), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n680), .B1(new_n859), .B2(new_n688), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n692), .A3(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n858), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT55), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n727), .A2(new_n857), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n608), .A2(new_n868), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n701), .A2(new_n602), .A3(new_n856), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n657), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n851), .B1(new_n676), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n719), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n471), .A2(new_n541), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n759), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n204), .B1(new_n882), .B2(new_n608), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n876), .A2(new_n421), .A3(new_n879), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT113), .Z(new_n885));
  NOR2_X1   g684(.A1(new_n609), .A2(G113gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(G1340gat));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n202), .A3(new_n701), .ZN(new_n890));
  OAI21_X1  g689(.A(G120gat), .B1(new_n881), .B2(new_n782), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1341gat));
  NAND3_X1  g691(.A1(new_n882), .A2(G127gat), .A3(new_n677), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  AOI21_X1  g695(.A(G127gat), .B1(new_n884), .B2(new_n677), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1342gat));
  OAI21_X1  g697(.A(G134gat), .B1(new_n881), .B2(new_n657), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT116), .Z(new_n900));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n208), .A3(new_n727), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT56), .Z(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1343gat));
  XNOR2_X1  g702(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n876), .B2(new_n415), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n701), .A2(new_n856), .A3(new_n602), .A4(KEYINPUT118), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n871), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n657), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(KEYINPUT119), .A3(new_n657), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n870), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n851), .B1(new_n914), .B2(new_n676), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n719), .A2(KEYINPUT57), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n905), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n716), .A2(new_n879), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n608), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(G141gat), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n876), .A2(new_n415), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n918), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n923), .A2(G141gat), .A3(new_n609), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n921), .B(new_n924), .C1(KEYINPUT121), .C2(new_n920), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT121), .ZN(new_n926));
  INV_X1    g725(.A(new_n904), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n649), .B(new_n857), .C1(new_n651), .C2(new_n656), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n929), .A2(new_n869), .B1(new_n873), .B2(new_n657), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n850), .B1(new_n930), .B2(new_n677), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n931), .B2(new_n719), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n676), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n850), .ZN(new_n934));
  INV_X1    g733(.A(new_n916), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n918), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT120), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n917), .A2(new_n939), .A3(new_n918), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n940), .A3(new_n608), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n926), .B1(new_n941), .B2(G141gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n925), .B1(new_n942), .B2(new_n920), .ZN(G1344gat));
  INV_X1    g742(.A(new_n923), .ZN(new_n944));
  INV_X1    g743(.A(G148gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n701), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT122), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G148gat), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n917), .A2(new_n939), .A3(new_n918), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n939), .B1(new_n917), .B2(new_n918), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n949), .B1(new_n952), .B2(new_n701), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n719), .A3(new_n927), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n910), .A2(new_n870), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n676), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n415), .B1(new_n956), .B2(new_n850), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n957), .B2(KEYINPUT57), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n937), .A2(new_n782), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n945), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n960), .A2(KEYINPUT123), .A3(new_n948), .ZN(new_n961));
  OAI21_X1  g760(.A(KEYINPUT123), .B1(new_n960), .B2(new_n948), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n947), .B1(new_n953), .B2(new_n963), .ZN(G1345gat));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n672), .A3(new_n677), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n951), .A3(new_n676), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n672), .ZN(G1346gat));
  NOR3_X1   g766(.A1(new_n923), .A2(G162gat), .A3(new_n657), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n950), .A2(new_n951), .A3(new_n657), .ZN(new_n970));
  INV_X1    g769(.A(G162gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G1347gat));
  NAND4_X1  g771(.A1(new_n877), .A2(new_n471), .A3(new_n541), .A4(new_n713), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n973), .A2(new_n247), .A3(new_n609), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n876), .A2(new_n703), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n975), .A2(new_n541), .A3(new_n415), .A4(new_n713), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n608), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n978), .B2(new_n247), .ZN(G1348gat));
  OAI21_X1  g778(.A(G176gat), .B1(new_n973), .B2(new_n782), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n701), .A2(new_n248), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT125), .ZN(G1349gat));
  OAI21_X1  g782(.A(G183gat), .B1(new_n973), .B2(new_n676), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n677), .A2(new_n273), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g786(.A(G190gat), .B1(new_n973), .B2(new_n657), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT61), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n977), .A2(new_n266), .A3(new_n727), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1351gat));
  NOR3_X1   g790(.A1(new_n716), .A2(new_n494), .A3(new_n415), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT126), .ZN(new_n994));
  AOI21_X1  g793(.A(G197gat), .B1(new_n994), .B2(new_n608), .ZN(new_n995));
  AND4_X1   g794(.A1(new_n471), .A2(new_n958), .A3(new_n541), .A4(new_n715), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n608), .A2(G197gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(G1352gat));
  NOR3_X1   g797(.A1(new_n993), .A2(G204gat), .A3(new_n782), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n996), .A2(new_n701), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G204gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1001), .A2(KEYINPUT62), .A3(new_n1002), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(G1353gat));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n360), .A3(new_n677), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n996), .A2(new_n677), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n1011), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1011), .B2(G211gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(G1354gat));
  NAND3_X1  g813(.A1(new_n994), .A2(new_n361), .A3(new_n727), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n727), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1015), .B1(new_n1017), .B2(new_n361), .ZN(G1355gat));
endmodule


