

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787;

  XNOR2_X1 U375 ( .A(n653), .B(n646), .ZN(n778) );
  INV_X1 U376 ( .A(n728), .ZN(n730) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n525) );
  OR2_X1 U378 ( .A1(n578), .A2(n577), .ZN(n728) );
  XNOR2_X1 U379 ( .A(n554), .B(KEYINPUT108), .ZN(n460) );
  AND2_X4 U380 ( .A1(n657), .A2(n400), .ZN(n756) );
  XNOR2_X2 U381 ( .A(n613), .B(KEYINPUT1), .ZN(n560) );
  NOR2_X1 U382 ( .A1(n557), .A2(n673), .ZN(n582) );
  XNOR2_X2 U383 ( .A(n493), .B(KEYINPUT0), .ZN(n572) );
  NAND2_X1 U384 ( .A1(n577), .A2(n578), .ZN(n375) );
  NOR2_X1 U385 ( .A1(n370), .A2(n355), .ZN(n369) );
  AND2_X1 U386 ( .A1(G472), .A2(n533), .ZN(n371) );
  NAND2_X1 U387 ( .A1(n652), .A2(n651), .ZN(n657) );
  NAND2_X1 U388 ( .A1(n401), .A2(n362), .ZN(n400) );
  XNOR2_X1 U389 ( .A(n374), .B(n365), .ZN(n662) );
  NOR2_X1 U390 ( .A1(n639), .A2(n728), .ZN(n374) );
  NOR2_X1 U391 ( .A1(n606), .A2(n605), .ZN(n628) );
  XNOR2_X1 U392 ( .A(n457), .B(n456), .ZN(n614) );
  XNOR2_X1 U393 ( .A(n464), .B(KEYINPUT19), .ZN(n627) );
  NAND2_X2 U394 ( .A1(n369), .A2(n372), .ZN(n679) );
  AND2_X1 U395 ( .A1(n403), .A2(n371), .ZN(n370) );
  XNOR2_X1 U396 ( .A(n532), .B(n481), .ZN(n748) );
  XNOR2_X1 U397 ( .A(n516), .B(n515), .ZN(n771) );
  XNOR2_X1 U398 ( .A(n501), .B(n484), .ZN(n516) );
  XNOR2_X1 U399 ( .A(n463), .B(G113), .ZN(n497) );
  INV_X1 U400 ( .A(G137), .ZN(n514) );
  INV_X1 U401 ( .A(n521), .ZN(n470) );
  NAND2_X1 U402 ( .A1(n423), .A2(n673), .ZN(n422) );
  NAND2_X1 U403 ( .A1(n357), .A2(n458), .ZN(n457) );
  AND2_X1 U404 ( .A1(n613), .A2(n612), .ZN(n458) );
  XNOR2_X1 U405 ( .A(n499), .B(KEYINPUT10), .ZN(n538) );
  NOR2_X1 U406 ( .A1(n603), .A2(n611), .ZN(n618) );
  OR2_X1 U407 ( .A1(n708), .A2(G902), .ZN(n469) );
  OR2_X1 U408 ( .A1(n403), .A2(G472), .ZN(n372) );
  INV_X2 U409 ( .A(G953), .ZN(n780) );
  NAND2_X1 U410 ( .A1(n476), .A2(KEYINPUT71), .ZN(n475) );
  INV_X1 U411 ( .A(KEYINPUT47), .ZN(n476) );
  AND2_X1 U412 ( .A1(n454), .A2(n455), .ZN(n448) );
  NOR2_X1 U413 ( .A1(n783), .A2(n662), .ZN(n447) );
  NAND2_X1 U414 ( .A1(n390), .A2(KEYINPUT88), .ZN(n389) );
  AND2_X1 U415 ( .A1(n460), .A2(n408), .ZN(n590) );
  INV_X1 U416 ( .A(KEYINPUT72), .ZN(n456) );
  XNOR2_X1 U417 ( .A(n380), .B(KEYINPUT9), .ZN(n379) );
  INV_X1 U418 ( .A(KEYINPUT101), .ZN(n380) );
  XNOR2_X1 U419 ( .A(G116), .B(KEYINPUT102), .ZN(n377) );
  NAND2_X1 U420 ( .A1(n690), .A2(n617), .ZN(n387) );
  NAND2_X1 U421 ( .A1(n634), .A2(n415), .ZN(n414) );
  XNOR2_X1 U422 ( .A(n642), .B(n598), .ZN(n689) );
  XNOR2_X1 U423 ( .A(n485), .B(n480), .ZN(n597) );
  INV_X1 U424 ( .A(KEYINPUT28), .ZN(n467) );
  NAND2_X1 U425 ( .A1(n604), .A2(n618), .ZN(n468) );
  NAND2_X2 U426 ( .A1(n394), .A2(n391), .ZN(n613) );
  AND2_X1 U427 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U428 ( .A1(n393), .A2(n533), .ZN(n392) );
  XNOR2_X1 U429 ( .A(n532), .B(n531), .ZN(n403) );
  XNOR2_X1 U430 ( .A(G140), .B(G128), .ZN(n546) );
  XOR2_X1 U431 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n504) );
  XNOR2_X1 U432 ( .A(n381), .B(n772), .ZN(n708) );
  XNOR2_X1 U433 ( .A(n382), .B(n385), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n383), .B(n497), .ZN(n382) );
  XNOR2_X1 U435 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n484) );
  XNOR2_X1 U436 ( .A(n499), .B(n517), .ZN(n407) );
  NAND2_X1 U437 ( .A1(n412), .A2(n409), .ZN(n639) );
  AND2_X1 U438 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U439 ( .A1(n411), .A2(n410), .ZN(n409) );
  NAND2_X1 U440 ( .A1(n689), .A2(n415), .ZN(n413) );
  BUF_X1 U441 ( .A(n560), .Z(n673) );
  INV_X1 U442 ( .A(KEYINPUT75), .ZN(n421) );
  OR2_X1 U443 ( .A1(n758), .A2(G902), .ZN(n465) );
  XNOR2_X1 U444 ( .A(n575), .B(n574), .ZN(n577) );
  XNOR2_X1 U445 ( .A(n679), .B(n555), .ZN(n620) );
  XNOR2_X1 U446 ( .A(n404), .B(n439), .ZN(n441) );
  XNOR2_X1 U447 ( .A(n500), .B(n497), .ZN(n439) );
  XNOR2_X1 U448 ( .A(n527), .B(n440), .ZN(n404) );
  XNOR2_X1 U449 ( .A(n462), .B(KEYINPUT16), .ZN(n440) );
  NOR2_X1 U450 ( .A1(n354), .A2(n429), .ZN(n420) );
  NAND2_X1 U451 ( .A1(n359), .A2(KEYINPUT119), .ZN(n418) );
  NOR2_X1 U452 ( .A1(n428), .A2(G953), .ZN(n427) );
  NOR2_X1 U453 ( .A1(n400), .A2(n429), .ZN(n428) );
  NOR2_X1 U454 ( .A1(n629), .A2(n785), .ZN(n455) );
  NAND2_X1 U455 ( .A1(n435), .A2(n636), .ZN(n637) );
  XNOR2_X1 U456 ( .A(n436), .B(KEYINPUT77), .ZN(n435) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n488) );
  OR2_X1 U458 ( .A1(G902), .A2(G237), .ZN(n486) );
  NAND2_X1 U459 ( .A1(n748), .A2(n524), .ZN(n396) );
  XOR2_X1 U460 ( .A(KEYINPUT5), .B(G113), .Z(n526) );
  XNOR2_X1 U461 ( .A(n433), .B(n384), .ZN(n383) );
  INV_X1 U462 ( .A(KEYINPUT99), .ZN(n384) );
  XNOR2_X1 U463 ( .A(KEYINPUT11), .B(G143), .ZN(n433) );
  XNOR2_X1 U464 ( .A(n434), .B(G122), .ZN(n432) );
  INV_X1 U465 ( .A(KEYINPUT12), .ZN(n434) );
  XNOR2_X1 U466 ( .A(G902), .B(KEYINPUT15), .ZN(n649) );
  INV_X1 U467 ( .A(KEYINPUT39), .ZN(n415) );
  NOR2_X1 U468 ( .A1(n689), .A2(n415), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n373), .B(n610), .ZN(n615) );
  INV_X1 U470 ( .A(G104), .ZN(n463) );
  INV_X1 U471 ( .A(G110), .ZN(n462) );
  XNOR2_X1 U472 ( .A(n461), .B(G119), .ZN(n527) );
  XNOR2_X1 U473 ( .A(G116), .B(KEYINPUT3), .ZN(n461) );
  XNOR2_X1 U474 ( .A(n378), .B(n376), .ZN(n506) );
  XNOR2_X1 U475 ( .A(n502), .B(n377), .ZN(n376) );
  XNOR2_X1 U476 ( .A(KEYINPUT7), .B(KEYINPUT103), .ZN(n502) );
  XOR2_X1 U477 ( .A(G107), .B(G122), .Z(n500) );
  XNOR2_X1 U478 ( .A(G140), .B(G131), .ZN(n521) );
  XNOR2_X1 U479 ( .A(G110), .B(G107), .ZN(n520) );
  OR2_X1 U480 ( .A1(n451), .A2(n449), .ZN(n687) );
  NAND2_X1 U481 ( .A1(n387), .A2(n356), .ZN(n386) );
  NAND2_X1 U482 ( .A1(n597), .A2(n617), .ZN(n464) );
  XNOR2_X1 U483 ( .A(n468), .B(n466), .ZN(n606) );
  XNOR2_X1 U484 ( .A(n467), .B(KEYINPUT109), .ZN(n466) );
  INV_X1 U485 ( .A(KEYINPUT62), .ZN(n402) );
  XNOR2_X1 U486 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U487 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U488 ( .A(n405), .B(n441), .ZN(n741) );
  XNOR2_X1 U489 ( .A(n353), .B(n406), .ZN(n405) );
  INV_X1 U490 ( .A(KEYINPUT35), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n558), .B(n459), .ZN(n408) );
  XNOR2_X1 U492 ( .A(n422), .B(n421), .ZN(n556) );
  NAND2_X1 U493 ( .A1(n582), .A2(n553), .ZN(n554) );
  NAND2_X1 U494 ( .A1(n443), .A2(n675), .ZN(n714) );
  XNOR2_X1 U495 ( .A(n583), .B(n444), .ZN(n443) );
  INV_X1 U496 ( .A(KEYINPUT86), .ZN(n444) );
  NAND2_X1 U497 ( .A1(n419), .A2(n417), .ZN(n705) );
  NAND2_X1 U498 ( .A1(n363), .A2(n430), .ZN(n419) );
  AND2_X1 U499 ( .A1(n416), .A2(n418), .ZN(n417) );
  XOR2_X1 U500 ( .A(n483), .B(n364), .Z(n353) );
  NAND2_X1 U501 ( .A1(n704), .A2(n703), .ZN(n354) );
  AND2_X1 U502 ( .A1(G902), .A2(n534), .ZN(n355) );
  XOR2_X1 U503 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n356) );
  NOR2_X2 U504 ( .A1(n602), .A2(n559), .ZN(n357) );
  XOR2_X1 U505 ( .A(KEYINPUT13), .B(G475), .Z(n358) );
  NAND2_X1 U506 ( .A1(n614), .A2(n615), .ZN(n634) );
  AND2_X1 U507 ( .A1(n702), .A2(n700), .ZN(n359) );
  NOR2_X1 U508 ( .A1(n689), .A2(n688), .ZN(n360) );
  OR2_X1 U509 ( .A1(n453), .A2(n450), .ZN(n361) );
  AND2_X1 U510 ( .A1(n655), .A2(KEYINPUT2), .ZN(n362) );
  AND2_X1 U511 ( .A1(n427), .A2(KEYINPUT119), .ZN(n363) );
  INV_X1 U512 ( .A(n690), .ZN(n453) );
  AND2_X1 U513 ( .A1(G224), .A2(n780), .ZN(n364) );
  XOR2_X1 U514 ( .A(n616), .B(KEYINPUT40), .Z(n365) );
  XOR2_X1 U515 ( .A(n565), .B(KEYINPUT34), .Z(n366) );
  AND2_X1 U516 ( .A1(n477), .A2(KEYINPUT47), .ZN(n367) );
  XOR2_X1 U517 ( .A(n403), .B(n402), .Z(n368) );
  OR2_X1 U518 ( .A1(n688), .A2(n356), .ZN(n450) );
  OR2_X1 U519 ( .A1(n679), .A2(n688), .ZN(n373) );
  INV_X1 U520 ( .A(n688), .ZN(n617) );
  XNOR2_X2 U521 ( .A(n375), .B(n576), .ZN(n733) );
  XNOR2_X2 U522 ( .A(n469), .B(n358), .ZN(n575) );
  XNOR2_X1 U523 ( .A(n501), .B(n379), .ZN(n378) );
  XNOR2_X2 U524 ( .A(G143), .B(G128), .ZN(n501) );
  XNOR2_X1 U525 ( .A(n432), .B(n498), .ZN(n385) );
  NAND2_X1 U526 ( .A1(n452), .A2(n386), .ZN(n451) );
  NAND2_X1 U527 ( .A1(n388), .A2(KEYINPUT44), .ZN(n588) );
  NAND2_X1 U528 ( .A1(n590), .A2(n389), .ZN(n388) );
  INV_X1 U529 ( .A(n424), .ZN(n390) );
  XNOR2_X2 U530 ( .A(n397), .B(n425), .ZN(n424) );
  OR2_X1 U531 ( .A1(n748), .A2(n392), .ZN(n391) );
  INV_X1 U532 ( .A(n524), .ZN(n393) );
  NAND2_X1 U533 ( .A1(n524), .A2(G902), .ZN(n395) );
  NAND2_X1 U534 ( .A1(n398), .A2(n632), .ZN(n397) );
  XNOR2_X1 U535 ( .A(n399), .B(n366), .ZN(n398) );
  NOR2_X1 U536 ( .A1(n671), .A2(n572), .ZN(n399) );
  NAND2_X1 U537 ( .A1(n670), .A2(n400), .ZN(n426) );
  INV_X1 U538 ( .A(n656), .ZN(n401) );
  XNOR2_X1 U539 ( .A(n407), .B(n516), .ZN(n406) );
  XNOR2_X1 U540 ( .A(n408), .B(G119), .ZN(G21) );
  INV_X1 U541 ( .A(n634), .ZN(n411) );
  NAND2_X1 U542 ( .A1(n426), .A2(n420), .ZN(n416) );
  AND2_X1 U543 ( .A1(n620), .A2(n602), .ZN(n423) );
  NAND2_X1 U544 ( .A1(n424), .A2(n591), .ZN(n592) );
  NOR2_X1 U545 ( .A1(n424), .A2(n591), .ZN(n585) );
  XNOR2_X1 U546 ( .A(n424), .B(G122), .ZN(G24) );
  INV_X1 U547 ( .A(n672), .ZN(n429) );
  NAND2_X1 U548 ( .A1(n431), .A2(n672), .ZN(n430) );
  INV_X1 U549 ( .A(n670), .ZN(n431) );
  NAND2_X1 U550 ( .A1(n437), .A2(n726), .ZN(n436) );
  NAND2_X1 U551 ( .A1(n631), .A2(KEYINPUT47), .ZN(n437) );
  XNOR2_X2 U552 ( .A(n438), .B(KEYINPUT105), .ZN(n692) );
  NOR2_X2 U553 ( .A1(n733), .A2(n730), .ZN(n438) );
  XNOR2_X1 U554 ( .A(n441), .B(G101), .ZN(n767) );
  XNOR2_X1 U555 ( .A(n551), .B(n550), .ZN(n758) );
  NAND2_X1 U556 ( .A1(n442), .A2(n588), .ZN(n589) );
  NOR2_X1 U557 ( .A1(n587), .A2(n586), .ZN(n442) );
  XNOR2_X1 U558 ( .A(n445), .B(n638), .ZN(n645) );
  NAND2_X1 U559 ( .A1(n448), .A2(n446), .ZN(n445) );
  XNOR2_X1 U560 ( .A(n447), .B(KEYINPUT46), .ZN(n446) );
  NAND2_X1 U561 ( .A1(n689), .A2(n356), .ZN(n452) );
  NOR2_X1 U562 ( .A1(n689), .A2(n361), .ZN(n449) );
  XNOR2_X1 U563 ( .A(n637), .B(KEYINPUT79), .ZN(n454) );
  XNOR2_X2 U564 ( .A(n465), .B(n552), .ZN(n602) );
  XNOR2_X2 U565 ( .A(n771), .B(n518), .ZN(n532) );
  INV_X1 U566 ( .A(KEYINPUT32), .ZN(n459) );
  XNOR2_X1 U567 ( .A(n460), .B(G110), .ZN(G12) );
  XNOR2_X2 U568 ( .A(G146), .B(G125), .ZN(n499) );
  INV_X1 U569 ( .A(n761), .ZN(n656) );
  NAND2_X1 U570 ( .A1(n647), .A2(n761), .ZN(n648) );
  XNOR2_X2 U571 ( .A(n596), .B(KEYINPUT45), .ZN(n761) );
  NAND2_X1 U572 ( .A1(n656), .A2(n663), .ZN(n666) );
  NAND2_X1 U573 ( .A1(n627), .A2(n492), .ZN(n493) );
  XNOR2_X1 U574 ( .A(n538), .B(n470), .ZN(n772) );
  NOR2_X1 U575 ( .A1(n727), .A2(n367), .ZN(n473) );
  NOR2_X1 U576 ( .A1(n474), .A2(n471), .ZN(n629) );
  NAND2_X1 U577 ( .A1(n473), .A2(n472), .ZN(n471) );
  NAND2_X1 U578 ( .A1(n626), .A2(n477), .ZN(n472) );
  NOR2_X1 U579 ( .A1(n626), .A2(n475), .ZN(n474) );
  INV_X1 U580 ( .A(KEYINPUT71), .ZN(n477) );
  XNOR2_X1 U581 ( .A(n692), .B(KEYINPUT81), .ZN(n626) );
  XNOR2_X1 U582 ( .A(n478), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U583 ( .A1(n479), .A2(n660), .ZN(n478) );
  XNOR2_X1 U584 ( .A(n658), .B(n368), .ZN(n479) );
  XNOR2_X1 U585 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U586 ( .A(n665), .B(n664), .ZN(n667) );
  AND2_X1 U587 ( .A1(G210), .A2(n486), .ZN(n480) );
  XOR2_X1 U588 ( .A(n523), .B(n522), .Z(n481) );
  XNOR2_X1 U589 ( .A(n526), .B(G131), .ZN(n528) );
  XNOR2_X1 U590 ( .A(n527), .B(n528), .ZN(n529) );
  INV_X1 U591 ( .A(n611), .ZN(n612) );
  INV_X1 U592 ( .A(KEYINPUT95), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n567), .B(KEYINPUT97), .ZN(n568) );
  INV_X1 U594 ( .A(n760), .ZN(n660) );
  XNOR2_X1 U595 ( .A(n569), .B(n568), .ZN(n734) );
  XNOR2_X1 U596 ( .A(KEYINPUT91), .B(KEYINPUT17), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n482), .B(KEYINPUT18), .ZN(n483) );
  XNOR2_X1 U598 ( .A(KEYINPUT67), .B(G101), .ZN(n517) );
  NAND2_X1 U599 ( .A1(n741), .A2(n649), .ZN(n485) );
  NAND2_X1 U600 ( .A1(G214), .A2(n486), .ZN(n487) );
  XOR2_X1 U601 ( .A(KEYINPUT92), .B(n487), .Z(n688) );
  XNOR2_X1 U602 ( .A(n488), .B(KEYINPUT14), .ZN(n489) );
  AND2_X1 U603 ( .A1(n489), .A2(G952), .ZN(n701) );
  AND2_X1 U604 ( .A1(n701), .A2(n780), .ZN(n700) );
  NAND2_X1 U605 ( .A1(G902), .A2(n489), .ZN(n599) );
  OR2_X1 U606 ( .A1(n780), .A2(G898), .ZN(n768) );
  NOR2_X1 U607 ( .A1(n599), .A2(n768), .ZN(n490) );
  NOR2_X1 U608 ( .A1(n700), .A2(n490), .ZN(n491) );
  XNOR2_X1 U609 ( .A(KEYINPUT93), .B(n491), .ZN(n492) );
  NAND2_X1 U610 ( .A1(n649), .A2(G234), .ZN(n494) );
  XNOR2_X1 U611 ( .A(n494), .B(KEYINPUT20), .ZN(n535) );
  NAND2_X1 U612 ( .A1(n535), .A2(G221), .ZN(n496) );
  XOR2_X1 U613 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n495) );
  XNOR2_X1 U614 ( .A(n496), .B(n495), .ZN(n676) );
  NAND2_X1 U615 ( .A1(n525), .A2(G214), .ZN(n498) );
  XNOR2_X1 U616 ( .A(G134), .B(n500), .ZN(n508) );
  NAND2_X1 U617 ( .A1(G234), .A2(n780), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n504), .B(n503), .ZN(n545) );
  NAND2_X1 U619 ( .A1(G217), .A2(n545), .ZN(n505) );
  XNOR2_X1 U620 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U621 ( .A(n508), .B(n507), .ZN(n752) );
  NOR2_X1 U622 ( .A1(G902), .A2(n752), .ZN(n510) );
  INV_X1 U623 ( .A(G478), .ZN(n509) );
  XNOR2_X1 U624 ( .A(n510), .B(n509), .ZN(n578) );
  NOR2_X1 U625 ( .A1(n575), .A2(n578), .ZN(n690) );
  NAND2_X1 U626 ( .A1(n676), .A2(n690), .ZN(n511) );
  NOR2_X1 U627 ( .A1(n572), .A2(n511), .ZN(n513) );
  XNOR2_X1 U628 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n512) );
  XNOR2_X1 U629 ( .A(n513), .B(n512), .ZN(n557) );
  XNOR2_X1 U630 ( .A(n514), .B(G134), .ZN(n515) );
  XNOR2_X1 U631 ( .A(n517), .B(G146), .ZN(n518) );
  NAND2_X1 U632 ( .A1(n780), .A2(G227), .ZN(n519) );
  XNOR2_X1 U633 ( .A(n519), .B(G104), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U635 ( .A(KEYINPUT70), .B(G469), .ZN(n524) );
  NAND2_X1 U636 ( .A1(n525), .A2(G210), .ZN(n530) );
  XNOR2_X1 U637 ( .A(n530), .B(n529), .ZN(n531) );
  INV_X1 U638 ( .A(G902), .ZN(n533) );
  INV_X1 U639 ( .A(G472), .ZN(n534) );
  XOR2_X1 U640 ( .A(KEYINPUT73), .B(KEYINPUT25), .Z(n537) );
  NAND2_X1 U641 ( .A1(n535), .A2(G217), .ZN(n536) );
  XNOR2_X1 U642 ( .A(n537), .B(n536), .ZN(n552) );
  XNOR2_X1 U643 ( .A(n538), .B(KEYINPUT24), .ZN(n544) );
  XOR2_X1 U644 ( .A(KEYINPUT94), .B(KEYINPUT82), .Z(n540) );
  XNOR2_X1 U645 ( .A(G137), .B(KEYINPUT23), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n540), .B(n539), .ZN(n542) );
  XNOR2_X1 U647 ( .A(n544), .B(n543), .ZN(n551) );
  NAND2_X1 U648 ( .A1(G221), .A2(n545), .ZN(n549) );
  XOR2_X1 U649 ( .A(G119), .B(G110), .Z(n547) );
  XNOR2_X1 U650 ( .A(n547), .B(n546), .ZN(n548) );
  AND2_X1 U651 ( .A1(n679), .A2(n602), .ZN(n553) );
  INV_X1 U652 ( .A(n602), .ZN(n675) );
  XNOR2_X1 U653 ( .A(KEYINPUT107), .B(KEYINPUT6), .ZN(n555) );
  NOR2_X1 U654 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U655 ( .A(n676), .ZN(n559) );
  NAND2_X1 U656 ( .A1(n560), .A2(n357), .ZN(n566) );
  INV_X1 U657 ( .A(n566), .ZN(n562) );
  INV_X1 U658 ( .A(n620), .ZN(n561) );
  NAND2_X1 U659 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U660 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n563) );
  XNOR2_X1 U661 ( .A(n564), .B(n563), .ZN(n671) );
  INV_X1 U662 ( .A(KEYINPUT74), .ZN(n565) );
  AND2_X1 U663 ( .A1(n578), .A2(n575), .ZN(n632) );
  OR2_X1 U664 ( .A1(n566), .A2(n679), .ZN(n682) );
  NOR2_X1 U665 ( .A1(n572), .A2(n682), .ZN(n569) );
  XNOR2_X1 U666 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n567) );
  INV_X1 U667 ( .A(n734), .ZN(n573) );
  AND2_X1 U668 ( .A1(n613), .A2(n357), .ZN(n570) );
  NAND2_X1 U669 ( .A1(n570), .A2(n679), .ZN(n571) );
  OR2_X1 U670 ( .A1(n572), .A2(n571), .ZN(n715) );
  NAND2_X1 U671 ( .A1(n573), .A2(n715), .ZN(n580) );
  INV_X1 U672 ( .A(KEYINPUT100), .ZN(n574) );
  INV_X1 U673 ( .A(KEYINPUT104), .ZN(n576) );
  INV_X1 U674 ( .A(n626), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U676 ( .A(n581), .B(KEYINPUT106), .ZN(n584) );
  NAND2_X1 U677 ( .A1(n582), .A2(n620), .ZN(n583) );
  NAND2_X1 U678 ( .A1(n584), .A2(n714), .ZN(n587) );
  NOR2_X1 U679 ( .A1(n585), .A2(KEYINPUT88), .ZN(n586) );
  XNOR2_X1 U680 ( .A(n589), .B(KEYINPUT87), .ZN(n595) );
  INV_X1 U681 ( .A(n590), .ZN(n593) );
  INV_X1 U682 ( .A(KEYINPUT44), .ZN(n591) );
  OR2_X1 U683 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U684 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U685 ( .A(n597), .ZN(n642) );
  INV_X1 U686 ( .A(KEYINPUT38), .ZN(n598) );
  OR2_X1 U687 ( .A1(n780), .A2(n599), .ZN(n600) );
  NOR2_X1 U688 ( .A1(n600), .A2(G900), .ZN(n601) );
  NOR2_X1 U689 ( .A1(n700), .A2(n601), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n602), .A2(n676), .ZN(n603) );
  INV_X1 U691 ( .A(n679), .ZN(n604) );
  INV_X1 U692 ( .A(n613), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n687), .A2(n628), .ZN(n609) );
  INV_X1 U694 ( .A(KEYINPUT112), .ZN(n607) );
  XNOR2_X1 U695 ( .A(n607), .B(KEYINPUT42), .ZN(n608) );
  XNOR2_X1 U696 ( .A(n609), .B(n608), .ZN(n783) );
  INV_X1 U697 ( .A(KEYINPUT30), .ZN(n610) );
  INV_X1 U698 ( .A(KEYINPUT110), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n621), .A2(n730), .ZN(n640) );
  NOR2_X1 U702 ( .A1(n642), .A2(n640), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT36), .B(n622), .ZN(n623) );
  AND2_X1 U704 ( .A1(n623), .A2(n673), .ZN(n625) );
  INV_X1 U705 ( .A(KEYINPUT113), .ZN(n624) );
  XNOR2_X1 U706 ( .A(n625), .B(n624), .ZN(n785) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n727) );
  NAND2_X1 U708 ( .A1(KEYINPUT47), .A2(n727), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT80), .ZN(n636) );
  INV_X1 U710 ( .A(n692), .ZN(n631) );
  INV_X1 U711 ( .A(n632), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n642), .A2(n633), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n635), .A2(n411), .ZN(n726) );
  XNOR2_X1 U714 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n638) );
  INV_X1 U715 ( .A(n733), .ZN(n723) );
  OR2_X1 U716 ( .A1(n639), .A2(n723), .ZN(n661) );
  OR2_X1 U717 ( .A1(n640), .A2(n673), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n641), .B(KEYINPUT43), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n737) );
  AND2_X1 U720 ( .A1(n661), .A2(n737), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n653) );
  INV_X1 U722 ( .A(KEYINPUT85), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n778), .A2(n649), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n648), .B(KEYINPUT84), .ZN(n652) );
  INV_X1 U725 ( .A(n649), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n650), .A2(KEYINPUT2), .ZN(n651) );
  BUF_X1 U727 ( .A(n653), .Z(n654) );
  INV_X1 U728 ( .A(n654), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n756), .A2(G472), .ZN(n658) );
  INV_X1 U730 ( .A(G952), .ZN(n659) );
  AND2_X1 U731 ( .A1(n659), .A2(G953), .ZN(n760) );
  XNOR2_X1 U732 ( .A(n661), .B(G134), .ZN(G36) );
  XOR2_X1 U733 ( .A(G131), .B(n662), .Z(G33) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n778), .A2(n663), .ZN(n665) );
  INV_X1 U736 ( .A(KEYINPUT83), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n669) );
  INV_X1 U738 ( .A(KEYINPUT76), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(n670) );
  INV_X1 U740 ( .A(n671), .ZN(n695) );
  NAND2_X1 U741 ( .A1(n687), .A2(n695), .ZN(n672) );
  NOR2_X1 U742 ( .A1(n673), .A2(n357), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(KEYINPUT50), .ZN(n681) );
  NOR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(KEYINPUT49), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n684) );
  INV_X1 U748 ( .A(n682), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(KEYINPUT51), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n698) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U754 ( .A1(n360), .A2(n692), .ZN(n693) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U758 ( .A(n699), .B(KEYINPUT52), .ZN(n702) );
  NAND2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U760 ( .A1(G953), .A2(KEYINPUT119), .ZN(n703) );
  XNOR2_X1 U761 ( .A(n705), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U762 ( .A1(n756), .A2(G475), .ZN(n710) );
  XOR2_X1 U763 ( .A(KEYINPUT66), .B(KEYINPUT90), .Z(n706) );
  XNOR2_X1 U764 ( .A(n706), .B(KEYINPUT59), .ZN(n707) );
  XNOR2_X1 U765 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X2 U766 ( .A1(n711), .A2(n760), .ZN(n713) );
  XNOR2_X1 U767 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n713), .B(n712), .ZN(G60) );
  XNOR2_X1 U769 ( .A(n714), .B(G101), .ZN(G3) );
  INV_X1 U770 ( .A(n715), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n720), .A2(n730), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n716), .B(G104), .ZN(G6) );
  XOR2_X1 U773 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n718) );
  XNOR2_X1 U774 ( .A(G107), .B(KEYINPUT114), .ZN(n717) );
  XNOR2_X1 U775 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U776 ( .A(KEYINPUT26), .B(n719), .Z(n722) );
  NAND2_X1 U777 ( .A1(n720), .A2(n733), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n722), .B(n721), .ZN(G9) );
  NOR2_X1 U779 ( .A1(n723), .A2(n727), .ZN(n725) );
  XNOR2_X1 U780 ( .A(G128), .B(KEYINPUT29), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n725), .B(n724), .ZN(G30) );
  XNOR2_X1 U782 ( .A(G143), .B(n726), .ZN(G45) );
  NOR2_X1 U783 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U784 ( .A(G146), .B(n729), .Z(G48) );
  NAND2_X1 U785 ( .A1(n734), .A2(n730), .ZN(n731) );
  XNOR2_X1 U786 ( .A(n731), .B(KEYINPUT116), .ZN(n732) );
  XNOR2_X1 U787 ( .A(G113), .B(n732), .ZN(G15) );
  XOR2_X1 U788 ( .A(G116), .B(KEYINPUT117), .Z(n736) );
  NAND2_X1 U789 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U790 ( .A(n736), .B(n735), .ZN(G18) );
  XNOR2_X1 U791 ( .A(G140), .B(n737), .ZN(G42) );
  NAND2_X1 U792 ( .A1(n756), .A2(G210), .ZN(n743) );
  XOR2_X1 U793 ( .A(KEYINPUT78), .B(KEYINPUT55), .Z(n739) );
  XNOR2_X1 U794 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n738) );
  XNOR2_X1 U795 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U796 ( .A(n741), .B(n740), .Z(n742) );
  XNOR2_X1 U797 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X2 U798 ( .A1(n744), .A2(n760), .ZN(n745) );
  XNOR2_X1 U799 ( .A(n745), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U800 ( .A1(n756), .A2(G469), .ZN(n750) );
  XNOR2_X1 U801 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n746) );
  XNOR2_X1 U802 ( .A(n746), .B(KEYINPUT57), .ZN(n747) );
  XNOR2_X1 U803 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U804 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n760), .A2(n751), .ZN(G54) );
  NAND2_X1 U806 ( .A1(n756), .A2(G478), .ZN(n754) );
  XOR2_X1 U807 ( .A(n752), .B(KEYINPUT123), .Z(n753) );
  XNOR2_X1 U808 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U809 ( .A1(n760), .A2(n755), .ZN(G63) );
  NAND2_X1 U810 ( .A1(n756), .A2(G217), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U812 ( .A1(n760), .A2(n759), .ZN(G66) );
  NAND2_X1 U813 ( .A1(n761), .A2(n780), .ZN(n765) );
  NAND2_X1 U814 ( .A1(G953), .A2(G224), .ZN(n762) );
  XNOR2_X1 U815 ( .A(KEYINPUT61), .B(n762), .ZN(n763) );
  NAND2_X1 U816 ( .A1(n763), .A2(G898), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n766), .B(KEYINPUT124), .ZN(n770) );
  NAND2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U820 ( .A(n770), .B(n769), .Z(G69) );
  XNOR2_X1 U821 ( .A(G227), .B(KEYINPUT126), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n772), .B(n771), .ZN(n776) );
  XOR2_X1 U823 ( .A(n773), .B(n776), .Z(n774) );
  NAND2_X1 U824 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U825 ( .A1(n775), .A2(G953), .ZN(n782) );
  XNOR2_X1 U826 ( .A(n776), .B(KEYINPUT125), .ZN(n777) );
  XNOR2_X1 U827 ( .A(n778), .B(n777), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n782), .A2(n781), .ZN(G72) );
  XNOR2_X1 U830 ( .A(G137), .B(n783), .ZN(n784) );
  XNOR2_X1 U831 ( .A(n784), .B(KEYINPUT127), .ZN(G39) );
  XNOR2_X1 U832 ( .A(n785), .B(KEYINPUT118), .ZN(n786) );
  XNOR2_X1 U833 ( .A(n786), .B(KEYINPUT37), .ZN(n787) );
  XNOR2_X1 U834 ( .A(G125), .B(n787), .ZN(G27) );
endmodule

