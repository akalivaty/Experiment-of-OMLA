//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT28), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT72), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT27), .B1(new_n206), .B2(KEYINPUT70), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G183gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n207), .B(new_n203), .C1(KEYINPUT70), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT71), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n210), .A2(KEYINPUT71), .A3(new_n211), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n216), .A2(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n220), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT73), .B1(new_n222), .B2(KEYINPUT26), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n224), .A3(new_n219), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n206), .A2(new_n203), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n214), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT64), .B1(new_n220), .B2(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n231), .B(new_n232), .C1(G169gat), .C2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n215), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n235), .A2(new_n236), .B1(KEYINPUT23), .B2(new_n220), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n206), .A2(new_n203), .A3(KEYINPUT24), .ZN(new_n240));
  XOR2_X1   g039(.A(G183gat), .B(G190gat), .Z(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(KEYINPUT24), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n234), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n216), .B2(new_n218), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n203), .A2(G183gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n206), .A2(G190gat), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n240), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT67), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n250), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n234), .A2(KEYINPUT25), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n248), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n230), .B2(new_n233), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT67), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT67), .B1(new_n235), .B2(new_n236), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n261), .A2(new_n264), .A3(KEYINPUT68), .A4(new_n242), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n247), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n247), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n229), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT75), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(new_n229), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n271), .A2(KEYINPUT78), .A3(new_n273), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n247), .A2(new_n266), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n229), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n275), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n266), .A2(new_n247), .B1(new_n214), .B2(new_n228), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n274), .C1(new_n287), .C2(KEYINPUT29), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G197gat), .B(G204gat), .Z(new_n291));
  NAND2_X1  g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT22), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(G211gat), .A2(G218gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n295), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n271), .A2(new_n283), .A3(new_n273), .A4(new_n274), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n275), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n304), .A2(KEYINPUT76), .A3(new_n299), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n280), .A2(KEYINPUT79), .A3(new_n300), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n312), .B(new_n313), .Z(new_n314));
  NAND4_X1  g113(.A1(new_n303), .A2(new_n310), .A3(new_n311), .A4(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n314), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(new_n316), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n310), .A3(new_n311), .A4(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n310), .A3(new_n311), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n314), .B(KEYINPUT80), .Z(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n317), .A2(new_n323), .A3(KEYINPUT89), .A4(new_n320), .ZN(new_n327));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT0), .ZN(new_n329));
  XNOR2_X1  g128(.A(G57gat), .B(G85gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G141gat), .B(G148gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(KEYINPUT2), .ZN(new_n336));
  XOR2_X1   g135(.A(G113gat), .B(G120gat), .Z(new_n337));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G155gat), .ZN(new_n342));
  INV_X1    g141(.A(G162gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT2), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT82), .ZN(new_n345));
  INV_X1    g144(.A(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G141gat), .ZN(new_n347));
  XOR2_X1   g146(.A(KEYINPUT81), .B(G141gat), .Z(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n349), .A3(new_n333), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n336), .B(new_n341), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n336), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n350), .A2(new_n351), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n341), .B(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n355), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT5), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT85), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n355), .A2(new_n366), .A3(KEYINPUT4), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n368), .A3(new_n341), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n355), .B2(KEYINPUT4), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n336), .B1(new_n353), .B2(new_n354), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n360), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n363), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n365), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n378));
  INV_X1    g177(.A(new_n375), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n341), .B(KEYINPUT84), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n358), .B2(new_n374), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n378), .B(new_n362), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n355), .A2(KEYINPUT4), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT86), .B1(new_n355), .B2(KEYINPUT4), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n358), .A2(new_n387), .A3(new_n368), .A4(new_n341), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n382), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n332), .B1(new_n377), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n383), .A2(new_n384), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT87), .B1(new_n355), .B2(KEYINPUT4), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n386), .B(new_n388), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n375), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n362), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT39), .B1(new_n361), .B2(new_n363), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT39), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n332), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n391), .B1(new_n401), .B2(KEYINPUT40), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(KEYINPUT40), .B2(new_n401), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n326), .A2(new_n327), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT31), .B(G50gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n298), .B1(new_n375), .B2(new_n283), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n298), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n297), .B1(new_n291), .B2(new_n294), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n283), .B1(new_n411), .B2(KEYINPUT88), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n374), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n413), .A2(new_n372), .B1(G228gat), .B2(G233gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT3), .B1(new_n298), .B2(new_n283), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n358), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(G228gat), .B(G233gat), .C1(new_n407), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n406), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G22gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n418), .A3(new_n406), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n422), .ZN(new_n425));
  INV_X1    g224(.A(new_n423), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(new_n419), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n367), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n370), .A2(new_n369), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n376), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT5), .A3(new_n364), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n394), .A2(new_n378), .A3(new_n376), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n331), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n391), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(KEYINPUT6), .B(new_n332), .C1(new_n377), .C2(new_n390), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n315), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n280), .A2(KEYINPUT79), .A3(new_n300), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT79), .B1(new_n280), .B2(new_n300), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n310), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n298), .B(new_n290), .C1(new_n278), .C2(new_n279), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n304), .A2(new_n298), .A3(new_n305), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT37), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n445), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n290), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n280), .A2(new_n299), .A3(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(KEYINPUT90), .A3(KEYINPUT37), .A4(new_n447), .ZN(new_n452));
  INV_X1    g251(.A(new_n322), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT38), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n439), .B1(new_n444), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n318), .B1(new_n321), .B2(KEYINPUT37), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n443), .B1(new_n442), .B2(new_n310), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n428), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n404), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n436), .A2(new_n437), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n317), .A2(new_n323), .A3(new_n462), .A4(new_n320), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n428), .ZN(new_n464));
  INV_X1    g263(.A(new_n341), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n270), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n341), .B(new_n229), .C1(new_n268), .C2(new_n269), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G227gat), .ZN(new_n469));
  INV_X1    g268(.A(G233gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT32), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(G71gat), .B(G99gat), .Z(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G43gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n466), .B2(new_n467), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n473), .B(new_n476), .C1(KEYINPUT33), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(KEYINPUT33), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT74), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT74), .ZN(new_n483));
  INV_X1    g282(.A(new_n481), .ZN(new_n484));
  NOR4_X1   g283(.A1(new_n477), .A2(new_n483), .A3(new_n479), .A4(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n478), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n472), .A3(new_n467), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT34), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n478), .B(new_n488), .C1(new_n482), .C2(new_n485), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(KEYINPUT36), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n464), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n326), .A2(new_n327), .ZN(new_n499));
  NOR4_X1   g298(.A1(new_n492), .A2(new_n428), .A3(KEYINPUT35), .A4(new_n438), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n323), .A2(new_n320), .ZN(new_n502));
  INV_X1    g301(.A(new_n428), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n490), .A2(new_n503), .A3(new_n491), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n502), .A2(new_n504), .A3(new_n462), .A4(new_n317), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n461), .A2(new_n498), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n508), .B(KEYINPUT94), .Z(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT95), .ZN(new_n512));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT92), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n513), .A2(KEYINPUT92), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT93), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n510), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n508), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n517), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT16), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n530));
  OAI221_X1 g329(.A(new_n529), .B1(new_n530), .B2(G8gat), .C1(new_n528), .C2(new_n527), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT96), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n531), .B(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n522), .A2(new_n525), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n526), .A2(KEYINPUT17), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT97), .Z(new_n543));
  AOI21_X1  g342(.A(KEYINPUT18), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n526), .B(new_n534), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n543), .B(KEYINPUT13), .Z(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(KEYINPUT18), .A3(new_n543), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  NOR2_X1   g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT98), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n554), .B(KEYINPUT91), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n507), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(G99gat), .ZN(new_n564));
  INV_X1    g363(.A(G106gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT8), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n563), .B(new_n566), .C1(G85gat), .C2(G92gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND3_X1  g368(.A1(new_n540), .A2(new_n538), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n536), .A2(new_n571), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT103), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT104), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n580), .B(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT99), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G71gat), .B(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(G64gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(KEYINPUT99), .A3(G57gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT100), .Z(new_n598));
  INV_X1    g397(.A(KEYINPUT9), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n596), .A2(new_n598), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n534), .B1(new_n589), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT102), .Z(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT101), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n603), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n589), .ZN(new_n609));
  XOR2_X1   g408(.A(G127gat), .B(G155gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n608), .B(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n569), .A2(new_n601), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n569), .A2(new_n601), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  AOI21_X1  g420(.A(new_n617), .B1(new_n621), .B2(new_n616), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n623), .B2(new_n621), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n626), .A2(new_n630), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n631), .B2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n588), .A2(new_n614), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n561), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n462), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n528), .ZN(G1324gat));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n499), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n532), .B2(new_n641), .ZN(new_n644));
  MUX2_X1   g443(.A(new_n643), .B(new_n644), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g444(.A(G15gat), .B1(new_n638), .B2(new_n496), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n492), .A2(G15gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n638), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n638), .A2(new_n503), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  AND2_X1   g450(.A1(new_n585), .A2(new_n587), .ZN(new_n652));
  INV_X1    g451(.A(new_n636), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n614), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT107), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n561), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(G29gat), .A3(new_n462), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n461), .A2(new_n498), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n501), .A2(new_n506), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(KEYINPUT109), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n497), .B1(new_n404), .B2(new_n460), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n499), .A2(new_n500), .B1(new_n505), .B2(KEYINPUT35), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n588), .A2(KEYINPUT44), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT44), .B1(new_n507), .B2(new_n588), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n559), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT110), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n462), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n679), .ZN(G1328gat));
  NOR3_X1   g479(.A1(new_n657), .A2(G36gat), .A3(new_n499), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT46), .ZN(new_n682));
  OAI21_X1  g481(.A(G36gat), .B1(new_n678), .B2(new_n499), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1329gat));
  AOI21_X1  g483(.A(new_n676), .B1(new_n671), .B2(new_n673), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT110), .B(new_n672), .C1(new_n669), .C2(new_n670), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n685), .A2(new_n686), .A3(new_n496), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT112), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n496), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n690), .A3(new_n677), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(G43gat), .ZN(new_n693));
  INV_X1    g492(.A(new_n657), .ZN(new_n694));
  INV_X1    g493(.A(new_n492), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n688), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n689), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G43gat), .B1(new_n674), .B2(new_n496), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n696), .A2(KEYINPUT47), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1330gat));
  OR3_X1    g501(.A1(new_n657), .A2(G50gat), .A3(new_n503), .ZN(new_n703));
  OAI21_X1  g502(.A(G50gat), .B1(new_n674), .B2(new_n503), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(KEYINPUT48), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G50gat), .B1(new_n678), .B2(new_n503), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(new_n703), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n707), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g507(.A(new_n614), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n652), .A2(new_n559), .A3(new_n709), .A4(new_n636), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n667), .A3(new_n663), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT113), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(KEYINPUT113), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n438), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n499), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(G1333gat));
  OR3_X1    g521(.A1(new_n714), .A2(G71gat), .A3(new_n492), .ZN(new_n723));
  OAI21_X1  g522(.A(G71gat), .B1(new_n714), .B2(new_n496), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(KEYINPUT50), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1334gat));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n503), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT114), .B(G78gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n559), .A2(new_n614), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n653), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n669), .B2(new_n670), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n438), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G85gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n507), .A2(new_n588), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n733), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n741), .A2(KEYINPUT115), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(KEYINPUT115), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT116), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n653), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n462), .A2(G85gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n737), .B1(new_n749), .B2(new_n750), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n636), .A2(new_n499), .A3(G92gat), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(new_n745), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n499), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G92gat), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G92gat), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT117), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n743), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n741), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n752), .B(KEYINPUT118), .Z(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n755), .A2(KEYINPUT117), .A3(new_n760), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT52), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n759), .A2(new_n767), .ZN(G1337gat));
  NAND2_X1  g567(.A1(new_n735), .A2(new_n690), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n564), .B1(new_n769), .B2(KEYINPUT120), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT120), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n695), .A2(new_n564), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n749), .B2(new_n772), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n636), .A2(G106gat), .A3(new_n503), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n745), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n565), .B1(new_n735), .B2(new_n428), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(KEYINPUT121), .ZN(new_n780));
  INV_X1    g579(.A(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT121), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n763), .A2(new_n781), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT53), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(G1339gat));
  OR2_X1    g584(.A1(new_n625), .A2(KEYINPUT54), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n622), .A2(new_n624), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n625), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n786), .A2(new_n630), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT55), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n632), .B1(new_n789), .B2(KEYINPUT55), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n541), .A2(new_n543), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n545), .A2(new_n546), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n553), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n556), .A2(new_n790), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n614), .B1(new_n652), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n559), .A2(new_n790), .A3(new_n791), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n556), .A2(new_n794), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n588), .B(new_n797), .C1(new_n636), .C2(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n796), .A2(new_n799), .B1(new_n637), .B2(new_n560), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n428), .A3(new_n492), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n754), .A2(new_n462), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n560), .ZN(new_n804));
  XOR2_X1   g603(.A(KEYINPUT122), .B(G113gat), .Z(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1340gat));
  INV_X1    g605(.A(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n653), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n614), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G127gat), .ZN(G1342gat));
  OR3_X1    g610(.A1(new_n803), .A2(G134gat), .A3(new_n588), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT56), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n803), .B2(new_n588), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(KEYINPUT56), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(G1343gat));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n800), .B2(new_n503), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n796), .A2(new_n799), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n637), .A2(new_n560), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT57), .A3(new_n428), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n496), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n348), .B1(new_n826), .B2(new_n560), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n428), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n824), .ZN(new_n829));
  INV_X1    g628(.A(G141gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n559), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n827), .B(new_n831), .C1(new_n834), .C2(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1344gat));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n346), .A3(new_n653), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n653), .A3(new_n825), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(G148gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(G148gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1345gat));
  OAI21_X1  g643(.A(G155gat), .B1(new_n826), .B2(new_n709), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n342), .A3(new_n614), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1346gat));
  NOR3_X1   g646(.A1(new_n826), .A2(new_n343), .A3(new_n588), .ZN(new_n848));
  AOI21_X1  g647(.A(G162gat), .B1(new_n829), .B2(new_n652), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1347gat));
  NAND2_X1  g649(.A1(new_n821), .A2(new_n503), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n499), .A2(new_n438), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n695), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(KEYINPUT124), .A3(new_n695), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(G169gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(new_n560), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n851), .A2(new_n854), .ZN(new_n860));
  AOI21_X1  g659(.A(G169gat), .B1(new_n860), .B2(new_n559), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(G1348gat));
  OAI21_X1  g661(.A(G176gat), .B1(new_n857), .B2(new_n636), .ZN(new_n863));
  INV_X1    g662(.A(G176gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n864), .A3(new_n653), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1349gat));
  NAND3_X1  g665(.A1(new_n855), .A2(new_n614), .A3(new_n856), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G183gat), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n614), .A2(new_n202), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT125), .B1(new_n860), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT60), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n203), .A3(new_n652), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n855), .A2(new_n652), .A3(new_n856), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(G190gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n877), .B2(G190gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(G1351gat));
  NAND2_X1  g680(.A1(new_n853), .A2(new_n496), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n828), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G197gat), .B1(new_n883), .B2(new_n559), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n818), .B2(new_n822), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n559), .A2(G197gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(G1352gat));
  NAND3_X1  g686(.A1(new_n885), .A2(KEYINPUT127), .A3(new_n653), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT126), .B(G204gat), .Z(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT127), .B1(new_n885), .B2(new_n653), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n883), .A2(new_n653), .A3(new_n889), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n891), .A2(new_n892), .B1(new_n895), .B2(new_n896), .ZN(G1353gat));
  INV_X1    g696(.A(G211gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n898), .A3(new_n614), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n885), .A2(new_n614), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT63), .B1(new_n900), .B2(G211gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1354gat));
  INV_X1    g702(.A(G218gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n904), .A3(new_n652), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n885), .A2(new_n652), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n904), .ZN(G1355gat));
endmodule


