

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U556 ( .A(n736), .ZN(n761) );
  NOR2_X2 U557 ( .A1(n525), .A2(n524), .ZN(n882) );
  AND2_X1 U558 ( .A1(n806), .A2(n805), .ZN(n807) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n769) );
  OR2_X1 U560 ( .A1(n791), .A2(KEYINPUT33), .ZN(n796) );
  OR2_X1 U561 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U562 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U563 ( .A(n752), .B(KEYINPUT29), .ZN(n753) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n522), .ZN(n877) );
  NOR2_X1 U565 ( .A1(G651), .A2(n627), .ZN(n650) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(G2104), .ZN(n522) );
  NAND2_X1 U567 ( .A1(G102), .A2(n877), .ZN(n523) );
  XNOR2_X1 U568 ( .A(KEYINPUT91), .B(n523), .ZN(n527) );
  INV_X1 U569 ( .A(G2105), .ZN(n525) );
  XOR2_X1 U570 ( .A(G2104), .B(KEYINPUT65), .Z(n524) );
  AND2_X1 U571 ( .A1(G126), .A2(n882), .ZN(n526) );
  NOR2_X1 U572 ( .A1(n527), .A2(n526), .ZN(n534) );
  XNOR2_X1 U573 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n528) );
  XNOR2_X1 U574 ( .A(n528), .B(KEYINPUT17), .ZN(n530) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  XNOR2_X2 U576 ( .A(n530), .B(n529), .ZN(n876) );
  NAND2_X1 U577 ( .A1(G138), .A2(n876), .ZN(n532) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U579 ( .A1(n881), .A2(G114), .ZN(n531) );
  AND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U582 ( .A(KEYINPUT92), .ZN(n535) );
  XNOR2_X1 U583 ( .A(n536), .B(n535), .ZN(n690) );
  BUF_X1 U584 ( .A(n690), .Z(G164) );
  INV_X1 U585 ( .A(G57), .ZN(G237) );
  INV_X1 U586 ( .A(G132), .ZN(G219) );
  INV_X1 U587 ( .A(G82), .ZN(G220) );
  INV_X1 U588 ( .A(G651), .ZN(n543) );
  NOR2_X1 U589 ( .A1(G543), .A2(n543), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n537), .Z(n649) );
  NAND2_X1 U591 ( .A1(G63), .A2(n649), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NAND2_X1 U593 ( .A1(G51), .A2(n650), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(n540), .ZN(n548) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U597 ( .A1(G89), .A2(n644), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n541), .B(KEYINPUT4), .ZN(n542) );
  XNOR2_X1 U599 ( .A(n542), .B(KEYINPUT80), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n627), .A2(n543), .ZN(n645) );
  NAND2_X1 U601 ( .A1(G76), .A2(n645), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U603 ( .A(n546), .B(KEYINPUT5), .Z(n547) );
  NOR2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT81), .B(n549), .Z(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n550), .Z(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G94), .A2(G452), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U610 ( .A1(G7), .A2(G661), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n552), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U612 ( .A(G223), .ZN(n829) );
  NAND2_X1 U613 ( .A1(n829), .A2(G567), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n553), .Z(G234) );
  NAND2_X1 U615 ( .A1(G56), .A2(n649), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT14), .ZN(n555) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(n555), .ZN(n563) );
  XOR2_X1 U618 ( .A(KEYINPUT74), .B(KEYINPUT12), .Z(n557) );
  NAND2_X1 U619 ( .A1(G81), .A2(n644), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n645), .A2(G68), .ZN(n558) );
  XNOR2_X1 U622 ( .A(KEYINPUT75), .B(n558), .ZN(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U624 ( .A(KEYINPUT13), .B(n561), .ZN(n562) );
  NOR2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G43), .A2(n650), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n1015) );
  INV_X1 U629 ( .A(G860), .ZN(n597) );
  OR2_X1 U630 ( .A1(n1015), .A2(n597), .ZN(G153) );
  NAND2_X1 U631 ( .A1(G64), .A2(n649), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G52), .A2(n650), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G90), .A2(n644), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G77), .A2(n645), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT70), .B(n574), .ZN(G171) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  NAND2_X1 U641 ( .A1(n644), .A2(G92), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G79), .A2(n645), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G54), .A2(n650), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U645 ( .A(KEYINPUT78), .B(n577), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G66), .A2(n649), .ZN(n578) );
  XNOR2_X1 U647 ( .A(KEYINPUT77), .B(n578), .ZN(n579) );
  NOR2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT15), .B(n583), .Z(n1010) );
  INV_X1 U651 ( .A(n1010), .ZN(n613) );
  NOR2_X1 U652 ( .A1(n613), .A2(G868), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT79), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G91), .A2(n644), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G65), .A2(n649), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G78), .A2(n645), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G53), .A2(n650), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U663 ( .A(KEYINPUT72), .B(n593), .Z(G299) );
  INV_X1 U664 ( .A(G868), .ZN(n665) );
  NOR2_X1 U665 ( .A1(G286), .A2(n665), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT82), .ZN(n596) );
  NOR2_X1 U667 ( .A1(G299), .A2(G868), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n597), .A2(G559), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n598), .A2(n613), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT16), .ZN(n600) );
  XOR2_X1 U672 ( .A(KEYINPUT83), .B(n600), .Z(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n1015), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G868), .A2(n613), .ZN(n601) );
  NOR2_X1 U675 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G282) );
  XOR2_X1 U677 ( .A(G2100), .B(KEYINPUT84), .Z(n612) );
  NAND2_X1 U678 ( .A1(n881), .A2(G111), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G135), .A2(n876), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n882), .A2(G123), .ZN(n606) );
  XOR2_X1 U682 ( .A(KEYINPUT18), .B(n606), .Z(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G99), .A2(n877), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n928) );
  XOR2_X1 U686 ( .A(G2096), .B(n928), .Z(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U688 ( .A1(n613), .A2(G559), .ZN(n662) );
  XNOR2_X1 U689 ( .A(n1015), .B(n662), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n614), .A2(G860), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G93), .A2(n644), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G67), .A2(n649), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G80), .A2(n645), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G55), .A2(n650), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n666) );
  XOR2_X1 U698 ( .A(n621), .B(n666), .Z(G145) );
  NAND2_X1 U699 ( .A1(n650), .A2(G49), .ZN(n622) );
  XOR2_X1 U700 ( .A(KEYINPUT85), .B(n622), .Z(n624) );
  NAND2_X1 U701 ( .A1(G651), .A2(G74), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(KEYINPUT86), .B(n625), .ZN(n626) );
  NOR2_X1 U704 ( .A1(n649), .A2(n626), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G88), .A2(n644), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G75), .A2(n645), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G62), .A2(n649), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G50), .A2(n650), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U713 ( .A(KEYINPUT87), .B(n634), .Z(n635) );
  NOR2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G86), .A2(n644), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G61), .A2(n649), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n645), .A2(G73), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n650), .A2(G48), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G85), .A2(n644), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G72), .A2(n645), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U726 ( .A(KEYINPUT69), .B(n648), .ZN(n654) );
  NAND2_X1 U727 ( .A1(G60), .A2(n649), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G47), .A2(n650), .ZN(n651) );
  AND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(G290) );
  XNOR2_X1 U731 ( .A(G288), .B(n1015), .ZN(n661) );
  XOR2_X1 U732 ( .A(n666), .B(KEYINPUT19), .Z(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(KEYINPUT88), .ZN(n658) );
  XNOR2_X1 U734 ( .A(G166), .B(G305), .ZN(n656) );
  INV_X1 U735 ( .A(G299), .ZN(n747) );
  XNOR2_X1 U736 ( .A(n656), .B(n747), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(G290), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n661), .B(n660), .ZN(n899) );
  XNOR2_X1 U740 ( .A(n899), .B(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n663), .A2(G868), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT89), .B(n664), .Z(n668) );
  NAND2_X1 U743 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U754 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U755 ( .A1(G96), .A2(n675), .ZN(n834) );
  NAND2_X1 U756 ( .A1(n834), .A2(G2106), .ZN(n679) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U758 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U759 ( .A1(G108), .A2(n677), .ZN(n835) );
  NAND2_X1 U760 ( .A1(n835), .A2(G567), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n836) );
  NOR2_X1 U762 ( .A1(n680), .A2(n836), .ZN(n681) );
  XNOR2_X1 U763 ( .A(n681), .B(KEYINPUT90), .ZN(n833) );
  NAND2_X1 U764 ( .A1(G36), .A2(n833), .ZN(G176) );
  NAND2_X1 U765 ( .A1(G137), .A2(n876), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n881), .A2(G113), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n689) );
  NAND2_X1 U768 ( .A1(n882), .A2(G125), .ZN(n684) );
  XNOR2_X1 U769 ( .A(n684), .B(KEYINPUT66), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G101), .A2(n877), .ZN(n685) );
  XOR2_X1 U771 ( .A(KEYINPUT23), .B(n685), .Z(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n689), .A2(n688), .ZN(G160) );
  XNOR2_X1 U774 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  XNOR2_X1 U775 ( .A(G1986), .B(G290), .ZN(n1003) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n690), .A2(G1384), .ZN(n691) );
  XNOR2_X1 U778 ( .A(n691), .B(KEYINPUT64), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n723), .A2(n721), .ZN(n824) );
  NAND2_X1 U780 ( .A1(n1003), .A2(n824), .ZN(n812) );
  NAND2_X1 U781 ( .A1(G131), .A2(n876), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G95), .A2(n877), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n881), .A2(G107), .ZN(n695) );
  NAND2_X1 U785 ( .A1(G119), .A2(n882), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n863) );
  INV_X1 U788 ( .A(G1991), .ZN(n951) );
  NOR2_X1 U789 ( .A1(n863), .A2(n951), .ZN(n707) );
  NAND2_X1 U790 ( .A1(n881), .A2(G117), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G141), .A2(n876), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n877), .A2(G105), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT38), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n882), .A2(G129), .ZN(n701) );
  XOR2_X1 U796 ( .A(KEYINPUT95), .B(n701), .Z(n702) );
  NAND2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n890) );
  INV_X1 U799 ( .A(G1996), .ZN(n817) );
  NOR2_X1 U800 ( .A1(n890), .A2(n817), .ZN(n706) );
  NOR2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n933) );
  INV_X1 U802 ( .A(n824), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n933), .A2(n708), .ZN(n816) );
  INV_X1 U804 ( .A(n816), .ZN(n719) );
  NAND2_X1 U805 ( .A1(G140), .A2(n876), .ZN(n710) );
  NAND2_X1 U806 ( .A1(G104), .A2(n877), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n711), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n881), .A2(G116), .ZN(n713) );
  NAND2_X1 U810 ( .A1(G128), .A2(n882), .ZN(n712) );
  NAND2_X1 U811 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U812 ( .A(n714), .B(KEYINPUT35), .Z(n715) );
  NOR2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U814 ( .A(KEYINPUT36), .B(n717), .Z(n718) );
  XOR2_X1 U815 ( .A(KEYINPUT94), .B(n718), .Z(n895) );
  XNOR2_X1 U816 ( .A(G2067), .B(KEYINPUT37), .ZN(n813) );
  NOR2_X1 U817 ( .A1(n895), .A2(n813), .ZN(n942) );
  NAND2_X1 U818 ( .A1(n824), .A2(n942), .ZN(n822) );
  NAND2_X1 U819 ( .A1(n719), .A2(n822), .ZN(n720) );
  XOR2_X1 U820 ( .A(n720), .B(KEYINPUT96), .Z(n810) );
  INV_X1 U821 ( .A(n721), .ZN(n722) );
  NOR2_X2 U822 ( .A1(n723), .A2(n722), .ZN(n736) );
  INV_X1 U823 ( .A(n761), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NAND2_X1 U825 ( .A1(n732), .A2(n957), .ZN(n724) );
  XNOR2_X1 U826 ( .A(n724), .B(KEYINPUT98), .ZN(n726) );
  XNOR2_X1 U827 ( .A(G1961), .B(KEYINPUT97), .ZN(n971) );
  INV_X1 U828 ( .A(n732), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n971), .A2(n755), .ZN(n725) );
  NAND2_X1 U830 ( .A1(n726), .A2(n725), .ZN(n766) );
  AND2_X1 U831 ( .A1(G171), .A2(n766), .ZN(n727) );
  XNOR2_X1 U832 ( .A(n727), .B(KEYINPUT99), .ZN(n754) );
  NOR2_X1 U833 ( .A1(n761), .A2(n817), .ZN(n728) );
  XNOR2_X1 U834 ( .A(n728), .B(KEYINPUT26), .ZN(n730) );
  AND2_X1 U835 ( .A1(n761), .A2(G1341), .ZN(n729) );
  NOR2_X1 U836 ( .A1(n1015), .A2(n731), .ZN(n741) );
  NAND2_X1 U837 ( .A1(G1348), .A2(n755), .ZN(n734) );
  NAND2_X1 U838 ( .A1(G2067), .A2(n732), .ZN(n733) );
  NAND2_X1 U839 ( .A1(n734), .A2(n733), .ZN(n742) );
  NOR2_X1 U840 ( .A1(n742), .A2(n1010), .ZN(n739) );
  NAND2_X1 U841 ( .A1(n736), .A2(G2072), .ZN(n735) );
  XNOR2_X1 U842 ( .A(n735), .B(KEYINPUT27), .ZN(n738) );
  INV_X1 U843 ( .A(G1956), .ZN(n979) );
  NOR2_X1 U844 ( .A1(n979), .A2(n736), .ZN(n737) );
  NOR2_X1 U845 ( .A1(n738), .A2(n737), .ZN(n748) );
  AND2_X1 U846 ( .A1(n748), .A2(n747), .ZN(n744) );
  OR2_X1 U847 ( .A1(n739), .A2(n744), .ZN(n740) );
  NOR2_X1 U848 ( .A1(n741), .A2(n740), .ZN(n746) );
  NAND2_X1 U849 ( .A1(n1010), .A2(n742), .ZN(n743) );
  NOR2_X1 U850 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U851 ( .A1(n746), .A2(n745), .ZN(n751) );
  NOR2_X1 U852 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U853 ( .A(n749), .B(KEYINPUT28), .Z(n750) );
  NAND2_X1 U854 ( .A1(n754), .A2(n753), .ZN(n779) );
  INV_X1 U855 ( .A(G8), .ZN(n760) );
  NAND2_X1 U856 ( .A1(G8), .A2(n761), .ZN(n803) );
  NOR2_X1 U857 ( .A1(G1971), .A2(n803), .ZN(n757) );
  NOR2_X1 U858 ( .A1(G2090), .A2(n755), .ZN(n756) );
  NOR2_X1 U859 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U860 ( .A1(n758), .A2(G303), .ZN(n759) );
  OR2_X1 U861 ( .A1(n760), .A2(n759), .ZN(n772) );
  AND2_X1 U862 ( .A1(n779), .A2(n772), .ZN(n771) );
  NOR2_X1 U863 ( .A1(G1966), .A2(n803), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G2084), .A2(n761), .ZN(n777) );
  NOR2_X1 U865 ( .A1(n781), .A2(n777), .ZN(n762) );
  NAND2_X1 U866 ( .A1(G8), .A2(n762), .ZN(n763) );
  XNOR2_X1 U867 ( .A(KEYINPUT100), .B(n763), .ZN(n764) );
  XNOR2_X1 U868 ( .A(n764), .B(KEYINPUT30), .ZN(n765) );
  NOR2_X1 U869 ( .A1(n765), .A2(G168), .ZN(n768) );
  NOR2_X1 U870 ( .A1(n766), .A2(G171), .ZN(n767) );
  NOR2_X1 U871 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U872 ( .A(n770), .B(n769), .ZN(n778) );
  NAND2_X1 U873 ( .A1(n771), .A2(n778), .ZN(n775) );
  INV_X1 U874 ( .A(n772), .ZN(n773) );
  OR2_X1 U875 ( .A1(n773), .A2(G286), .ZN(n774) );
  NAND2_X1 U876 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U877 ( .A(n776), .B(KEYINPUT32), .ZN(n785) );
  NAND2_X1 U878 ( .A1(G8), .A2(n777), .ZN(n783) );
  AND2_X1 U879 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U880 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U881 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n801) );
  NOR2_X1 U883 ( .A1(G1976), .A2(G288), .ZN(n998) );
  NOR2_X1 U884 ( .A1(G1971), .A2(G303), .ZN(n786) );
  NOR2_X1 U885 ( .A1(n998), .A2(n786), .ZN(n787) );
  XOR2_X1 U886 ( .A(KEYINPUT101), .B(n787), .Z(n788) );
  NAND2_X1 U887 ( .A1(n801), .A2(n788), .ZN(n789) );
  NAND2_X1 U888 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NAND2_X1 U889 ( .A1(n789), .A2(n1000), .ZN(n790) );
  NOR2_X1 U890 ( .A1(n790), .A2(n803), .ZN(n791) );
  XOR2_X1 U891 ( .A(G1981), .B(G305), .Z(n1018) );
  INV_X1 U892 ( .A(n1018), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n998), .A2(KEYINPUT33), .ZN(n792) );
  NOR2_X1 U894 ( .A1(n792), .A2(n803), .ZN(n793) );
  NOR2_X1 U895 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U896 ( .A1(n796), .A2(n795), .ZN(n808) );
  NOR2_X1 U897 ( .A1(G1981), .A2(G305), .ZN(n797) );
  XOR2_X1 U898 ( .A(n797), .B(KEYINPUT24), .Z(n798) );
  OR2_X1 U899 ( .A1(n803), .A2(n798), .ZN(n806) );
  NOR2_X1 U900 ( .A1(G2090), .A2(G303), .ZN(n799) );
  NAND2_X1 U901 ( .A1(G8), .A2(n799), .ZN(n800) );
  NAND2_X1 U902 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U903 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U904 ( .A(n804), .B(KEYINPUT102), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  AND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n827) );
  NAND2_X1 U908 ( .A1(n895), .A2(n813), .ZN(n939) );
  XNOR2_X1 U909 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n820) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n814) );
  AND2_X1 U911 ( .A1(n951), .A2(n863), .ZN(n931) );
  NOR2_X1 U912 ( .A1(n814), .A2(n931), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n818) );
  AND2_X1 U914 ( .A1(n817), .A2(n890), .ZN(n935) );
  NOR2_X1 U915 ( .A1(n818), .A2(n935), .ZN(n819) );
  XOR2_X1 U916 ( .A(n820), .B(n819), .Z(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n939), .A2(n823), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(n829), .A2(G2106), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT107), .B(n830), .Z(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U925 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G188) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G325) );
  XOR2_X1 U929 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U930 ( .A(n836), .ZN(G319) );
  XOR2_X1 U931 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U932 ( .A(KEYINPUT109), .B(G2678), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U934 ( .A(KEYINPUT42), .B(G2090), .Z(n840) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U938 ( .A(G2100), .B(G2096), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n846) );
  XOR2_X1 U940 ( .A(G2078), .B(G2084), .Z(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1971), .B(G1956), .Z(n848) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1976), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U945 ( .A(n849), .B(G2474), .Z(n851) );
  XNOR2_X1 U946 ( .A(G1981), .B(G1966), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U948 ( .A(KEYINPUT41), .B(G1961), .Z(n853) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U952 ( .A1(n881), .A2(G112), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G136), .A2(n876), .ZN(n856) );
  NAND2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U955 ( .A1(n882), .A2(G124), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G100), .A2(n877), .ZN(n859) );
  NAND2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U959 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n865) );
  XNOR2_X1 U961 ( .A(n863), .B(KEYINPUT114), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n894) );
  NAND2_X1 U963 ( .A1(n881), .A2(G118), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G130), .A2(n882), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G142), .A2(n876), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G106), .A2(n877), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT45), .B(n870), .ZN(n871) );
  XNOR2_X1 U970 ( .A(KEYINPUT111), .B(n871), .ZN(n872) );
  NOR2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U972 ( .A(G162), .B(n874), .Z(n875) );
  XNOR2_X1 U973 ( .A(n928), .B(n875), .ZN(n889) );
  NAND2_X1 U974 ( .A1(G139), .A2(n876), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G103), .A2(n877), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U977 ( .A(KEYINPUT112), .B(n880), .ZN(n888) );
  NAND2_X1 U978 ( .A1(n881), .A2(G115), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U981 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(n886), .ZN(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n923) );
  XOR2_X1 U984 ( .A(n889), .B(n923), .Z(n892) );
  XNOR2_X1 U985 ( .A(G160), .B(n890), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U988 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U990 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n1010), .ZN(n900) );
  XNOR2_X1 U992 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n901), .B(G171), .ZN(n902) );
  NOR2_X1 U994 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2451), .B(KEYINPUT106), .Z(n904) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2446), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U998 ( .A(G2435), .B(KEYINPUT105), .Z(n906) );
  XNOR2_X1 U999 ( .A(G2438), .B(G2454), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1001 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1002 ( .A(G2427), .B(KEYINPUT104), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n913) );
  XOR2_X1 U1004 ( .A(G1341), .B(G1348), .Z(n911) );
  XNOR2_X1 U1005 ( .A(G2430), .B(n911), .ZN(n912) );
  XOR2_X1 U1006 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1007 ( .A1(G14), .A2(n914), .ZN(n921) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n915) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  XNOR2_X1 U1011 ( .A(n916), .B(KEYINPUT115), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(G225) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1017 ( .A(G120), .ZN(G236) );
  INV_X1 U1018 ( .A(G96), .ZN(G221) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  INV_X1 U1021 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(G2078), .B(KEYINPUT119), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(n922), .B(G164), .ZN(n926) );
  XOR2_X1 U1024 ( .A(G2072), .B(KEYINPUT118), .Z(n924) );
  XNOR2_X1 U1025 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n927), .Z(n945) );
  XNOR2_X1 U1028 ( .A(G160), .B(G2084), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n936), .B(KEYINPUT51), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT117), .B(n943), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n967), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G25), .B(n951), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n952), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G26), .B(G2067), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1053 ( .A(G27), .B(n957), .Z(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1061 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n970), .ZN(n1028) );
  XNOR2_X1 U1064 ( .A(G5), .B(n971), .ZN(n992) );
  XOR2_X1 U1065 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n978) );
  XNOR2_X1 U1066 ( .A(G1976), .B(G23), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1069 ( .A(G1986), .B(KEYINPUT124), .Z(n974) );
  XNOR2_X1 U1070 ( .A(G24), .B(n974), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n978), .B(n977), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G20), .B(n979), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT59), .B(G1348), .Z(n984) );
  XNOR2_X1 U1079 ( .A(G4), .B(n984), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT123), .B(n987), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(KEYINPUT60), .B(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G21), .B(G1966), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(KEYINPUT61), .B(n995), .Z(n996) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n996), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(n997), .Z(n1026) );
  XNOR2_X1 U1090 ( .A(KEYINPUT56), .B(G16), .ZN(n1024) );
  INV_X1 U1091 ( .A(n998), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT121), .ZN(n1014) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G299), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G1971), .B(KEYINPUT122), .ZN(n1004) );
  XNOR2_X1 U1097 ( .A(n1004), .B(G303), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(G301), .B(G1961), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(n1005), .B(KEYINPUT120), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G1348), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G1341), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G168), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(n1020), .B(KEYINPUT57), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(n1031), .B(KEYINPUT62), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(KEYINPUT127), .B(n1032), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

