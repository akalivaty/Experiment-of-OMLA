

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756;

  BUF_X1 U372 ( .A(n590), .Z(n597) );
  NAND2_X1 U373 ( .A1(G214), .A2(n471), .ZN(n692) );
  XNOR2_X2 U374 ( .A(n455), .B(n454), .ZN(n456) );
  AND2_X2 U375 ( .A1(n636), .A2(KEYINPUT86), .ZN(n592) );
  AND2_X2 U376 ( .A1(n377), .A2(n375), .ZN(n374) );
  NAND2_X2 U377 ( .A1(n751), .A2(n657), .ZN(n573) );
  NOR2_X1 U378 ( .A1(n532), .A2(n533), .ZN(n568) );
  NAND2_X1 U379 ( .A1(n516), .A2(n692), .ZN(n395) );
  XNOR2_X2 U380 ( .A(KEYINPUT18), .B(KEYINPUT77), .ZN(n398) );
  XNOR2_X2 U381 ( .A(n450), .B(G134), .ZN(n461) );
  XNOR2_X2 U382 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n457) );
  INV_X1 U383 ( .A(n677), .ZN(n575) );
  XNOR2_X1 U384 ( .A(n391), .B(n630), .ZN(n631) );
  AND2_X1 U385 ( .A1(n388), .A2(n385), .ZN(n384) );
  INV_X1 U386 ( .A(n604), .ZN(n351) );
  NAND2_X1 U387 ( .A1(n681), .A2(n680), .ZN(n677) );
  XNOR2_X2 U388 ( .A(n367), .B(KEYINPUT45), .ZN(n725) );
  NOR2_X2 U389 ( .A1(n617), .A2(n616), .ZN(n367) );
  XNOR2_X2 U390 ( .A(n741), .B(G146), .ZN(n380) );
  XNOR2_X2 U391 ( .A(n460), .B(n461), .ZN(n741) );
  OR2_X2 U392 ( .A1(n362), .A2(n390), .ZN(n391) );
  XOR2_X2 U393 ( .A(KEYINPUT68), .B(G101), .Z(n462) );
  XNOR2_X1 U394 ( .A(n439), .B(n438), .ZN(n467) );
  NAND2_X1 U395 ( .A1(n437), .A2(n436), .ZN(n439) );
  XNOR2_X1 U396 ( .A(KEYINPUT3), .B(G119), .ZN(n438) );
  NOR2_X1 U397 ( .A1(G953), .A2(G237), .ZN(n463) );
  XNOR2_X1 U398 ( .A(n457), .B(n379), .ZN(n449) );
  INV_X1 U399 ( .A(KEYINPUT79), .ZN(n379) );
  XNOR2_X1 U400 ( .A(n365), .B(n577), .ZN(n604) );
  OR2_X1 U401 ( .A1(n637), .A2(G902), .ZN(n470) );
  XNOR2_X1 U402 ( .A(n446), .B(n445), .ZN(n733) );
  NAND2_X1 U403 ( .A1(n444), .A2(n443), .ZN(n446) );
  XNOR2_X1 U404 ( .A(KEYINPUT76), .B(G110), .ZN(n445) );
  XNOR2_X1 U405 ( .A(n467), .B(n401), .ZN(n734) );
  XNOR2_X1 U406 ( .A(n440), .B(G122), .ZN(n401) );
  XNOR2_X1 U407 ( .A(n742), .B(n409), .ZN(n422) );
  XNOR2_X1 U408 ( .A(n458), .B(n410), .ZN(n409) );
  XNOR2_X1 U409 ( .A(n402), .B(n733), .ZN(n477) );
  XNOR2_X1 U410 ( .A(n462), .B(KEYINPUT72), .ZN(n402) );
  INV_X1 U411 ( .A(KEYINPUT39), .ZN(n363) );
  AND2_X1 U412 ( .A1(n386), .A2(n584), .ZN(n385) );
  NAND2_X1 U413 ( .A1(n605), .A2(n387), .ZN(n386) );
  INV_X1 U414 ( .A(n361), .ZN(n387) );
  NOR2_X1 U415 ( .A1(n678), .A2(KEYINPUT103), .ZN(n376) );
  NAND2_X1 U416 ( .A1(n568), .A2(n680), .ZN(n389) );
  INV_X1 U417 ( .A(KEYINPUT64), .ZN(n430) );
  XNOR2_X1 U418 ( .A(n412), .B(G125), .ZN(n447) );
  INV_X1 U419 ( .A(G146), .ZN(n412) );
  XNOR2_X1 U420 ( .A(G113), .B(G122), .ZN(n410) );
  XNOR2_X1 U421 ( .A(n421), .B(G131), .ZN(n458) );
  XNOR2_X1 U422 ( .A(G143), .B(G104), .ZN(n417) );
  XOR2_X1 U423 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n418) );
  XOR2_X1 U424 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n416) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n501) );
  XNOR2_X1 U426 ( .A(n433), .B(G478), .ZN(n532) );
  XNOR2_X1 U427 ( .A(n372), .B(KEYINPUT0), .ZN(n582) );
  XNOR2_X1 U428 ( .A(n380), .B(n468), .ZN(n637) );
  XNOR2_X1 U429 ( .A(G128), .B(G110), .ZN(n482) );
  XOR2_X1 U430 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n483) );
  XNOR2_X1 U431 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U432 ( .A(KEYINPUT24), .ZN(n484) );
  XNOR2_X1 U433 ( .A(G119), .B(G137), .ZN(n485) );
  XNOR2_X1 U434 ( .A(n431), .B(n394), .ZN(n489) );
  INV_X1 U435 ( .A(KEYINPUT8), .ZN(n394) );
  XNOR2_X1 U436 ( .A(n447), .B(n411), .ZN(n742) );
  XNOR2_X1 U437 ( .A(G140), .B(KEYINPUT10), .ZN(n411) );
  XNOR2_X1 U438 ( .A(G116), .B(G122), .ZN(n425) );
  NAND2_X1 U439 ( .A1(n489), .A2(G217), .ZN(n393) );
  XNOR2_X1 U440 ( .A(G107), .B(KEYINPUT7), .ZN(n426) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n427) );
  XNOR2_X1 U442 ( .A(n734), .B(n477), .ZN(n370) );
  INV_X1 U443 ( .A(KEYINPUT1), .ZN(n404) );
  XNOR2_X1 U444 ( .A(n524), .B(KEYINPUT105), .ZN(n525) );
  AND2_X1 U445 ( .A1(n508), .A2(n507), .ZN(n530) );
  AND2_X1 U446 ( .A1(n506), .A2(n414), .ZN(n507) );
  XNOR2_X1 U447 ( .A(n408), .B(n407), .ZN(n533) );
  XNOR2_X1 U448 ( .A(G475), .B(n424), .ZN(n407) );
  OR2_X1 U449 ( .A1(n621), .A2(G902), .ZN(n408) );
  BUF_X1 U450 ( .A(n599), .Z(n403) );
  XNOR2_X1 U451 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U452 ( .A(n380), .B(n478), .ZN(n645) );
  INV_X1 U453 ( .A(G140), .ZN(n474) );
  NAND2_X1 U454 ( .A1(n492), .A2(G210), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n368), .B(KEYINPUT40), .ZN(n752) );
  NOR2_X1 U456 ( .A1(n552), .A2(n531), .ZN(n368) );
  NAND2_X1 U457 ( .A1(n384), .A2(n382), .ZN(n585) );
  NAND2_X1 U458 ( .A1(n383), .A2(n387), .ZN(n382) );
  NOR2_X1 U459 ( .A1(n376), .A2(n358), .ZN(n375) );
  AND2_X1 U460 ( .A1(n598), .A2(n361), .ZN(n352) );
  AND2_X1 U461 ( .A1(n678), .A2(KEYINPUT103), .ZN(n353) );
  XOR2_X1 U462 ( .A(n480), .B(G469), .Z(n354) );
  XOR2_X1 U463 ( .A(n389), .B(KEYINPUT101), .Z(n355) );
  BUF_X1 U464 ( .A(n582), .Z(n605) );
  AND2_X1 U465 ( .A1(n572), .A2(n406), .ZN(n356) );
  AND2_X1 U466 ( .A1(n396), .A2(n678), .ZN(n357) );
  NAND2_X1 U467 ( .A1(n571), .A2(n406), .ZN(n358) );
  AND2_X1 U468 ( .A1(n528), .A2(n635), .ZN(n359) );
  OR2_X1 U469 ( .A1(n549), .A2(n413), .ZN(n360) );
  XNOR2_X1 U470 ( .A(n684), .B(n521), .ZN(n609) );
  XOR2_X1 U471 ( .A(KEYINPUT80), .B(KEYINPUT34), .Z(n361) );
  NAND2_X2 U472 ( .A1(n374), .A2(n373), .ZN(n657) );
  XNOR2_X1 U473 ( .A(n581), .B(n580), .ZN(n709) );
  NOR2_X2 U474 ( .A1(n362), .A2(n619), .ZN(n644) );
  AND2_X1 U475 ( .A1(n362), .A2(n713), .ZN(n714) );
  XNOR2_X2 U476 ( .A(n618), .B(KEYINPUT2), .ZN(n362) );
  XNOR2_X1 U477 ( .A(n364), .B(n363), .ZN(n552) );
  NAND2_X1 U478 ( .A1(n530), .A2(n693), .ZN(n364) );
  NAND2_X1 U479 ( .A1(n351), .A2(n609), .ZN(n581) );
  NAND2_X1 U480 ( .A1(n575), .A2(n576), .ZN(n365) );
  AND2_X1 U481 ( .A1(n366), .A2(n359), .ZN(n551) );
  NOR2_X1 U482 ( .A1(n542), .A2(n360), .ZN(n366) );
  NOR2_X2 U483 ( .A1(n725), .A2(n743), .ZN(n618) );
  XNOR2_X2 U484 ( .A(n369), .B(n456), .ZN(n516) );
  XNOR2_X2 U485 ( .A(n569), .B(KEYINPUT22), .ZN(n396) );
  OR2_X2 U486 ( .A1(n627), .A2(n492), .ZN(n369) );
  XNOR2_X1 U487 ( .A(n371), .B(n370), .ZN(n627) );
  XNOR2_X1 U488 ( .A(n452), .B(n451), .ZN(n371) );
  NOR2_X2 U489 ( .A1(n582), .A2(n355), .ZN(n569) );
  NAND2_X1 U490 ( .A1(n567), .A2(n566), .ZN(n372) );
  XNOR2_X2 U491 ( .A(n395), .B(KEYINPUT19), .ZN(n567) );
  OR2_X1 U492 ( .A1(n396), .A2(KEYINPUT103), .ZN(n373) );
  NAND2_X1 U493 ( .A1(n396), .A2(n353), .ZN(n377) );
  XNOR2_X2 U494 ( .A(n378), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U495 ( .A1(n396), .A2(n356), .ZN(n378) );
  XNOR2_X2 U496 ( .A(n381), .B(G143), .ZN(n450) );
  XNOR2_X2 U497 ( .A(G128), .B(KEYINPUT66), .ZN(n381) );
  INV_X1 U498 ( .A(n709), .ZN(n383) );
  NAND2_X1 U499 ( .A1(n709), .A2(n352), .ZN(n388) );
  XNOR2_X1 U500 ( .A(n392), .B(n432), .ZN(n715) );
  XNOR2_X1 U501 ( .A(n393), .B(n461), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X2 U503 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n397) );
  XNOR2_X1 U504 ( .A(n399), .B(n447), .ZN(n400) );
  XNOR2_X1 U505 ( .A(n400), .B(n448), .ZN(n452) );
  NAND2_X1 U506 ( .A1(n567), .A2(n405), .ZN(n517) );
  XNOR2_X2 U507 ( .A(n599), .B(n404), .ZN(n576) );
  NAND2_X1 U508 ( .A1(n536), .A2(n405), .ZN(n537) );
  INV_X1 U509 ( .A(n403), .ZN(n405) );
  XNOR2_X2 U510 ( .A(n481), .B(n354), .ZN(n599) );
  INV_X1 U511 ( .A(n681), .ZN(n406) );
  BUF_X1 U512 ( .A(n627), .Z(n629) );
  XNOR2_X1 U513 ( .A(n590), .B(n574), .ZN(n586) );
  XNOR2_X2 U514 ( .A(n430), .B(G953), .ZN(n745) );
  AND2_X1 U515 ( .A1(KEYINPUT47), .A2(n548), .ZN(n413) );
  OR2_X1 U516 ( .A1(n564), .A2(n505), .ZN(n414) );
  INV_X1 U517 ( .A(KEYINPUT87), .ZN(n574) );
  INV_X1 U518 ( .A(KEYINPUT46), .ZN(n540) );
  NOR2_X1 U519 ( .A1(n589), .A2(n588), .ZN(n595) );
  XNOR2_X1 U520 ( .A(n487), .B(n486), .ZN(n488) );
  OR2_X1 U521 ( .A1(n745), .A2(G952), .ZN(n640) );
  INV_X1 U522 ( .A(KEYINPUT60), .ZN(n625) );
  NAND2_X1 U523 ( .A1(G214), .A2(n463), .ZN(n415) );
  XNOR2_X1 U524 ( .A(n416), .B(n415), .ZN(n420) );
  XNOR2_X1 U525 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U526 ( .A(n420), .B(n419), .Z(n423) );
  INV_X1 U527 ( .A(KEYINPUT69), .ZN(n421) );
  XNOR2_X1 U528 ( .A(n423), .B(n422), .ZN(n621) );
  INV_X1 U529 ( .A(KEYINPUT13), .ZN(n424) );
  XNOR2_X1 U530 ( .A(n425), .B(KEYINPUT99), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U532 ( .A(n429), .B(n428), .Z(n432) );
  NAND2_X1 U533 ( .A1(n745), .A2(G234), .ZN(n431) );
  INV_X1 U534 ( .A(G902), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n715), .A2(n479), .ZN(n433) );
  NAND2_X1 U536 ( .A1(n533), .A2(n532), .ZN(n583) );
  XOR2_X1 U537 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n440) );
  INV_X1 U538 ( .A(G116), .ZN(n434) );
  NAND2_X1 U539 ( .A1(G113), .A2(n434), .ZN(n437) );
  INV_X1 U540 ( .A(G113), .ZN(n435) );
  NAND2_X1 U541 ( .A1(n435), .A2(G116), .ZN(n436) );
  INV_X1 U542 ( .A(G107), .ZN(n441) );
  NAND2_X1 U543 ( .A1(G104), .A2(n441), .ZN(n444) );
  INV_X1 U544 ( .A(G104), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n442), .A2(G107), .ZN(n443) );
  NAND2_X1 U546 ( .A1(G224), .A2(n745), .ZN(n448) );
  XOR2_X1 U547 ( .A(n450), .B(n449), .Z(n451) );
  INV_X1 U548 ( .A(KEYINPUT15), .ZN(n453) );
  XNOR2_X1 U549 ( .A(n453), .B(G902), .ZN(n492) );
  XOR2_X1 U550 ( .A(KEYINPUT91), .B(KEYINPUT81), .Z(n455) );
  OR2_X1 U551 ( .A1(G237), .A2(G902), .ZN(n471) );
  NAND2_X1 U552 ( .A1(G210), .A2(n471), .ZN(n454) );
  BUF_X2 U553 ( .A(n516), .Z(n556) );
  XNOR2_X1 U554 ( .A(n457), .B(G137), .ZN(n459) );
  XNOR2_X1 U555 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U556 ( .A(n462), .B(KEYINPUT5), .Z(n465) );
  NAND2_X1 U557 ( .A1(n463), .A2(G210), .ZN(n464) );
  XNOR2_X1 U558 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U559 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U560 ( .A(G472), .B(KEYINPUT73), .Z(n469) );
  XNOR2_X2 U561 ( .A(n470), .B(n469), .ZN(n520) );
  XNOR2_X2 U562 ( .A(n520), .B(KEYINPUT102), .ZN(n570) );
  NAND2_X1 U563 ( .A1(n570), .A2(n692), .ZN(n473) );
  XOR2_X1 U564 ( .A(KEYINPUT106), .B(KEYINPUT30), .Z(n472) );
  XNOR2_X1 U565 ( .A(n473), .B(n472), .ZN(n508) );
  NAND2_X1 U566 ( .A1(n745), .A2(G227), .ZN(n475) );
  XNOR2_X1 U567 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U568 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U569 ( .A1(n645), .A2(n479), .ZN(n481) );
  INV_X1 U570 ( .A(KEYINPUT71), .ZN(n480) );
  XNOR2_X1 U571 ( .A(n483), .B(n482), .ZN(n487) );
  XOR2_X1 U572 ( .A(n742), .B(n488), .Z(n491) );
  NAND2_X1 U573 ( .A1(G221), .A2(n489), .ZN(n490) );
  XNOR2_X1 U574 ( .A(n491), .B(n490), .ZN(n720) );
  NOR2_X1 U575 ( .A1(n720), .A2(G902), .ZN(n496) );
  XOR2_X1 U576 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n494) );
  INV_X1 U577 ( .A(n492), .ZN(n619) );
  NAND2_X1 U578 ( .A1(G234), .A2(n619), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n494), .B(n493), .ZN(n498) );
  NAND2_X1 U580 ( .A1(n498), .A2(G217), .ZN(n495) );
  XNOR2_X1 U581 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X2 U582 ( .A(n497), .B(KEYINPUT25), .ZN(n681) );
  NAND2_X1 U583 ( .A1(n498), .A2(G221), .ZN(n500) );
  INV_X1 U584 ( .A(KEYINPUT21), .ZN(n499) );
  XNOR2_X1 U585 ( .A(n500), .B(n499), .ZN(n680) );
  NOR2_X1 U586 ( .A1(n403), .A2(n677), .ZN(n506) );
  XNOR2_X1 U587 ( .A(n501), .B(KEYINPUT14), .ZN(n502) );
  NAND2_X1 U588 ( .A1(G952), .A2(n502), .ZN(n707) );
  NOR2_X1 U589 ( .A1(G953), .A2(n707), .ZN(n564) );
  INV_X1 U590 ( .A(n745), .ZN(n503) );
  AND2_X1 U591 ( .A1(G902), .A2(n502), .ZN(n561) );
  NAND2_X1 U592 ( .A1(n503), .A2(n561), .ZN(n504) );
  NOR2_X1 U593 ( .A1(G900), .A2(n504), .ZN(n505) );
  NAND2_X1 U594 ( .A1(n556), .A2(n530), .ZN(n509) );
  NOR2_X1 U595 ( .A1(n583), .A2(n509), .ZN(n662) );
  XNOR2_X1 U596 ( .A(KEYINPUT85), .B(n662), .ZN(n512) );
  INV_X1 U597 ( .A(n532), .ZN(n510) );
  NOR2_X1 U598 ( .A1(n510), .A2(n533), .ZN(n658) );
  INV_X1 U599 ( .A(n658), .ZN(n672) );
  NAND2_X1 U600 ( .A1(n533), .A2(n510), .ZN(n531) );
  NAND2_X1 U601 ( .A1(n672), .A2(n531), .ZN(n696) );
  NAND2_X1 U602 ( .A1(n696), .A2(KEYINPUT83), .ZN(n511) );
  NAND2_X1 U603 ( .A1(n512), .A2(n511), .ZN(n519) );
  NAND2_X1 U604 ( .A1(n414), .A2(n680), .ZN(n513) );
  NOR2_X1 U605 ( .A1(n681), .A2(n513), .ZN(n523) );
  AND2_X1 U606 ( .A1(n570), .A2(n523), .ZN(n515) );
  XNOR2_X1 U607 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n514) );
  XNOR2_X1 U608 ( .A(n515), .B(n514), .ZN(n538) );
  NOR2_X1 U609 ( .A1(n538), .A2(n517), .ZN(n659) );
  INV_X1 U610 ( .A(n659), .ZN(n663) );
  NOR2_X1 U611 ( .A1(KEYINPUT82), .A2(n663), .ZN(n518) );
  NOR2_X1 U612 ( .A1(n519), .A2(n518), .ZN(n528) );
  INV_X1 U613 ( .A(n556), .ZN(n529) );
  XNOR2_X1 U614 ( .A(KEYINPUT104), .B(n531), .ZN(n667) );
  BUF_X2 U615 ( .A(n520), .Z(n684) );
  INV_X1 U616 ( .A(KEYINPUT6), .ZN(n521) );
  INV_X1 U617 ( .A(n609), .ZN(n578) );
  NOR2_X1 U618 ( .A1(n667), .A2(n578), .ZN(n522) );
  NAND2_X1 U619 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U620 ( .A1(n525), .A2(n692), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n529), .A2(n554), .ZN(n526) );
  XNOR2_X1 U622 ( .A(n526), .B(KEYINPUT36), .ZN(n527) );
  NAND2_X1 U623 ( .A1(n527), .A2(n576), .ZN(n635) );
  XNOR2_X1 U624 ( .A(KEYINPUT38), .B(n529), .ZN(n693) );
  NAND2_X1 U625 ( .A1(n693), .A2(n692), .ZN(n697) );
  INV_X1 U626 ( .A(n568), .ZN(n695) );
  NOR2_X1 U627 ( .A1(n697), .A2(n695), .ZN(n535) );
  XNOR2_X1 U628 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n535), .B(n534), .ZN(n710) );
  INV_X1 U630 ( .A(n710), .ZN(n536) );
  NOR2_X1 U631 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U632 ( .A(n539), .B(KEYINPUT42), .ZN(n756) );
  NOR2_X1 U633 ( .A1(n752), .A2(n756), .ZN(n541) );
  XNOR2_X1 U634 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U635 ( .A(KEYINPUT84), .B(n696), .ZN(n607) );
  NAND2_X1 U636 ( .A1(n659), .A2(n607), .ZN(n543) );
  NAND2_X1 U637 ( .A1(KEYINPUT82), .A2(n543), .ZN(n544) );
  NOR2_X1 U638 ( .A1(KEYINPUT83), .A2(n544), .ZN(n545) );
  NOR2_X1 U639 ( .A1(KEYINPUT47), .A2(n545), .ZN(n549) );
  NAND2_X1 U640 ( .A1(KEYINPUT82), .A2(n663), .ZN(n547) );
  OR2_X1 U641 ( .A1(n696), .A2(KEYINPUT83), .ZN(n546) );
  NAND2_X1 U642 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U643 ( .A(KEYINPUT48), .B(KEYINPUT70), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n551), .B(n550), .ZN(n559) );
  OR2_X1 U645 ( .A1(n552), .A2(n672), .ZN(n553) );
  XNOR2_X1 U646 ( .A(KEYINPUT109), .B(n553), .ZN(n754) );
  NOR2_X1 U647 ( .A1(n554), .A2(n576), .ZN(n555) );
  XNOR2_X1 U648 ( .A(n555), .B(KEYINPUT43), .ZN(n557) );
  NOR2_X1 U649 ( .A1(n557), .A2(n556), .ZN(n675) );
  NOR2_X1 U650 ( .A1(n754), .A2(n675), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n559), .A2(n558), .ZN(n743) );
  INV_X1 U652 ( .A(G953), .ZN(n560) );
  NOR2_X1 U653 ( .A1(G898), .A2(n560), .ZN(n737) );
  NAND2_X1 U654 ( .A1(n561), .A2(n737), .ZN(n562) );
  XOR2_X1 U655 ( .A(KEYINPUT92), .B(n562), .Z(n563) );
  NOR2_X1 U656 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U657 ( .A(KEYINPUT93), .B(n565), .ZN(n566) );
  INV_X1 U658 ( .A(n570), .ZN(n571) );
  INV_X1 U659 ( .A(n576), .ZN(n678) );
  NOR2_X1 U660 ( .A1(n678), .A2(n609), .ZN(n572) );
  XNOR2_X2 U661 ( .A(n573), .B(KEYINPUT88), .ZN(n590) );
  INV_X1 U662 ( .A(KEYINPUT75), .ZN(n577) );
  INV_X1 U663 ( .A(KEYINPUT89), .ZN(n579) );
  XNOR2_X1 U664 ( .A(n579), .B(KEYINPUT33), .ZN(n580) );
  INV_X1 U665 ( .A(n605), .ZN(n598) );
  INV_X1 U666 ( .A(n583), .ZN(n584) );
  XNOR2_X2 U667 ( .A(n585), .B(KEYINPUT35), .ZN(n636) );
  NOR2_X1 U668 ( .A1(n586), .A2(n636), .ZN(n589) );
  NOR2_X1 U669 ( .A1(KEYINPUT67), .A2(KEYINPUT44), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n587), .A2(KEYINPUT86), .ZN(n588) );
  INV_X1 U671 ( .A(KEYINPUT67), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n591), .A2(KEYINPUT44), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U675 ( .A1(n595), .A2(n594), .ZN(n617) );
  NOR2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n613) );
  NAND2_X1 U677 ( .A1(n598), .A2(n575), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n600), .A2(n403), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT96), .ZN(n603) );
  INV_X1 U680 ( .A(n684), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n653) );
  NAND2_X1 U682 ( .A1(n351), .A2(n684), .ZN(n688) );
  NOR2_X1 U683 ( .A1(n688), .A2(n605), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT31), .ZN(n671) );
  NAND2_X1 U685 ( .A1(n653), .A2(n671), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n609), .A2(n406), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n357), .A2(n610), .ZN(n650) );
  NAND2_X1 U689 ( .A1(n611), .A2(n650), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n615) );
  OR2_X1 U691 ( .A1(n636), .A2(KEYINPUT86), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n644), .A2(G475), .ZN(n623) );
  XOR2_X1 U694 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n620) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n624), .A2(n640), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(G60) );
  XOR2_X1 U698 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n628) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(n630) );
  INV_X1 U700 ( .A(n640), .ZN(n724) );
  NOR2_X2 U701 ( .A1(n631), .A2(n724), .ZN(n633) );
  XNOR2_X1 U702 ( .A(KEYINPUT56), .B(KEYINPUT120), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(G51) );
  XOR2_X1 U704 ( .A(G125), .B(KEYINPUT37), .Z(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(G27) );
  XOR2_X1 U706 ( .A(n636), .B(G122), .Z(G24) );
  NAND2_X1 U707 ( .A1(n644), .A2(G472), .ZN(n639) );
  XOR2_X1 U708 ( .A(KEYINPUT62), .B(n637), .Z(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U711 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(G57) );
  BUF_X2 U713 ( .A(n644), .Z(n719) );
  NAND2_X1 U714 ( .A1(n719), .A2(G469), .ZN(n648) );
  XOR2_X1 U715 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n646) );
  XOR2_X1 U716 ( .A(n646), .B(n645), .Z(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n649), .A2(n724), .ZN(G54) );
  XNOR2_X1 U719 ( .A(G101), .B(n650), .ZN(G3) );
  NOR2_X1 U720 ( .A1(n667), .A2(n653), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT110), .B(n651), .Z(n652) );
  XNOR2_X1 U722 ( .A(G104), .B(n652), .ZN(G6) );
  NOR2_X1 U723 ( .A1(n672), .A2(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U726 ( .A(G107), .B(n656), .ZN(G9) );
  XNOR2_X1 U727 ( .A(G110), .B(n657), .ZN(G12) );
  XOR2_X1 U728 ( .A(G128), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n661), .B(n660), .ZN(G30) );
  XOR2_X1 U731 ( .A(G143), .B(n662), .Z(G45) );
  NOR2_X1 U732 ( .A1(n667), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U735 ( .A(G146), .B(n666), .ZN(G48) );
  NOR2_X1 U736 ( .A1(n667), .A2(n671), .ZN(n669) );
  XNOR2_X1 U737 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U739 ( .A(G113), .B(n670), .ZN(G15) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n674) );
  XNOR2_X1 U741 ( .A(G116), .B(KEYINPUT115), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(G18) );
  XNOR2_X1 U743 ( .A(G140), .B(n675), .ZN(n676) );
  XNOR2_X1 U744 ( .A(n676), .B(KEYINPUT117), .ZN(G42) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n679), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U748 ( .A(KEYINPUT49), .B(n682), .Z(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U752 ( .A(n689), .B(KEYINPUT118), .ZN(n690) );
  XNOR2_X1 U753 ( .A(KEYINPUT51), .B(n690), .ZN(n691) );
  NOR2_X1 U754 ( .A1(n710), .A2(n691), .ZN(n704) );
  NOR2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n700) );
  INV_X1 U757 ( .A(n696), .ZN(n698) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U760 ( .A(KEYINPUT119), .B(n701), .ZN(n702) );
  AND2_X1 U761 ( .A1(n709), .A2(n702), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U765 ( .A1(n708), .A2(G953), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n383), .A2(n710), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U768 ( .A(n714), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U769 ( .A1(n719), .A2(G478), .ZN(n717) );
  XOR2_X1 U770 ( .A(KEYINPUT122), .B(n715), .Z(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n724), .A2(n718), .ZN(G63) );
  NAND2_X1 U773 ( .A1(n719), .A2(G217), .ZN(n722) );
  XOR2_X1 U774 ( .A(n720), .B(KEYINPUT123), .Z(n721) );
  XNOR2_X1 U775 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(G66) );
  BUF_X1 U777 ( .A(n725), .Z(n726) );
  NOR2_X1 U778 ( .A1(n726), .A2(G953), .ZN(n732) );
  XOR2_X1 U779 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n728) );
  NAND2_X1 U780 ( .A1(G224), .A2(G953), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT124), .B(n729), .ZN(n730) );
  AND2_X1 U783 ( .A1(n730), .A2(G898), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n739) );
  XOR2_X1 U785 ( .A(n734), .B(G101), .Z(n735) );
  XNOR2_X1 U786 ( .A(n733), .B(n735), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U788 ( .A(n739), .B(n738), .Z(n740) );
  XNOR2_X1 U789 ( .A(KEYINPUT126), .B(n740), .ZN(G69) );
  XOR2_X1 U790 ( .A(n741), .B(n742), .Z(n746) );
  XNOR2_X1 U791 ( .A(n743), .B(n746), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n745), .A2(n744), .ZN(n750) );
  XNOR2_X1 U793 ( .A(n746), .B(G227), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U795 ( .A1(G953), .A2(n748), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n750), .A2(n749), .ZN(G72) );
  XNOR2_X1 U797 ( .A(n751), .B(G119), .ZN(G21) );
  XNOR2_X1 U798 ( .A(G131), .B(KEYINPUT127), .ZN(n753) );
  XNOR2_X1 U799 ( .A(n753), .B(n752), .ZN(G33) );
  XOR2_X1 U800 ( .A(G134), .B(n754), .Z(n755) );
  XNOR2_X1 U801 ( .A(KEYINPUT116), .B(n755), .ZN(G36) );
  XOR2_X1 U802 ( .A(G137), .B(n756), .Z(G39) );
endmodule

