//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n465), .A2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  OR2_X1    g054(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n477), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n474), .A2(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n464), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n478), .A2(new_n482), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  INV_X1    g065(.A(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n478), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G136), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n469), .A2(new_n470), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(KEYINPUT68), .A3(G136), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n489), .B1(new_n494), .B2(new_n497), .ZN(G162));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n462), .A2(new_n463), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n500), .A2(new_n468), .A3(new_n471), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n480), .A2(G138), .A3(new_n481), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n503), .B2(new_n495), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  AND2_X1   g084(.A1(G126), .A2(G2105), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n478), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n469), .B2(new_n470), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT69), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  NAND2_X1  g091(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT74), .ZN(new_n524));
  OAI21_X1  g099(.A(G651), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT70), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n519), .A2(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g106(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT6), .B1(KEYINPUT70), .B2(G651), .ZN(new_n533));
  OAI211_X1 g108(.A(G50), .B(G543), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(new_n530), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n536), .A2(new_n537), .A3(G50), .A4(G543), .ZN(new_n538));
  AOI221_X4 g113(.A(new_n526), .B1(new_n531), .B2(G88), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n531), .A2(G88), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT73), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n525), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n546), .B(new_n525), .C1(new_n539), .C2(new_n542), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G303));
  INV_X1    g124(.A(G303), .ZN(G166));
  NAND2_X1  g125(.A1(new_n531), .A2(G89), .ZN(new_n551));
  NAND3_X1  g126(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n554));
  AND2_X1   g129(.A1(G63), .A2(G651), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n553), .A2(new_n554), .B1(new_n521), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n518), .B1(new_n529), .B2(new_n530), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT76), .B(G51), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n551), .A2(new_n556), .A3(new_n559), .ZN(G286));
  INV_X1    g135(.A(G286), .ZN(G168));
  INV_X1    g136(.A(new_n557), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT77), .B(G52), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n521), .A2(new_n536), .ZN(new_n564));
  INV_X1    g139(.A(G90), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n562), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G651), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n566), .A2(new_n569), .ZN(G171));
  AOI22_X1  g145(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n568), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n557), .A2(G43), .ZN(new_n573));
  INV_X1    g148(.A(G81), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  NAND4_X1  g152(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND4_X1  g155(.A1(G319), .A2(G483), .A3(G661), .A4(new_n580), .ZN(G188));
  NAND2_X1  g156(.A1(new_n557), .A2(G53), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT9), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT78), .B(G65), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(new_n584), .B1(G78), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G91), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n585), .A2(new_n568), .B1(new_n564), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  NAND2_X1  g165(.A1(new_n531), .A2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n557), .A2(G49), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n519), .B2(new_n520), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n597), .B2(KEYINPUT79), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  AOI211_X1 g174(.A(new_n599), .B(new_n596), .C1(new_n519), .C2(new_n520), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g176(.A(G48), .B(G543), .C1(new_n532), .C2(new_n533), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n536), .A2(KEYINPUT80), .A3(G48), .A4(G543), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n604), .A2(new_n605), .B1(G86), .B2(new_n531), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n601), .A2(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(new_n521), .ZN(new_n609));
  INV_X1    g184(.A(G60), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n568), .B1(new_n611), .B2(KEYINPUT81), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT81), .B2(new_n611), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n531), .A2(G85), .B1(new_n557), .B2(G47), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n521), .A2(new_n536), .A3(G92), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT10), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n609), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(G54), .B2(new_n557), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n616), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(G168), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n627), .B2(G168), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  OR2_X1    g207(.A1(new_n572), .A2(new_n575), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n627), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n623), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g212(.A1(new_n468), .A2(new_n471), .A3(new_n476), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2100), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n644));
  OR3_X1    g219(.A1(new_n464), .A2(new_n644), .A3(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n464), .B2(G111), .ZN(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n645), .A2(new_n646), .A3(G2104), .A4(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n487), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n649), .A2(G123), .B1(G135), .B2(new_n496), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n642), .A2(new_n643), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n673), .B2(new_n670), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT86), .Z(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT87), .B(KEYINPUT88), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1981), .B(G1986), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n695), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G35), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G162), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT29), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G2090), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  NOR2_X1   g282(.A1(G4), .A2(G16), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n624), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1348), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT27), .B(G1996), .Z(new_n712));
  NOR2_X1   g287(.A1(G29), .A2(G32), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  INV_X1    g290(.A(G129), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n487), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n476), .A2(G105), .ZN(new_n718));
  INV_X1    g293(.A(G141), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n492), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT99), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n713), .B1(new_n723), .B2(G29), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n707), .B(new_n711), .C1(new_n712), .C2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n702), .A2(G33), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT25), .ZN(new_n728));
  INV_X1    g303(.A(G139), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n492), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n468), .A2(new_n471), .A3(G127), .ZN(new_n732));
  INV_X1    g307(.A(G115), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n475), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n735), .A2(new_n482), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n726), .B1(new_n738), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2072), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n706), .B2(KEYINPUT103), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n743), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n576), .B2(new_n743), .ZN(new_n747));
  OAI22_X1  g322(.A1(G1961), .A2(new_n745), .B1(new_n747), .B2(G1341), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n724), .B2(new_n712), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n702), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G160), .B2(new_n702), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT97), .B(G2084), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G27), .A2(G29), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G164), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G1341), .B2(new_n747), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n749), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n743), .A2(G21), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G286), .B2(G16), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT100), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n651), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT30), .B(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(new_n702), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n745), .A2(G1961), .B1(new_n764), .B2(new_n763), .ZN(new_n775));
  AND4_X1   g350(.A1(new_n766), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT102), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n725), .A2(new_n742), .A3(new_n761), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n705), .A2(G2090), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n743), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT104), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT23), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1956), .ZN(new_n785));
  AOI21_X1  g360(.A(KEYINPUT105), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n777), .B2(new_n776), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n702), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n649), .A2(G128), .B1(G140), .B2(new_n496), .ZN(new_n790));
  OAI221_X1 g365(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n790), .A2(KEYINPUT93), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n796), .A2(KEYINPUT94), .A3(G29), .ZN(new_n797));
  AOI21_X1  g372(.A(KEYINPUT94), .B1(new_n796), .B2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n789), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n780), .A2(KEYINPUT105), .A3(new_n785), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n739), .A2(new_n740), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n779), .A2(new_n787), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n743), .A2(G6), .ZN(new_n807));
  INV_X1    g382(.A(G305), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n743), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT91), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  MUX2_X1   g388(.A(G23), .B(G288), .S(G16), .Z(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT92), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n812), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(G16), .A2(G22), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G303), .B2(new_n743), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(G1971), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(G1971), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n649), .A2(G119), .B1(G131), .B2(new_n496), .ZN(new_n827));
  OAI221_X1 g402(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT89), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(G29), .Z(new_n831));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G1991), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n743), .A2(G24), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n743), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT90), .B(G1986), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n826), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n824), .A2(new_n825), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT36), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n826), .A4(new_n840), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n806), .B1(new_n843), .B2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(new_n806), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(new_n624), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n568), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n557), .A2(G55), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n564), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n576), .A2(new_n858), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n572), .A2(new_n575), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n852), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n858), .A2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(G145));
  NAND2_X1  g446(.A1(new_n796), .A2(G164), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n796), .A2(G164), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n640), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n796), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n515), .ZN(new_n877));
  INV_X1    g452(.A(new_n640), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n649), .A2(G130), .B1(G142), .B2(new_n496), .ZN(new_n881));
  OAI221_X1 g456(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n829), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n738), .A2(new_n721), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n738), .B2(new_n723), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n875), .A2(new_n879), .A3(new_n884), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n886), .B2(new_n889), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n651), .B(G160), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NOR3_X1   g473(.A1(new_n545), .A2(new_n548), .A3(new_n808), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G288), .ZN(new_n901));
  AOI21_X1  g476(.A(G305), .B1(new_n544), .B2(new_n547), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n901), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n899), .B2(new_n902), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n904), .A2(new_n906), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n635), .A2(new_n861), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n635), .A2(new_n861), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n623), .A2(G299), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n618), .A2(new_n583), .A3(new_n588), .A4(new_n622), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n915), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n908), .B1(new_n904), .B2(new_n906), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n923), .A2(new_n924), .B1(KEYINPUT108), .B2(new_n921), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n922), .A4(new_n910), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G868), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n858), .A2(G868), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n627), .B1(new_n925), .B2(new_n928), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT109), .B1(new_n935), .B2(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n933), .ZN(G331));
  XNOR2_X1  g513(.A(G171), .B(G168), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n861), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(KEYINPUT110), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n939), .B2(new_n861), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n939), .A2(new_n861), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n913), .A2(new_n914), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(G171), .B(G286), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n862), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n918), .B(new_n919), .C1(new_n950), .C2(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n904), .A2(new_n906), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n951), .A2(new_n948), .B1(new_n904), .B2(new_n906), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT111), .B1(new_n958), .B2(G37), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT43), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n947), .A2(new_n940), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n941), .A2(new_n943), .A3(new_n945), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n920), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n953), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n964), .B(new_n895), .C1(new_n953), .C2(new_n952), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n957), .B2(new_n959), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n515), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n976));
  INV_X1    g551(.A(G2084), .ZN(new_n977));
  XOR2_X1   g552(.A(KEYINPUT112), .B(G40), .Z(new_n978));
  NOR3_X1   g553(.A1(new_n474), .A2(new_n483), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n505), .B2(new_n514), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n976), .A2(new_n977), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n985), .B(G1384), .C1(new_n505), .C2(new_n514), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n472), .A2(new_n473), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n482), .ZN(new_n988));
  INV_X1    g563(.A(new_n483), .ZN(new_n989));
  INV_X1    g564(.A(new_n978), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n984), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n983), .B(G168), .C1(new_n992), .C2(G1966), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G8), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n975), .A2(new_n985), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n979), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n764), .ZN(new_n998));
  AOI21_X1  g573(.A(G168), .B1(new_n998), .B2(new_n983), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n998), .B2(new_n983), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT51), .B1(new_n1002), .B2(KEYINPUT124), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT124), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1008), .A2(new_n977), .B1(new_n997), .B2(new_n764), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n994), .B1(new_n1010), .B2(KEYINPUT51), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n544), .A2(G8), .A3(new_n547), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n544), .A2(KEYINPUT55), .A3(G8), .A4(new_n547), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1008), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n997), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1001), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1008), .A2(new_n1018), .B1(new_n997), .B2(new_n1020), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1015), .B(new_n1016), .C1(new_n1024), .C2(new_n1001), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n601), .A2(new_n606), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n601), .A2(new_n606), .A3(KEYINPUT118), .A4(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n601), .B1(new_n606), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n604), .A2(new_n605), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n531), .A2(G86), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(G1981), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT120), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1032), .A2(new_n1044), .A3(KEYINPUT49), .A4(new_n1038), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n975), .A2(new_n991), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n1001), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1040), .A2(new_n1043), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n591), .A2(G1976), .A3(new_n592), .A4(new_n593), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT116), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT117), .B(G1976), .Z(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1047), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n995), .A2(new_n1059), .A3(new_n979), .A4(new_n996), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n976), .A2(new_n979), .A3(new_n982), .ZN(new_n1061));
  INV_X1    g636(.A(G1961), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1058), .A2(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n992), .A2(KEYINPUT53), .A3(new_n1059), .ZN(new_n1064));
  AOI21_X1  g639(.A(G301), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1026), .A2(new_n1057), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1010), .B(KEYINPUT51), .C1(new_n994), .C2(new_n999), .ZN(new_n1068));
  INV_X1    g643(.A(new_n994), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1003), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1012), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT126), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1002), .A2(G168), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1023), .A2(new_n1048), .A3(new_n1025), .A4(new_n1056), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT63), .B1(new_n1081), .B2(new_n1078), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G288), .A2(G1976), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1048), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1032), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1085), .A2(new_n1047), .B1(new_n1077), .B2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1080), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1012), .A2(new_n1067), .A3(new_n1089), .A4(new_n1072), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT9), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n582), .B(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT121), .B(KEYINPUT57), .C1(new_n1092), .C2(new_n587), .ZN(new_n1093));
  OR2_X1    g668(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g669(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n583), .A2(new_n588), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n995), .A2(new_n979), .A3(new_n996), .A4(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1061), .A2(new_n710), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1046), .A2(new_n800), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n623), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1104), .A2(new_n623), .A3(new_n1105), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1106), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1107), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n979), .A2(new_n980), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1996), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n995), .A2(new_n1119), .A3(new_n979), .A4(new_n996), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(KEYINPUT122), .A3(new_n1115), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n633), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1122), .B(new_n1123), .C1(KEYINPUT123), .C2(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  NOR2_X1   g700(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1110), .A2(new_n1113), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1103), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n623), .A2(KEYINPUT60), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1104), .A2(new_n1105), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1108), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1060), .A2(new_n1058), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1059), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n995), .A2(G160), .A3(new_n996), .A4(new_n1138), .ZN(new_n1139));
  AND4_X1   g714(.A1(G301), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1065), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT125), .B(new_n1135), .C1(new_n1065), .C2(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1081), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1063), .A2(G301), .A3(new_n1064), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1063), .A2(new_n1139), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1135), .B1(new_n1148), .B2(G171), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1068), .A2(new_n1070), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1134), .A2(new_n1145), .A3(new_n1146), .A4(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1074), .A2(new_n1088), .A3(new_n1090), .A4(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n991), .A2(new_n980), .A3(KEYINPUT45), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1119), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n723), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT114), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n796), .B(G2067), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n721), .A2(new_n1119), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n832), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n829), .B(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1153), .ZN(new_n1164));
  AND2_X1   g739(.A1(G290), .A2(G1986), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1153), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT113), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1161), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT115), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1152), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n721), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1153), .B1(new_n1158), .B2(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1155), .A2(KEYINPUT46), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1155), .A2(KEYINPUT46), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT47), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n830), .A2(new_n1162), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1161), .A2(new_n1179), .B1(new_n800), .B2(new_n876), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1153), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1161), .A2(new_n1183), .A3(new_n1164), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1166), .A2(new_n1153), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT48), .Z(new_n1187));
  NOR2_X1   g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1182), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1172), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g765(.A1(G227), .A2(new_n460), .ZN(new_n1192));
  NOR3_X1   g766(.A1(G229), .A2(G401), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g767(.A(new_n1193), .B(new_n897), .C1(new_n970), .C2(new_n971), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


