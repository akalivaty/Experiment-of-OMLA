

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732;

  NOR2_X1 U378 ( .A1(n514), .A2(n513), .ZN(n630) );
  AND2_X4 U379 ( .A1(n592), .A2(n591), .ZN(n692) );
  NAND2_X2 U380 ( .A1(n726), .A2(n622), .ZN(n396) );
  XNOR2_X2 U381 ( .A(n398), .B(n421), .ZN(n726) );
  NOR2_X2 U382 ( .A1(n677), .A2(n520), .ZN(n507) );
  XNOR2_X2 U383 ( .A(n389), .B(n505), .ZN(n677) );
  XNOR2_X2 U384 ( .A(n566), .B(KEYINPUT79), .ZN(n627) );
  NAND2_X1 U385 ( .A1(n586), .A2(n424), .ZN(n592) );
  OR2_X1 U386 ( .A1(n653), .A2(n654), .ZN(n518) );
  XNOR2_X1 U387 ( .A(n393), .B(n392), .ZN(n694) );
  XNOR2_X1 U388 ( .A(n449), .B(n358), .ZN(n392) );
  XNOR2_X1 U389 ( .A(n712), .B(n394), .ZN(n393) );
  XOR2_X1 U390 ( .A(KEYINPUT10), .B(n450), .Z(n712) );
  INV_X2 U391 ( .A(G953), .ZN(n718) );
  XNOR2_X1 U392 ( .A(n558), .B(n466), .ZN(n563) );
  INV_X1 U393 ( .A(n457), .ZN(n407) );
  XNOR2_X1 U394 ( .A(n480), .B(KEYINPUT4), .ZN(n713) );
  XNOR2_X1 U395 ( .A(G146), .B(G125), .ZN(n461) );
  INV_X1 U396 ( .A(KEYINPUT45), .ZN(n420) );
  NOR2_X1 U397 ( .A1(n513), .A2(n508), .ZN(n544) );
  XNOR2_X1 U398 ( .A(n378), .B(KEYINPUT69), .ZN(n377) );
  XOR2_X1 U399 ( .A(KEYINPUT74), .B(KEYINPUT98), .Z(n430) );
  XNOR2_X1 U400 ( .A(G137), .B(KEYINPUT5), .ZN(n429) );
  XNOR2_X1 U401 ( .A(n433), .B(n432), .ZN(n409) );
  XNOR2_X1 U402 ( .A(G137), .B(G140), .ZN(n447) );
  XOR2_X1 U403 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n446) );
  XNOR2_X1 U404 ( .A(n367), .B(n374), .ZN(n402) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n374) );
  NAND2_X1 U406 ( .A1(n375), .A2(n377), .ZN(n367) );
  XNOR2_X1 U407 ( .A(n376), .B(n364), .ZN(n375) );
  XNOR2_X1 U408 ( .A(n713), .B(n411), .ZN(n436) );
  XNOR2_X1 U409 ( .A(n426), .B(n412), .ZN(n411) );
  INV_X1 U410 ( .A(KEYINPUT65), .ZN(n412) );
  XNOR2_X1 U411 ( .A(n428), .B(n427), .ZN(n457) );
  XOR2_X1 U412 ( .A(G113), .B(G119), .Z(n428) );
  XNOR2_X1 U413 ( .A(n479), .B(n478), .ZN(n371) );
  XNOR2_X1 U414 ( .A(n436), .B(n410), .ZN(n464) );
  INV_X1 U415 ( .A(n707), .ZN(n410) );
  INV_X1 U416 ( .A(KEYINPUT95), .ZN(n395) );
  XNOR2_X1 U417 ( .A(n368), .B(n460), .ZN(n418) );
  XNOR2_X1 U418 ( .A(n459), .B(n419), .ZN(n368) );
  INV_X1 U419 ( .A(KEYINPUT18), .ZN(n419) );
  XNOR2_X1 U420 ( .A(n414), .B(n457), .ZN(n705) );
  XNOR2_X1 U421 ( .A(n479), .B(n415), .ZN(n414) );
  XNOR2_X1 U422 ( .A(n416), .B(KEYINPUT16), .ZN(n415) );
  INV_X1 U423 ( .A(KEYINPUT72), .ZN(n416) );
  NAND2_X1 U424 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U425 ( .A(n404), .B(n403), .ZN(n540) );
  INV_X1 U426 ( .A(KEYINPUT39), .ZN(n403) );
  NOR2_X1 U427 ( .A1(n571), .A2(n543), .ZN(n404) );
  NAND2_X1 U428 ( .A1(n573), .A2(n639), .ZN(n558) );
  XNOR2_X1 U429 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n499) );
  NOR2_X1 U430 ( .A1(n694), .A2(G902), .ZN(n455) );
  XNOR2_X1 U431 ( .A(n502), .B(KEYINPUT90), .ZN(n503) );
  XOR2_X1 U432 ( .A(G131), .B(G134), .Z(n437) );
  XNOR2_X1 U433 ( .A(n583), .B(KEYINPUT85), .ZN(n668) );
  NOR2_X1 U434 ( .A1(n401), .A2(n400), .ZN(n399) );
  INV_X1 U435 ( .A(n637), .ZN(n400) );
  XNOR2_X1 U436 ( .A(G122), .B(G140), .ZN(n490) );
  XOR2_X1 U437 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n491) );
  XNOR2_X1 U438 ( .A(G143), .B(G113), .ZN(n488) );
  XOR2_X1 U439 ( .A(G104), .B(G131), .Z(n489) );
  AND2_X1 U440 ( .A1(G227), .A2(n718), .ZN(n425) );
  NOR2_X1 U441 ( .A1(n641), .A2(n388), .ZN(n387) );
  INV_X1 U442 ( .A(n647), .ZN(n372) );
  NOR2_X1 U443 ( .A1(n563), .A2(n471), .ZN(n473) );
  XNOR2_X1 U444 ( .A(n408), .B(n406), .ZN(n607) );
  XNOR2_X1 U445 ( .A(n431), .B(n407), .ZN(n406) );
  XNOR2_X1 U446 ( .A(n436), .B(n409), .ZN(n408) );
  XNOR2_X1 U447 ( .A(G128), .B(G119), .ZN(n443) );
  XNOR2_X1 U448 ( .A(n448), .B(n422), .ZN(n394) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n584) );
  NAND2_X1 U450 ( .A1(n382), .A2(n639), .ZN(n642) );
  NOR2_X1 U451 ( .A1(n538), .A2(n545), .ZN(n405) );
  XNOR2_X1 U452 ( .A(KEYINPUT30), .B(KEYINPUT106), .ZN(n536) );
  XOR2_X1 U453 ( .A(n498), .B(n497), .Z(n514) );
  NOR2_X1 U454 ( .A1(G902), .A2(n601), .ZN(n497) );
  XOR2_X1 U455 ( .A(G104), .B(KEYINPUT75), .Z(n435) );
  XNOR2_X1 U456 ( .A(n477), .B(n371), .ZN(n483) );
  XNOR2_X1 U457 ( .A(n413), .B(n464), .ZN(n685) );
  XNOR2_X1 U458 ( .A(n705), .B(n417), .ZN(n413) );
  XOR2_X1 U459 ( .A(KEYINPUT93), .B(n597), .Z(n697) );
  XNOR2_X1 U460 ( .A(KEYINPUT42), .B(n552), .ZN(n730) );
  NOR2_X1 U461 ( .A1(n577), .A2(n558), .ZN(n559) );
  XNOR2_X1 U462 ( .A(n390), .B(n365), .ZN(n727) );
  XNOR2_X1 U463 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n421) );
  NAND2_X1 U464 ( .A1(n361), .A2(n397), .ZN(n622) );
  AND2_X1 U465 ( .A1(n546), .A2(n548), .ZN(n397) );
  NOR2_X1 U466 ( .A1(n527), .A2(n546), .ZN(n614) );
  AND2_X1 U467 ( .A1(n554), .A2(n524), .ZN(n525) );
  XNOR2_X1 U468 ( .A(KEYINPUT81), .B(n575), .ZN(n357) );
  XNOR2_X1 U469 ( .A(n441), .B(G469), .ZN(n515) );
  XOR2_X1 U470 ( .A(n444), .B(n443), .Z(n358) );
  XOR2_X1 U471 ( .A(G116), .B(G146), .Z(n359) );
  AND2_X1 U472 ( .A1(n728), .A2(n569), .ZN(n360) );
  AND2_X1 U473 ( .A1(n524), .A2(n654), .ZN(n361) );
  AND2_X1 U474 ( .A1(G210), .A2(n465), .ZN(n362) );
  INV_X1 U475 ( .A(n548), .ZN(n651) );
  NAND2_X1 U476 ( .A1(n544), .A2(n372), .ZN(n363) );
  XNOR2_X1 U477 ( .A(KEYINPUT46), .B(KEYINPUT87), .ZN(n364) );
  XOR2_X1 U478 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n365) );
  XNOR2_X1 U479 ( .A(n473), .B(n472), .ZN(n506) );
  XNOR2_X1 U480 ( .A(n602), .B(n603), .ZN(n604) );
  OR2_X2 U481 ( .A1(n506), .A2(n363), .ZN(n500) );
  NAND2_X1 U482 ( .A1(n366), .A2(n668), .ZN(n586) );
  XNOR2_X1 U483 ( .A(n369), .B(KEYINPUT84), .ZN(n366) );
  NOR2_X2 U484 ( .A1(n598), .A2(n697), .ZN(n600) );
  NOR2_X1 U485 ( .A1(n387), .A2(KEYINPUT41), .ZN(n384) );
  NAND2_X1 U486 ( .A1(n383), .A2(n380), .ZN(n676) );
  OR2_X1 U487 ( .A1(n727), .A2(KEYINPUT44), .ZN(n511) );
  NAND2_X1 U488 ( .A1(n685), .A2(n584), .ZN(n379) );
  NOR2_X2 U489 ( .A1(n670), .A2(n584), .ZN(n369) );
  XNOR2_X1 U490 ( .A(n370), .B(n613), .ZN(G57) );
  NOR2_X2 U491 ( .A1(n611), .A2(n697), .ZN(n370) );
  NOR2_X1 U492 ( .A1(n528), .A2(n614), .ZN(n529) );
  NOR2_X2 U493 ( .A1(n604), .A2(n697), .ZN(n606) );
  XNOR2_X1 U494 ( .A(n373), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U495 ( .A1(n688), .A2(n697), .ZN(n373) );
  NAND2_X1 U496 ( .A1(n730), .A2(n732), .ZN(n376) );
  NAND2_X1 U497 ( .A1(n360), .A2(n357), .ZN(n378) );
  XNOR2_X2 U498 ( .A(n379), .B(n362), .ZN(n573) );
  AND2_X1 U499 ( .A1(n387), .A2(KEYINPUT41), .ZN(n381) );
  INV_X1 U500 ( .A(n543), .ZN(n382) );
  NOR2_X1 U501 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U502 ( .A1(n543), .A2(n386), .ZN(n385) );
  INV_X1 U503 ( .A(KEYINPUT41), .ZN(n386) );
  INV_X1 U504 ( .A(n639), .ZN(n388) );
  NOR2_X2 U505 ( .A1(n518), .A2(n554), .ZN(n389) );
  XNOR2_X1 U506 ( .A(n504), .B(KEYINPUT67), .ZN(n653) );
  NAND2_X1 U507 ( .A1(n391), .A2(n509), .ZN(n390) );
  XNOR2_X1 U508 ( .A(n507), .B(KEYINPUT34), .ZN(n391) );
  XNOR2_X1 U509 ( .A(n461), .B(n395), .ZN(n462) );
  XNOR2_X1 U510 ( .A(n396), .B(n503), .ZN(n510) );
  NAND2_X1 U511 ( .A1(n524), .A2(n501), .ZN(n398) );
  XNOR2_X1 U512 ( .A(n463), .B(n418), .ZN(n417) );
  NAND2_X1 U513 ( .A1(n402), .A2(n638), .ZN(n590) );
  NAND2_X1 U514 ( .A1(n402), .A2(n399), .ZN(n583) );
  INV_X1 U515 ( .A(n638), .ZN(n401) );
  NAND2_X1 U516 ( .A1(n405), .A2(n539), .ZN(n571) );
  XNOR2_X2 U517 ( .A(n531), .B(n420), .ZN(n670) );
  XNOR2_X2 U518 ( .A(n500), .B(n499), .ZN(n524) );
  BUF_X1 U519 ( .A(n506), .Z(n520) );
  XNOR2_X2 U520 ( .A(n458), .B(G122), .ZN(n479) );
  XNOR2_X2 U521 ( .A(G116), .B(G107), .ZN(n458) );
  XOR2_X1 U522 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n422) );
  XNOR2_X1 U523 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n423) );
  OR2_X1 U524 ( .A1(n585), .A2(n584), .ZN(n424) );
  XNOR2_X1 U525 ( .A(n437), .B(n359), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n715), .B(n425), .ZN(n439) );
  XNOR2_X1 U527 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U528 ( .A(KEYINPUT92), .ZN(n442) );
  INV_X1 U529 ( .A(n668), .ZN(n716) );
  XNOR2_X1 U530 ( .A(n464), .B(n440), .ZN(n594) );
  INV_X1 U531 ( .A(n570), .ZN(n509) );
  XNOR2_X1 U532 ( .A(n608), .B(KEYINPUT109), .ZN(n609) );
  XNOR2_X1 U533 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U534 ( .A(n610), .B(n609), .ZN(n611) );
  XOR2_X1 U535 ( .A(G101), .B(KEYINPUT66), .Z(n426) );
  XNOR2_X2 U536 ( .A(G143), .B(G128), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n427) );
  XNOR2_X1 U538 ( .A(n430), .B(n429), .ZN(n431) );
  NOR2_X1 U539 ( .A1(G953), .A2(G237), .ZN(n485) );
  NAND2_X1 U540 ( .A1(n485), .A2(G210), .ZN(n432) );
  NOR2_X1 U541 ( .A1(n607), .A2(G902), .ZN(n434) );
  XNOR2_X2 U542 ( .A(G472), .B(n434), .ZN(n548) );
  XOR2_X1 U543 ( .A(n548), .B(KEYINPUT6), .Z(n554) );
  XNOR2_X1 U544 ( .A(G110), .B(n435), .ZN(n707) );
  XNOR2_X1 U545 ( .A(n437), .B(n447), .ZN(n715) );
  XOR2_X1 U546 ( .A(G146), .B(G107), .Z(n438) );
  NOR2_X1 U547 ( .A1(n594), .A2(G902), .ZN(n441) );
  XNOR2_X2 U548 ( .A(n515), .B(KEYINPUT1), .ZN(n654) );
  XNOR2_X1 U549 ( .A(n654), .B(n442), .ZN(n560) );
  XOR2_X1 U550 ( .A(KEYINPUT24), .B(G110), .Z(n444) );
  NAND2_X1 U551 ( .A1(G234), .A2(n718), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n446), .B(n445), .ZN(n476) );
  NAND2_X1 U553 ( .A1(G221), .A2(n476), .ZN(n449) );
  XNOR2_X1 U554 ( .A(n447), .B(KEYINPUT96), .ZN(n448) );
  INV_X1 U555 ( .A(n461), .ZN(n450) );
  XOR2_X1 U556 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n453) );
  NAND2_X1 U557 ( .A1(n584), .A2(G234), .ZN(n451) );
  XNOR2_X1 U558 ( .A(n451), .B(KEYINPUT20), .ZN(n474) );
  NAND2_X1 U559 ( .A1(n474), .A2(G217), .ZN(n452) );
  XNOR2_X1 U560 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X2 U561 ( .A(n455), .B(n454), .ZN(n546) );
  AND2_X1 U562 ( .A1(n560), .A2(n546), .ZN(n456) );
  AND2_X1 U563 ( .A1(n554), .A2(n456), .ZN(n501) );
  INV_X1 U564 ( .A(KEYINPUT19), .ZN(n466) );
  XOR2_X1 U565 ( .A(KEYINPUT77), .B(KEYINPUT94), .Z(n460) );
  NAND2_X1 U566 ( .A1(G224), .A2(n718), .ZN(n459) );
  XNOR2_X1 U567 ( .A(n462), .B(KEYINPUT17), .ZN(n463) );
  OR2_X1 U568 ( .A1(G237), .A2(G902), .ZN(n465) );
  NAND2_X1 U569 ( .A1(G214), .A2(n465), .ZN(n639) );
  XOR2_X1 U570 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n468) );
  NAND2_X1 U571 ( .A1(G234), .A2(G237), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U573 ( .A1(G952), .A2(n469), .ZN(n667) );
  NOR2_X1 U574 ( .A1(G953), .A2(n667), .ZN(n535) );
  NAND2_X1 U575 ( .A1(G902), .A2(n469), .ZN(n532) );
  OR2_X1 U576 ( .A1(n718), .A2(G898), .ZN(n709) );
  NOR2_X1 U577 ( .A1(n532), .A2(n709), .ZN(n470) );
  NOR2_X1 U578 ( .A1(n535), .A2(n470), .ZN(n471) );
  INV_X1 U579 ( .A(KEYINPUT0), .ZN(n472) );
  NAND2_X1 U580 ( .A1(G221), .A2(n474), .ZN(n475) );
  XNOR2_X1 U581 ( .A(KEYINPUT21), .B(n475), .ZN(n647) );
  XOR2_X1 U582 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n478) );
  NAND2_X1 U583 ( .A1(G217), .A2(n476), .ZN(n477) );
  XNOR2_X1 U584 ( .A(G134), .B(KEYINPUT9), .ZN(n481) );
  XNOR2_X1 U585 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U586 ( .A(n483), .B(n482), .ZN(n690) );
  NOR2_X1 U587 ( .A1(G902), .A2(n690), .ZN(n484) );
  XOR2_X1 U588 ( .A(G478), .B(n484), .Z(n513) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(G475), .ZN(n498) );
  XOR2_X1 U590 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n487) );
  NAND2_X1 U591 ( .A1(G214), .A2(n485), .ZN(n486) );
  XNOR2_X1 U592 ( .A(n487), .B(n486), .ZN(n495) );
  XNOR2_X1 U593 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U594 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U595 ( .A(n493), .B(n492), .Z(n494) );
  XNOR2_X1 U596 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n712), .B(n496), .ZN(n601) );
  INV_X1 U598 ( .A(n514), .ZN(n508) );
  NOR2_X1 U599 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n502) );
  NOR2_X1 U600 ( .A1(n546), .A2(n647), .ZN(n504) );
  XNOR2_X1 U601 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n505) );
  NAND2_X1 U602 ( .A1(n513), .A2(n508), .ZN(n570) );
  NAND2_X1 U603 ( .A1(n510), .A2(n727), .ZN(n512) );
  NAND2_X1 U604 ( .A1(n512), .A2(n511), .ZN(n530) );
  AND2_X1 U605 ( .A1(n514), .A2(n513), .ZN(n634) );
  NOR2_X1 U606 ( .A1(n634), .A2(n630), .ZN(n643) );
  NOR2_X1 U607 ( .A1(n653), .A2(n515), .ZN(n539) );
  INV_X1 U608 ( .A(n539), .ZN(n517) );
  OR2_X1 U609 ( .A1(n651), .A2(n520), .ZN(n516) );
  NOR2_X1 U610 ( .A1(n517), .A2(n516), .ZN(n617) );
  NOR2_X1 U611 ( .A1(n518), .A2(n548), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n519), .B(KEYINPUT99), .ZN(n659) );
  NOR2_X1 U613 ( .A1(n520), .A2(n659), .ZN(n522) );
  XOR2_X1 U614 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n521) );
  XNOR2_X1 U615 ( .A(n522), .B(n521), .ZN(n635) );
  NOR2_X1 U616 ( .A1(n617), .A2(n635), .ZN(n523) );
  NOR2_X1 U617 ( .A1(n643), .A2(n523), .ZN(n528) );
  XNOR2_X1 U618 ( .A(n525), .B(KEYINPUT88), .ZN(n526) );
  NAND2_X1 U619 ( .A1(n526), .A2(n654), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n530), .A2(n529), .ZN(n531) );
  OR2_X1 U621 ( .A1(n718), .A2(n532), .ZN(n533) );
  NOR2_X1 U622 ( .A1(G900), .A2(n533), .ZN(n534) );
  NOR2_X1 U623 ( .A1(n535), .A2(n534), .ZN(n545) );
  NAND2_X1 U624 ( .A1(n639), .A2(n651), .ZN(n537) );
  XNOR2_X1 U625 ( .A(n537), .B(n536), .ZN(n538) );
  INV_X1 U626 ( .A(n573), .ZN(n581) );
  XOR2_X1 U627 ( .A(KEYINPUT38), .B(n581), .Z(n543) );
  NAND2_X1 U628 ( .A1(n540), .A2(n634), .ZN(n637) );
  AND2_X1 U629 ( .A1(n540), .A2(n630), .ZN(n542) );
  XNOR2_X1 U630 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n541) );
  XNOR2_X1 U631 ( .A(n542), .B(n541), .ZN(n732) );
  INV_X1 U632 ( .A(n544), .ZN(n641) );
  INV_X1 U633 ( .A(n676), .ZN(n551) );
  NOR2_X1 U634 ( .A1(n647), .A2(n545), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n547), .A2(n546), .ZN(n553) );
  NOR2_X1 U636 ( .A1(n548), .A2(n553), .ZN(n549) );
  XOR2_X1 U637 ( .A(KEYINPUT28), .B(n549), .Z(n550) );
  NOR2_X1 U638 ( .A1(n515), .A2(n550), .ZN(n564) );
  NAND2_X1 U639 ( .A1(n551), .A2(n564), .ZN(n552) );
  INV_X1 U640 ( .A(n553), .ZN(n557) );
  INV_X1 U641 ( .A(n630), .ZN(n555) );
  NOR2_X1 U642 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U643 ( .A1(n557), .A2(n556), .ZN(n577) );
  XNOR2_X1 U644 ( .A(KEYINPUT36), .B(n559), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U646 ( .A(n562), .B(KEYINPUT108), .ZN(n728) );
  INV_X1 U647 ( .A(n563), .ZN(n565) );
  NAND2_X1 U648 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U649 ( .A(n627), .B(KEYINPUT47), .Z(n568) );
  NAND2_X1 U650 ( .A1(n627), .A2(n643), .ZN(n567) );
  NAND2_X1 U651 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U652 ( .A1(KEYINPUT47), .A2(n643), .ZN(n574) );
  NOR2_X1 U653 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n626) );
  NAND2_X1 U655 ( .A1(n574), .A2(n626), .ZN(n575) );
  INV_X1 U656 ( .A(n654), .ZN(n576) );
  NOR2_X1 U657 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n639), .A2(n578), .ZN(n580) );
  XOR2_X1 U659 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n579) );
  XNOR2_X1 U660 ( .A(n580), .B(n579), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n638) );
  INV_X1 U662 ( .A(KEYINPUT2), .ZN(n585) );
  INV_X1 U663 ( .A(n670), .ZN(n698) );
  NAND2_X1 U664 ( .A1(KEYINPUT2), .A2(n637), .ZN(n587) );
  XOR2_X1 U665 ( .A(KEYINPUT80), .B(n587), .Z(n588) );
  NAND2_X1 U666 ( .A1(n698), .A2(n588), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n673) );
  INV_X1 U668 ( .A(n673), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n692), .A2(G469), .ZN(n596) );
  XOR2_X1 U670 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n593) );
  XNOR2_X1 U671 ( .A(n596), .B(n595), .ZN(n598) );
  NOR2_X1 U672 ( .A1(G952), .A2(n718), .ZN(n597) );
  INV_X1 U673 ( .A(KEYINPUT121), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n600), .B(n599), .ZN(G54) );
  XOR2_X1 U675 ( .A(n601), .B(KEYINPUT59), .Z(n603) );
  NAND2_X1 U676 ( .A1(n692), .A2(G475), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT60), .B(KEYINPUT64), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(G60) );
  NAND2_X1 U679 ( .A1(n692), .A2(G472), .ZN(n610) );
  XOR2_X1 U680 ( .A(n607), .B(KEYINPUT62), .Z(n608) );
  XNOR2_X1 U681 ( .A(KEYINPUT63), .B(KEYINPUT110), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT91), .ZN(n613) );
  XOR2_X1 U683 ( .A(G101), .B(n614), .Z(G3) );
  XOR2_X1 U684 ( .A(G104), .B(KEYINPUT111), .Z(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n630), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(G6) );
  XNOR2_X1 U687 ( .A(G107), .B(KEYINPUT112), .ZN(n621) );
  XOR2_X1 U688 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n619) );
  NAND2_X1 U689 ( .A1(n617), .A2(n634), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G9) );
  XNOR2_X1 U692 ( .A(G110), .B(n622), .ZN(G12) );
  XOR2_X1 U693 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n624) );
  NAND2_X1 U694 ( .A1(n627), .A2(n634), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(n625) );
  XOR2_X1 U696 ( .A(G128), .B(n625), .Z(G30) );
  XNOR2_X1 U697 ( .A(G143), .B(n626), .ZN(G45) );
  NAND2_X1 U698 ( .A1(n627), .A2(n630), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(KEYINPUT114), .ZN(n629) );
  XNOR2_X1 U700 ( .A(G146), .B(n629), .ZN(G48) );
  XOR2_X1 U701 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n632) );
  NAND2_X1 U702 ( .A1(n630), .A2(n635), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U704 ( .A(G113), .B(n633), .ZN(G15) );
  NAND2_X1 U705 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n636), .B(G116), .ZN(G18) );
  XNOR2_X1 U707 ( .A(G134), .B(n637), .ZN(G36) );
  XNOR2_X1 U708 ( .A(G140), .B(n638), .ZN(G42) );
  NOR2_X1 U709 ( .A1(n382), .A2(n639), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n645) );
  NOR2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U712 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n677), .A2(n646), .ZN(n664) );
  XOR2_X1 U714 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n649) );
  NAND2_X1 U715 ( .A1(n647), .A2(n546), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(KEYINPUT118), .ZN(n658) );
  XOR2_X1 U719 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n656) );
  NAND2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U723 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U724 ( .A(KEYINPUT51), .B(n661), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n676), .A2(n662), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U727 ( .A(n665), .B(KEYINPUT52), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n667), .A2(n666), .ZN(n682) );
  XOR2_X1 U729 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n669) );
  NAND2_X1 U730 ( .A1(n716), .A2(n669), .ZN(n675) );
  AND2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U732 ( .A(KEYINPUT83), .B(n671), .Z(n672) );
  NOR2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n680) );
  NOR2_X1 U735 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U736 ( .A1(G953), .A2(n678), .ZN(n679) );
  NAND2_X1 U737 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U738 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U739 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n684), .B(n683), .ZN(G75) );
  NAND2_X1 U741 ( .A1(n692), .A2(G210), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n685), .B(n423), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U744 ( .A1(G478), .A2(n692), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n697), .A2(n691), .ZN(G63) );
  NAND2_X1 U747 ( .A1(n692), .A2(G217), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n693), .B(KEYINPUT122), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n697), .A2(n696), .ZN(G66) );
  NAND2_X1 U751 ( .A1(n698), .A2(n718), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n699), .B(KEYINPUT124), .ZN(n704) );
  XOR2_X1 U753 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n701) );
  NAND2_X1 U754 ( .A1(G224), .A2(G953), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n702), .A2(G898), .ZN(n703) );
  NAND2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n711) );
  XOR2_X1 U758 ( .A(n705), .B(G101), .Z(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U761 ( .A(n711), .B(n710), .Z(G69) );
  XOR2_X1 U762 ( .A(n713), .B(n712), .Z(n714) );
  XOR2_X1 U763 ( .A(n715), .B(n714), .Z(n721) );
  XOR2_X1 U764 ( .A(KEYINPUT125), .B(n721), .Z(n717) );
  XNOR2_X1 U765 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U767 ( .A(n720), .B(KEYINPUT126), .ZN(n725) );
  XNOR2_X1 U768 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n723), .A2(G953), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(G72) );
  XNOR2_X1 U772 ( .A(n726), .B(G119), .ZN(G21) );
  XNOR2_X1 U773 ( .A(n727), .B(G122), .ZN(G24) );
  XOR2_X1 U774 ( .A(G125), .B(n728), .Z(n729) );
  XNOR2_X1 U775 ( .A(KEYINPUT37), .B(n729), .ZN(G27) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(n731) );
  XNOR2_X1 U777 ( .A(KEYINPUT127), .B(n731), .ZN(G39) );
  XNOR2_X1 U778 ( .A(G131), .B(n732), .ZN(G33) );
endmodule

