//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT2), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT75), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n208), .A2(new_n209), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G211gat), .B(G218gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT72), .B(G197gat), .ZN(new_n219));
  INV_X1    g018(.A(G204gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n221), .A2(new_n218), .A3(new_n225), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT29), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n217), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n216), .A3(new_n230), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n204), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n240));
  INV_X1    g039(.A(new_n228), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n226), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT73), .A3(new_n228), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n203), .B1(new_n245), .B2(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n233), .A2(new_n236), .A3(new_n217), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT77), .B(new_n217), .C1(new_n229), .C2(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n239), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G22gat), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n202), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT31), .B(G50gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n253), .A2(new_n254), .ZN(new_n260));
  AOI211_X1 g059(.A(G22gat), .B(new_n239), .C1(new_n252), .C2(new_n246), .ZN(new_n261));
  OAI22_X1  g060(.A1(new_n255), .A2(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n253), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G22gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n253), .A2(new_n254), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n202), .A3(new_n265), .A4(new_n258), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G113gat), .B(G120gat), .Z(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n249), .A2(new_n235), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n214), .A2(new_n216), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(KEYINPUT65), .A3(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n275), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n216), .A3(new_n214), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n276), .A2(new_n281), .A3(new_n282), .A4(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n217), .A2(new_n275), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n284), .ZN(new_n290));
  INV_X1    g089(.A(new_n282), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT0), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G85gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  AOI21_X1  g096(.A(new_n283), .B1(new_n217), .B2(KEYINPUT3), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n291), .B1(new_n298), .B2(new_n235), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n278), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n285), .B1(new_n300), .B2(new_n217), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n283), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n288), .A4(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n293), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n293), .A2(new_n303), .ZN(new_n307));
  INV_X1    g106(.A(new_n297), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT6), .ZN(new_n312));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(KEYINPUT24), .ZN(new_n321));
  INV_X1    g120(.A(G169gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(KEYINPUT24), .A3(new_n320), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(KEYINPUT27), .B(G183gat), .Z(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G190gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT64), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT64), .B(KEYINPUT28), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n331), .B2(G190gat), .ZN(new_n336));
  OR3_X1    g135(.A1(new_n324), .A2(new_n317), .A3(KEYINPUT26), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n317), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n334), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n330), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G226gat), .ZN(new_n341));
  INV_X1    g140(.A(G233gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n330), .A2(new_n339), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n345), .A2(new_n343), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n244), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n343), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n348), .B(new_n234), .C1(new_n343), .C2(new_n340), .ZN(new_n349));
  AOI211_X1 g148(.A(KEYINPUT30), .B(new_n316), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n349), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n315), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n316), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n310), .A2(new_n312), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n267), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n345), .A2(new_n278), .A3(new_n280), .ZN(new_n358));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n300), .A2(new_n330), .A3(new_n339), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n366));
  XOR2_X1   g165(.A(G15gat), .B(G43gat), .Z(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT68), .ZN(new_n368));
  XOR2_X1   g167(.A(G71gat), .B(G99gat), .Z(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT66), .B(KEYINPUT33), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n362), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n370), .A2(KEYINPUT69), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n370), .A2(KEYINPUT69), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(new_n371), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n363), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n360), .B1(new_n358), .B2(new_n361), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT34), .ZN(new_n380));
  OR3_X1    g179(.A1(new_n379), .A2(KEYINPUT70), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n379), .B2(KEYINPUT70), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n373), .A2(new_n381), .A3(new_n382), .A4(new_n377), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT36), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT71), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n389), .A3(new_n385), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT36), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(KEYINPUT71), .A3(new_n383), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n357), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n307), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n293), .A2(KEYINPUT81), .A3(new_n303), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n308), .A3(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n398), .A2(new_n355), .A3(new_n351), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n290), .A2(new_n291), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT80), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT39), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n276), .A2(new_n301), .A3(new_n302), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(new_n291), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n402), .A3(new_n291), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(new_n297), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n406), .B2(new_n297), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n405), .B(KEYINPUT40), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT40), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n399), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT82), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n347), .A2(KEYINPUT37), .A3(new_n349), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n316), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(KEYINPUT84), .A3(new_n316), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT83), .B1(new_n352), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n423), .B(KEYINPUT37), .C1(new_n347), .C2(new_n349), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n419), .B(new_n420), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT38), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n316), .B1(new_n347), .B2(new_n349), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n422), .A2(new_n424), .ZN(new_n428));
  INV_X1    g227(.A(new_n344), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n348), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n421), .B1(new_n430), .B2(new_n233), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n348), .A3(new_n245), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT38), .B(new_n315), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n398), .A2(new_n306), .B1(new_n311), .B2(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n426), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n399), .A2(new_n437), .A3(new_n410), .A4(new_n413), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n415), .A2(new_n436), .A3(new_n267), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n390), .A2(new_n392), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT35), .B1(new_n262), .B2(new_n266), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n398), .A2(new_n306), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n312), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n355), .A2(new_n351), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT85), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n354), .A2(KEYINPUT30), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(new_n427), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n350), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n435), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n440), .B(new_n441), .C1(new_n445), .C2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n387), .A2(new_n267), .A3(new_n356), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n394), .A2(new_n439), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT15), .ZN(new_n456));
  INV_X1    g255(.A(G43gat), .ZN(new_n457));
  INV_X1    g256(.A(G50gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G43gat), .A2(G50gat), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n464));
  AOI21_X1  g263(.A(G50gat), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n467));
  AOI21_X1  g266(.A(G43gat), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n456), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT14), .B(G29gat), .ZN(new_n470));
  INV_X1    g269(.A(G36gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n461), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n474), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n470), .B2(new_n471), .ZN(new_n478));
  INV_X1    g277(.A(new_n461), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT17), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n464), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n458), .B1(new_n482), .B2(new_n462), .ZN(new_n483));
  INV_X1    g282(.A(new_n467), .ZN(new_n484));
  NOR2_X1   g283(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n457), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT15), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n487), .B2(new_n478), .ZN(new_n488));
  INV_X1    g287(.A(new_n480), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT17), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n254), .A2(G15gat), .ZN(new_n493));
  INV_X1    g292(.A(G15gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT16), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(G1gat), .B1(new_n493), .B2(new_n495), .ZN(new_n499));
  XOR2_X1   g298(.A(KEYINPUT90), .B(G8gat), .Z(new_n500));
  NOR3_X1   g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n494), .A2(G22gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n254), .A2(G15gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT88), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n499), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n507), .B2(new_n510), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT91), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n498), .A2(new_n499), .A3(new_n509), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n509), .B(new_n496), .C1(new_n503), .C2(new_n504), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G8gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT89), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n502), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n492), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n476), .A2(new_n480), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n514), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n455), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n476), .A2(KEYINPUT17), .A3(new_n480), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n490), .B1(new_n488), .B2(new_n489), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n522), .B1(new_n521), .B2(new_n502), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT91), .B(new_n501), .C1(new_n519), .C2(new_n520), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n514), .A2(new_n525), .B1(G229gat), .B2(G233gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(KEYINPUT18), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n514), .B(new_n525), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n527), .B(KEYINPUT13), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n529), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G197gat), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT11), .B(G169gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT12), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n529), .A2(new_n537), .A3(new_n546), .A4(new_n540), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n541), .A2(KEYINPUT92), .A3(new_n547), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n551), .A2(KEYINPUT93), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT93), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n557));
  OR2_X1    g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(G57gat), .A2(G64gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n558), .B(new_n559), .C1(new_n566), .C2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n563), .A3(new_n557), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G127gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n571), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n556), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n576), .A2(new_n577), .A3(new_n556), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n514), .A2(new_n581), .A3(KEYINPUT95), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT95), .B1(new_n514), .B2(new_n581), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n205), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n584), .A2(new_n586), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n579), .A2(new_n580), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OR3_X1    g389(.A1(new_n576), .A2(new_n556), .A3(new_n577), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n578), .A4(new_n587), .ZN(new_n593));
  AND2_X1   g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(KEYINPUT8), .A3(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G99gat), .B(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n603), .A2(new_n607), .A3(new_n612), .A4(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n532), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n525), .A2(new_n620), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n598), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n597), .A3(new_n624), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n590), .A2(new_n593), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n620), .A2(new_n569), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n567), .A2(new_n563), .A3(new_n557), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n563), .B1(new_n567), .B2(new_n557), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n617), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n613), .A2(new_n638), .A3(new_n615), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n616), .A2(KEYINPUT98), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n636), .A2(new_n637), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n640), .A2(new_n569), .A3(new_n617), .A4(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT99), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n632), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  INV_X1    g446(.A(new_n632), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n638), .B1(new_n613), .B2(new_n615), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n637), .B1(new_n650), .B2(new_n639), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n642), .A2(KEYINPUT99), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n647), .B(new_n648), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n620), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n646), .B1(new_n655), .B2(new_n645), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  OAI21_X1  g458(.A(new_n631), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n645), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n653), .B2(new_n654), .ZN(new_n663));
  OAI211_X1 g462(.A(KEYINPUT101), .B(new_n661), .C1(new_n663), .C2(new_n646), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n662), .ZN(new_n666));
  INV_X1    g465(.A(new_n654), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n644), .B2(new_n647), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n666), .B(new_n659), .C1(new_n668), .C2(new_n662), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n645), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n672), .A2(KEYINPUT100), .A3(new_n666), .A4(new_n659), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n660), .A2(new_n664), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n630), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n454), .A2(new_n555), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n310), .A2(new_n312), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT102), .B(G1gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND4_X1  g481(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n448), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n448), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  OAI221_X1 g485(.A(new_n683), .B1(new_n508), .B2(new_n685), .C1(new_n686), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g486(.A(new_n676), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n388), .A2(new_n393), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n676), .A2(new_n494), .A3(new_n440), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n454), .A2(new_n555), .ZN(new_n693));
  INV_X1    g492(.A(new_n267), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n675), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT104), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  OAI21_X1  g500(.A(new_n666), .B1(new_n668), .B2(new_n662), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT101), .B1(new_n702), .B2(new_n661), .ZN(new_n703));
  INV_X1    g502(.A(new_n664), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT100), .B1(new_n656), .B2(new_n659), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n663), .A2(new_n670), .A3(new_n646), .A4(new_n661), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n590), .A2(new_n593), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n627), .A2(new_n629), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n693), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n473), .A3(new_n678), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n394), .A2(new_n439), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n451), .A2(new_n453), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n709), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(KEYINPUT44), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n454), .B2(new_n709), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n551), .A2(new_n552), .ZN(new_n722));
  INV_X1    g521(.A(new_n708), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n674), .ZN(new_n724));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724), .B2(new_n677), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n713), .A2(new_n725), .ZN(G1328gat));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n471), .A3(new_n448), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT46), .Z(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n724), .B2(new_n444), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1329gat));
  NAND2_X1  g529(.A1(new_n463), .A2(new_n464), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n724), .B2(new_n689), .ZN(new_n732));
  INV_X1    g531(.A(new_n440), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n731), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n711), .A2(new_n734), .B1(KEYINPUT105), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n737), .B(new_n738), .Z(G1330gat));
  OAI22_X1  g538(.A1(new_n724), .A2(new_n267), .B1(new_n485), .B2(new_n484), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT48), .B1(new_n740), .B2(KEYINPUT106), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n710), .A2(new_n466), .A3(new_n467), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n695), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n741), .B(new_n743), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n551), .A2(new_n552), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n716), .A2(new_n745), .A3(new_n630), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n707), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n678), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g549(.A1(new_n674), .A2(new_n444), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT49), .B(G64gat), .Z(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n747), .A2(new_n756), .A3(new_n689), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT107), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n747), .B2(new_n733), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT50), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n694), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n722), .A2(new_n708), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n716), .A2(new_n717), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT51), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT108), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n604), .A2(new_n606), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n677), .A2(new_n674), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n767), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n674), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n721), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n771), .B1(new_n776), .B2(new_n677), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(G1336gat));
  NAND4_X1  g577(.A1(new_n718), .A2(new_n720), .A3(new_n448), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  INV_X1    g580(.A(new_n751), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n780), .B(new_n781), .C1(new_n769), .C2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n454), .A2(new_n709), .A3(new_n774), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n768), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n783), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n780), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n786), .B1(new_n793), .B2(KEYINPUT52), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT110), .B(new_n781), .C1(new_n792), .C2(new_n780), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n785), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT111), .B(new_n785), .C1(new_n794), .C2(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1337gat));
  NOR3_X1   g599(.A1(new_n733), .A2(G99gat), .A3(new_n674), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n770), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G99gat), .B1(new_n776), .B2(new_n689), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n776), .B2(new_n267), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OR3_X1    g605(.A1(new_n267), .A2(G106gat), .A3(new_n674), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n805), .B(new_n806), .C1(new_n769), .C2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n267), .A2(G106gat), .A3(new_n674), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n791), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n806), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n813), .B(new_n659), .C1(new_n663), .C2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n668), .B2(new_n662), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n653), .A2(new_n662), .A3(new_n654), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT112), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n814), .B1(new_n655), .B2(new_n645), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n817), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n815), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n671), .A2(new_n673), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT112), .B1(new_n816), .B2(new_n818), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n820), .A3(new_n817), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n659), .B1(new_n663), .B2(new_n814), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT55), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n825), .A2(new_n830), .A3(new_n745), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n527), .B1(new_n535), .B2(new_n526), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n538), .A2(new_n539), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n545), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n550), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n674), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n836), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n707), .A2(KEYINPUT113), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n709), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n829), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n826), .B2(new_n827), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n823), .B(new_n824), .C1(new_n843), .C2(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n717), .A2(new_n838), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n708), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n675), .A2(new_n722), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT114), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851));
  INV_X1    g650(.A(new_n849), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n837), .B(new_n839), .C1(new_n844), .C2(new_n745), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n846), .B1(new_n853), .B2(new_n709), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n851), .B(new_n852), .C1(new_n854), .C2(new_n708), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n850), .A2(new_n678), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n694), .A2(new_n386), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n448), .ZN(new_n859));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n722), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n677), .A2(new_n448), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n733), .A2(new_n694), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n850), .A2(new_n855), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT115), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n553), .A2(new_n554), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(G113gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n860), .B1(new_n864), .B2(new_n866), .ZN(G1340gat));
  NAND3_X1  g666(.A1(new_n864), .A2(G120gat), .A3(new_n707), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n858), .A2(new_n448), .A3(new_n674), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(G120gat), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n868), .B(new_n872), .C1(G120gat), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n864), .A2(G127gat), .A3(new_n708), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n877));
  AOI21_X1  g676(.A(G127gat), .B1(new_n859), .B2(new_n708), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1342gat));
  NOR2_X1   g678(.A1(new_n448), .A2(new_n709), .ZN(new_n880));
  INV_X1    g679(.A(G134gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n858), .A2(new_n882), .B1(new_n883), .B2(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n884), .B(new_n885), .Z(new_n886));
  AND2_X1   g685(.A1(new_n864), .A2(new_n717), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n881), .B2(new_n887), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n707), .A2(new_n838), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n555), .B2(new_n844), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n709), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n847), .B1(new_n891), .B2(KEYINPUT119), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n723), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n852), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n267), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n850), .A2(new_n694), .A3(new_n855), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n895), .A2(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n689), .A2(new_n861), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G141gat), .B1(new_n901), .B2(new_n555), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n267), .B1(new_n388), .B2(new_n393), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT120), .Z(new_n904));
  AND3_X1   g703(.A1(new_n856), .A2(new_n444), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n555), .A2(G141gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT58), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n899), .A2(new_n745), .A3(new_n900), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n909), .A2(G141gat), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1344gat));
  NAND3_X1  g711(.A1(new_n856), .A2(new_n444), .A3(new_n904), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT59), .B1(new_n913), .B2(new_n674), .ZN(new_n914));
  INV_X1    g713(.A(G148gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n900), .A2(KEYINPUT59), .A3(new_n674), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n899), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n674), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT121), .B1(new_n865), .B2(new_n675), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n555), .A2(new_n697), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n846), .B1(new_n890), .B2(new_n709), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n708), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n267), .B1(new_n925), .B2(KEYINPUT122), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(new_n923), .C1(new_n924), .C2(new_n708), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT57), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n850), .A2(new_n855), .A3(new_n897), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n919), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n918), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n918), .A3(new_n935), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1345gat));
  OAI21_X1  g736(.A(G155gat), .B1(new_n901), .B2(new_n723), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n905), .A2(new_n205), .A3(new_n708), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1346gat));
  OAI21_X1  g739(.A(G162gat), .B1(new_n901), .B2(new_n709), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n856), .A2(new_n206), .A3(new_n880), .A4(new_n904), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n678), .A2(new_n444), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n850), .A2(new_n855), .A3(new_n862), .A4(new_n945), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n946), .A2(new_n322), .A3(new_n555), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n850), .A2(new_n855), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n678), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(new_n857), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n448), .A3(new_n722), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n951), .B2(new_n322), .ZN(G1348gat));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n323), .A3(new_n751), .ZN(new_n953));
  OAI21_X1  g752(.A(G176gat), .B1(new_n946), .B2(new_n674), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(G1349gat));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n959));
  OAI21_X1  g758(.A(G183gat), .B1(new_n946), .B2(new_n723), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n950), .A2(new_n448), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n723), .A2(new_n331), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n963), .B(new_n964), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n946), .B2(new_n709), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT61), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n709), .A2(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n961), .B2(new_n968), .ZN(G1351gat));
  AND2_X1   g768(.A1(new_n689), .A2(new_n945), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n929), .B2(new_n930), .ZN(new_n971));
  INV_X1    g770(.A(G197gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(new_n555), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n949), .A2(new_n903), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n974), .A2(new_n444), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n722), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n973), .B1(new_n976), .B2(new_n972), .ZN(G1352gat));
  NOR2_X1   g776(.A1(new_n782), .A2(G204gat), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  OR3_X1    g778(.A1(new_n974), .A2(KEYINPUT62), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n971), .B2(new_n674), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT62), .B1(new_n974), .B2(new_n979), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n975), .A2(new_n223), .A3(new_n708), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n708), .B(new_n970), .C1(new_n929), .C2(new_n930), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n984), .B(new_n990), .C1(new_n986), .C2(new_n987), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1354gat));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n224), .A3(new_n717), .ZN(new_n993));
  OAI21_X1  g792(.A(G218gat), .B1(new_n971), .B2(new_n709), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1355gat));
endmodule


