//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(G58), .A2(G68), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n212), .A2(G50), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n209), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  AOI211_X1 g0023(.A(new_n215), .B(new_n223), .C1(KEYINPUT1), .C2(new_n221), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(G226), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G20), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G33), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  AOI22_X1  g0044(.A1(new_n243), .A2(G77), .B1(G20), .B2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT70), .B1(new_n206), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n253), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT68), .B(G1), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n241), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n244), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT11), .B1(new_n249), .B2(new_n255), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT68), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT68), .A2(G1), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n263), .A2(G13), .A3(G20), .A4(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G68), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT12), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n261), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT14), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n252), .B1(G33), .B2(G41), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g0074(.A(KEYINPUT69), .B(G1698), .Z(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G226), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G232), .A2(G1698), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G97), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n250), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n271), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(G1), .B(G13), .C1(new_n250), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G41), .A2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n283), .A2(new_n284), .A3(G274), .A4(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT68), .A2(G1), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT68), .A2(G1), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n271), .B1(new_n291), .B2(new_n286), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n288), .B1(G238), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n281), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n281), .B2(new_n293), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n270), .B(G169), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n294), .B(KEYINPUT13), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n270), .B1(new_n300), .B2(G169), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n269), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G200), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(new_n268), .C1(new_n305), .C2(new_n300), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n274), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n241), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  OR2_X1    g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n309), .B1(new_n312), .B2(G20), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n241), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(G68), .B(new_n308), .C1(new_n315), .C2(KEYINPUT76), .ZN(new_n316));
  INV_X1    g0116(.A(G58), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n244), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(new_n211), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(G20), .B1(G159), .B2(new_n247), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT16), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n312), .A2(new_n309), .A3(G20), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n274), .B2(new_n241), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT16), .A3(new_n320), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(new_n255), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n329));
  XOR2_X1   g0129(.A(new_n329), .B(KEYINPUT8), .Z(new_n330));
  NAND2_X1  g0130(.A1(new_n260), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n265), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n323), .A2(new_n328), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT80), .ZN(new_n335));
  OAI211_X1 g0135(.A(G232), .B(new_n283), .C1(new_n257), .C2(new_n285), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT78), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n287), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n337), .B1(new_n336), .B2(new_n287), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT79), .A2(G190), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT79), .A2(G190), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n312), .A2(G226), .A3(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OR2_X1    g0148(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n272), .C2(new_n273), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n271), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT77), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n355), .A3(new_n271), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n345), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n340), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n358), .A3(new_n338), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n334), .A2(new_n335), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT17), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n334), .A2(new_n335), .A3(new_n362), .A4(KEYINPUT17), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n352), .A2(new_n355), .A3(new_n271), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n355), .B1(new_n352), .B2(new_n271), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n339), .A2(new_n340), .A3(G179), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n369), .A2(new_n370), .B1(new_n371), .B2(new_n359), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n331), .A2(new_n333), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT16), .B1(new_n316), .B2(new_n320), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n327), .A2(new_n255), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT18), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n365), .A2(new_n366), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n275), .A2(G232), .A3(new_n312), .ZN(new_n382));
  INV_X1    g0182(.A(G1698), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n310), .B2(new_n311), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G238), .ZN(new_n385));
  INV_X1    g0185(.A(G107), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n382), .B(new_n385), .C1(new_n386), .C2(new_n312), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n271), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n288), .B1(G244), .B2(new_n292), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n305), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT8), .B(G58), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n392), .A2(new_n248), .B1(new_n241), .B2(new_n203), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n242), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n255), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT73), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n265), .A2(G77), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n259), .B2(G77), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n391), .B(new_n400), .C1(G200), .C2(new_n390), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n371), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n388), .A2(new_n299), .A3(new_n389), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR4_X1   g0205(.A1(new_n307), .A2(new_n381), .A3(new_n401), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n265), .A2(new_n246), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n259), .B2(new_n246), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT72), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n330), .A2(new_n243), .ZN(new_n411));
  INV_X1    g0211(.A(G150), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n411), .B1(new_n412), .B2(new_n248), .C1(new_n241), .C2(new_n202), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n255), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(KEYINPUT9), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n312), .B1(new_n348), .B2(new_n383), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n349), .A2(G222), .A3(new_n350), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n271), .B1(G77), .B2(new_n312), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n292), .A2(G226), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n418), .A2(new_n419), .A3(new_n287), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G190), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT9), .B1(new_n410), .B2(new_n414), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n407), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n410), .A2(new_n414), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n427), .A2(KEYINPUT75), .A3(new_n415), .A4(new_n421), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n420), .A2(new_n360), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT10), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n422), .A2(new_n423), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT74), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n429), .A2(KEYINPUT10), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n427), .A2(new_n415), .A3(new_n421), .A4(new_n435), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT74), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n425), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n420), .A2(new_n299), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G169), .B2(new_n420), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n406), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT5), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G41), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(G41), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n263), .A2(new_n449), .A3(G45), .A4(new_n264), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT83), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n283), .A2(G274), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n447), .B2(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n291), .A2(KEYINPUT83), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n312), .A2(G257), .A3(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G294), .ZN(new_n459));
  INV_X1    g0259(.A(G250), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n351), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n271), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT93), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n271), .B1(new_n452), .B2(new_n456), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(G264), .ZN(new_n465));
  OAI21_X1  g0265(.A(G45), .B1(new_n282), .B2(KEYINPUT5), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n451), .B1(new_n257), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n448), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n456), .A3(new_n468), .ZN(new_n469));
  AND4_X1   g0269(.A1(new_n463), .A2(new_n469), .A3(G264), .A4(new_n283), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n457), .B(new_n462), .C1(new_n465), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n461), .A2(new_n271), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(G264), .A3(new_n283), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT93), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n469), .A2(new_n463), .A3(G264), .A4(new_n283), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G190), .A3(new_n457), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n241), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n386), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(G20), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(KEYINPUT88), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n241), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(KEYINPUT88), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n488), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n312), .A2(new_n241), .A3(G87), .A4(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n484), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n493), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n255), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT25), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n265), .B2(G107), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT91), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT90), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n291), .A2(G13), .A3(G20), .A4(new_n386), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(new_n497), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT91), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n503), .A3(new_n497), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n332), .A2(KEYINPUT90), .A3(KEYINPUT25), .A4(new_n386), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n499), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n265), .B1(new_n250), .B2(new_n257), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n255), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G107), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n472), .A2(new_n478), .A3(new_n496), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n471), .A2(new_n299), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n371), .B1(new_n477), .B2(new_n457), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g0316(.A(new_n495), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n255), .B1(new_n492), .B2(new_n493), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n516), .B1(new_n519), .B2(new_n510), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n496), .A2(new_n511), .A3(KEYINPUT92), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n512), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT94), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n520), .B(new_n521), .C1(new_n513), .C2(new_n514), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(KEYINPUT94), .A3(new_n512), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G20), .B1(G33), .B2(G283), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT81), .B(G97), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G33), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G20), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n255), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n265), .A2(G116), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n508), .B2(G116), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n371), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n469), .A2(G270), .A3(new_n283), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n274), .A2(G303), .ZN(new_n544));
  OAI211_X1 g0344(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n349), .A2(new_n350), .ZN(new_n546));
  OAI21_X1  g0346(.A(G257), .B1(new_n272), .B2(new_n273), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT86), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n548), .A2(new_n549), .A3(new_n271), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n548), .B2(new_n271), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n457), .B(new_n543), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT21), .B1(new_n542), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n541), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n299), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n542), .A2(new_n552), .A3(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT87), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n542), .A2(new_n552), .A3(new_n559), .A4(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n552), .A2(G200), .ZN(new_n562));
  INV_X1    g0362(.A(new_n554), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n562), .B(new_n563), .C1(new_n343), .C2(new_n552), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n556), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  INV_X1    g0366(.A(G244), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n351), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n384), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n312), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n271), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n469), .A2(G257), .A3(new_n283), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n457), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G169), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n299), .B2(new_n574), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT84), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n279), .A2(KEYINPUT81), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n386), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n386), .A2(KEYINPUT6), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n531), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n279), .A2(new_n386), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G20), .B1(G77), .B2(new_n247), .ZN(new_n591));
  OAI211_X1 g0391(.A(G107), .B(new_n308), .C1(new_n315), .C2(KEYINPUT76), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n255), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n265), .A2(G97), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n508), .B2(G97), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n577), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n254), .A2(new_n252), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n591), .A2(new_n592), .B1(new_n251), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n596), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n599), .A2(KEYINPUT84), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n576), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n599), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n574), .A2(G200), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n305), .C2(new_n574), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n453), .A2(G45), .A3(new_n291), .ZN(new_n606));
  OAI211_X1 g0406(.A(G250), .B(new_n283), .C1(new_n257), .C2(new_n454), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n384), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n275), .A2(G238), .A3(new_n312), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n283), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n360), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n608), .A2(new_n611), .A3(new_n305), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n312), .A2(new_n241), .A3(G68), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n531), .A2(new_n242), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(KEYINPUT19), .ZN(new_n618));
  AOI21_X1  g0418(.A(G20), .B1(new_n280), .B2(KEYINPUT19), .ZN(new_n619));
  NOR2_X1   g0419(.A1(G87), .A2(G107), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n531), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n255), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n332), .A2(new_n394), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(G87), .B2(new_n508), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n394), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n508), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n622), .A2(new_n628), .A3(new_n623), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT85), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n612), .A2(G179), .ZN(new_n631));
  OAI21_X1  g0431(.A(G169), .B1(new_n608), .B2(new_n611), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(KEYINPUT85), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n602), .A2(new_n605), .A3(new_n626), .A4(new_n635), .ZN(new_n636));
  NOR4_X1   g0436(.A1(new_n446), .A2(new_n529), .A3(new_n565), .A4(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n378), .A2(new_n380), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n306), .A2(new_n405), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n303), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n365), .A2(new_n366), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n431), .A2(KEYINPUT10), .B1(new_n436), .B2(new_n438), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n445), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n615), .A2(new_n625), .B1(new_n633), .B2(new_n629), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n602), .A2(new_n512), .A3(new_n605), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n496), .A2(new_n511), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n513), .B2(new_n514), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT95), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n471), .A2(G169), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n299), .B2(new_n471), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n653), .B2(new_n648), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n556), .A2(new_n561), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n635), .A2(new_n626), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n658), .B2(new_n602), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n633), .A2(new_n629), .ZN(new_n660));
  INV_X1    g0460(.A(new_n603), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n576), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n646), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n645), .B1(new_n446), .B2(new_n666), .ZN(G369));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n241), .A2(G13), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n291), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n656), .B(new_n564), .C1(new_n563), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n556), .A2(new_n561), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n554), .A3(new_n675), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n668), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n526), .A2(KEYINPUT94), .A3(new_n512), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT94), .B1(new_n526), .B2(new_n512), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n681), .A2(new_n682), .B1(new_n522), .B2(new_n676), .ZN(new_n683));
  INV_X1    g0483(.A(new_n526), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n675), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n653), .A2(new_n651), .A3(new_n648), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n675), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n675), .B1(new_n556), .B2(new_n561), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n528), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n207), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n531), .A2(new_n533), .A3(new_n620), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(new_n284), .ZN(new_n697));
  INV_X1    g0497(.A(new_n214), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n695), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND3_X1  g0500(.A1(new_n656), .A2(KEYINPUT97), .A3(new_n526), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT97), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n678), .B2(new_n684), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n647), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n663), .B1(new_n658), .B2(new_n602), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT96), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n646), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n662), .A2(KEYINPUT96), .A3(KEYINPUT26), .A4(new_n646), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n660), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n676), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n565), .A2(new_n636), .A3(new_n675), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n528), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n477), .A2(new_n612), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n543), .A2(new_n457), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(G179), .C1(new_n551), .C2(new_n550), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n574), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT30), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n574), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n555), .A2(new_n477), .A3(new_n612), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n612), .A2(G179), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n471), .A2(new_n552), .A3(new_n574), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n675), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n714), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n734), .B(new_n676), .C1(new_n657), .C2(new_n665), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n712), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n700), .B1(new_n737), .B2(G1), .ZN(G364));
  NAND2_X1  g0538(.A1(new_n677), .A2(new_n679), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n284), .B1(new_n669), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n695), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n677), .A2(new_n668), .A3(new_n679), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n740), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT98), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT104), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n252), .B1(G20), .B2(new_n371), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n241), .A2(new_n299), .A3(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n344), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n241), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n754), .A2(G322), .B1(G303), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G20), .A3(new_n305), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n312), .B1(new_n761), .B2(G329), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n758), .B(new_n762), .C1(new_n763), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n752), .A2(new_n305), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n343), .A2(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n769), .A2(G311), .B1(new_n771), .B2(G326), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(G317), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT33), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT33), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n755), .A2(new_n305), .A3(G200), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n772), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT103), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n779), .A2(new_n386), .ZN(new_n783));
  INV_X1    g0583(.A(G87), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n312), .B1(new_n756), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(new_n754), .C2(G58), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n771), .A2(G50), .B1(G97), .B2(new_n765), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n769), .A2(G77), .B1(G68), .B2(new_n773), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT101), .B(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n760), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT102), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n751), .B1(new_n782), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n750), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n694), .A2(new_n274), .ZN(new_n799));
  NAND2_X1  g0599(.A1(G355), .A2(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G355), .A2(KEYINPUT99), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n802), .B1(G116), .B2(new_n207), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n694), .A2(new_n312), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n698), .B2(new_n454), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n454), .B2(new_n236), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n744), .B(new_n794), .C1(new_n798), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n797), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n739), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n748), .A2(new_n749), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n749), .B1(new_n748), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  AOI21_X1  g0617(.A(new_n676), .B1(new_n397), .B2(new_n399), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n404), .B1(new_n401), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n405), .A2(new_n676), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n666), .B2(new_n675), .ZN(new_n822));
  INV_X1    g0622(.A(new_n821), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n676), .B(new_n823), .C1(new_n657), .C2(new_n665), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n743), .B1(new_n825), .B2(new_n733), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n733), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n750), .A2(new_n795), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n744), .B1(new_n203), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n274), .B1(new_n830), .B2(new_n760), .C1(new_n766), .C2(new_n279), .ZN(new_n831));
  INV_X1    g0631(.A(new_n771), .ZN(new_n832));
  INV_X1    g0632(.A(G303), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n832), .A2(new_n833), .B1(new_n386), .B2(new_n756), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n753), .A2(new_n763), .B1(new_n533), .B2(new_n768), .ZN(new_n835));
  INV_X1    g0635(.A(new_n773), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n836), .A2(new_n778), .B1(new_n779), .B2(new_n784), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n312), .B1(new_n839), .B2(new_n760), .C1(new_n766), .C2(new_n317), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n246), .A2(new_n756), .B1(new_n779), .B2(new_n244), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n754), .A2(G143), .B1(G150), .B2(new_n773), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n832), .C1(new_n768), .C2(new_n789), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n840), .B(new_n841), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n838), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n829), .B1(new_n751), .B2(new_n848), .C1(new_n823), .C2(new_n796), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n827), .A2(new_n849), .ZN(G384));
  OR3_X1    g0650(.A1(new_n214), .A2(new_n203), .A3(new_n318), .ZN(new_n851));
  INV_X1    g0651(.A(new_n201), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(G68), .ZN(new_n853));
  AOI211_X1 g0653(.A(G13), .B(new_n291), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT105), .Z(new_n855));
  INV_X1    g0655(.A(KEYINPUT36), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n533), .B(new_n210), .C1(new_n590), .C2(KEYINPUT35), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(KEYINPUT35), .B2(new_n590), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n291), .A2(new_n669), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n268), .A2(new_n676), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n303), .A2(new_n306), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n303), .B2(new_n306), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n824), .B2(new_n820), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n326), .B2(new_n320), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n373), .B1(new_n375), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n359), .A2(new_n371), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n370), .A2(new_n354), .A3(new_n356), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n357), .A2(new_n361), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n872), .B(KEYINPUT106), .C1(new_n873), .C2(new_n376), .ZN(new_n874));
  INV_X1    g0674(.A(new_n673), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n334), .A2(new_n362), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT106), .B1(new_n878), .B2(new_n872), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n376), .A2(new_n875), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n878), .A2(new_n377), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n876), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n381), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n334), .A2(new_n362), .B1(new_n372), .B2(new_n869), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n889), .B2(KEYINPUT106), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n878), .A2(new_n872), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n881), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n883), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n886), .B(KEYINPUT38), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n867), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n638), .A2(new_n673), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(KEYINPUT107), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n878), .A2(new_n377), .A3(new_n882), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n883), .ZN(new_n903));
  INV_X1    g0703(.A(new_n381), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n882), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT39), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT107), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n884), .A2(new_n908), .A3(KEYINPUT38), .A4(new_n886), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n896), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n911), .B2(new_n887), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n303), .A2(new_n675), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n898), .B(new_n899), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n446), .B1(new_n712), .B2(new_n735), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n644), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT108), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n675), .C1(new_n720), .C2(new_n726), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n728), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n714), .A2(new_n923), .A3(new_n731), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n823), .B1(new_n864), .B2(new_n865), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n924), .B(new_n926), .C1(new_n911), .C2(new_n887), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n905), .A2(new_n906), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n900), .A2(new_n909), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n730), .B1(new_n713), .B2(new_n528), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n925), .B1(new_n932), .B2(new_n923), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(KEYINPUT40), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n446), .B1(new_n932), .B2(new_n923), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n668), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n861), .B1(new_n919), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n940), .A2(new_n941), .B1(new_n919), .B2(new_n939), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n860), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OAI21_X1  g0744(.A(new_n646), .B1(new_n625), .B2(new_n676), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n660), .A2(new_n625), .A3(new_n676), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n797), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n798), .B1(new_n207), .B2(new_n394), .C1(new_n232), .C2(new_n806), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n743), .ZN(new_n951));
  INV_X1    g0751(.A(new_n779), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n769), .A2(G283), .B1(new_n952), .B2(new_n581), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n763), .B2(new_n836), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n756), .A2(new_n533), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT46), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n274), .B1(new_n774), .B2(new_n760), .C1(new_n766), .C2(new_n386), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n832), .A2(new_n830), .B1(new_n753), .B2(new_n833), .ZN(new_n958));
  NOR4_X1   g0758(.A1(new_n954), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n771), .A2(G143), .B1(G68), .B2(new_n765), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n836), .B2(new_n789), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n312), .B1(new_n753), .B2(new_n412), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n952), .A2(G77), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n852), .B2(new_n768), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n756), .A2(new_n317), .B1(new_n843), .B2(new_n760), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT112), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n959), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT47), .Z(new_n969));
  AOI21_X1  g0769(.A(new_n951), .B1(new_n969), .B2(new_n750), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n949), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT111), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n662), .A2(new_n675), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n602), .A2(new_n605), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n603), .A2(new_n676), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n973), .B1(new_n692), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n691), .B1(new_n681), .B2(new_n682), .ZN(new_n979));
  INV_X1    g0779(.A(new_n690), .ZN(new_n980));
  AND4_X1   g0780(.A1(new_n973), .A2(new_n979), .A3(new_n980), .A4(new_n977), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n972), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n980), .ZN(new_n983));
  INV_X1    g0783(.A(new_n977), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT111), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n692), .A2(new_n973), .A3(new_n977), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT45), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n692), .B2(new_n977), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n982), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n687), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n691), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n683), .A2(new_n685), .A3(new_n995), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n996), .A2(new_n740), .A3(new_n979), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n740), .B1(new_n996), .B2(new_n979), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n736), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n982), .A2(new_n987), .A3(new_n687), .A4(new_n991), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n994), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n737), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n695), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n742), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n687), .A2(new_n984), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT43), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n948), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n977), .A2(new_n684), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n675), .B1(new_n1012), .B2(new_n602), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n528), .A2(new_n691), .A3(new_n977), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1015), .B2(KEYINPUT42), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT42), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1009), .B(new_n1011), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1019), .A3(new_n1010), .A4(new_n948), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1008), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1011), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1009), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n1007), .A3(new_n1021), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n971), .B1(new_n1006), .B2(new_n1028), .ZN(G387));
  AOI211_X1 g0829(.A(G45), .B(new_n696), .C1(G68), .C2(G77), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n392), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n806), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n229), .B2(new_n454), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n799), .A2(new_n696), .B1(new_n386), .B2(new_n694), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT114), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n797), .B(new_n750), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n744), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n330), .A2(new_n773), .B1(G159), .B2(new_n771), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n627), .A2(new_n765), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n244), .C2(new_n768), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n312), .B1(new_n412), .B2(new_n760), .C1(new_n753), .C2(new_n246), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n203), .A2(new_n756), .B1(new_n779), .B2(new_n279), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n757), .A2(G294), .B1(new_n765), .B2(G283), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n771), .A2(G322), .B1(G311), .B2(new_n773), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n833), .B2(new_n768), .C1(new_n774), .C2(new_n753), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n312), .B1(new_n761), .B2(G326), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n533), .B2(new_n779), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1056), .B2(KEYINPUT49), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1047), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1041), .B1(new_n1061), .B2(new_n751), .C1(new_n686), .C2(new_n812), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n695), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1000), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n999), .A2(new_n736), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n999), .A2(new_n741), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n1002), .A2(new_n695), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1000), .B1(new_n994), .B2(new_n1001), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT119), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n994), .A2(new_n1001), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1000), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT119), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n695), .A4(new_n1002), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n994), .A2(new_n742), .A3(new_n1001), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n798), .B1(new_n207), .B2(new_n531), .C1(new_n239), .C2(new_n806), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n743), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n766), .A2(new_n203), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n201), .B2(new_n773), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n392), .B2(new_n768), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT117), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n274), .B1(new_n761), .B2(G143), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n244), .B2(new_n756), .C1(new_n784), .C2(new_n779), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT116), .ZN(new_n1089));
  INV_X1    g0889(.A(G159), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n832), .A2(new_n412), .B1(new_n753), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1086), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT118), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n832), .A2(new_n774), .B1(new_n753), .B2(new_n830), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n312), .B(new_n783), .C1(G322), .C2(new_n761), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n769), .A2(G294), .B1(G303), .B2(new_n773), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n757), .A2(G283), .B1(new_n765), .B2(G116), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1082), .B1(new_n1103), .B2(new_n750), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n812), .B2(new_n977), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1080), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1079), .A2(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n914), .A2(new_n795), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n828), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n743), .B1(new_n330), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n756), .A2(new_n412), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT53), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n771), .A2(G128), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n852), .B2(new_n779), .C1(new_n839), .C2(new_n753), .ZN(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n312), .B1(new_n1116), .B2(new_n760), .C1(new_n836), .C2(new_n843), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n766), .A2(new_n1090), .B1(new_n768), .B2(new_n1118), .ZN(new_n1119));
  OR4_X1    g0919(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n274), .B1(new_n756), .B2(new_n784), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1121), .B(new_n1083), .C1(G107), .C2(new_n773), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n832), .A2(new_n778), .B1(new_n753), .B2(new_n533), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n581), .B2(new_n769), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n779), .A2(new_n244), .B1(new_n763), .B2(new_n760), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT122), .Z(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1111), .B1(new_n1128), .B2(new_n750), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1109), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n915), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n824), .A2(new_n820), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n866), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n915), .B(KEYINPUT120), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n931), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n676), .B(new_n819), .C1(new_n704), .C2(new_n710), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n866), .B1(new_n1137), .B2(new_n820), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1134), .A2(new_n913), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n924), .A2(G330), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n925), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n732), .A2(new_n1133), .A3(G330), .A4(new_n823), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n1136), .B2(new_n1138), .C1(new_n913), .C2(new_n1134), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1130), .B1(new_n1145), .B2(new_n741), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n732), .A2(G330), .A3(new_n823), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n668), .B1(new_n932), .B2(new_n923), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1149), .A2(new_n866), .B1(new_n1150), .B2(new_n926), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1132), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1143), .A2(new_n820), .A3(new_n1137), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1133), .B1(new_n1150), .B2(new_n823), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1151), .A2(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1140), .A2(new_n446), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n917), .A2(new_n1156), .A3(new_n644), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1145), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n695), .B1(new_n1145), .B2(new_n1158), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1147), .B1(new_n1160), .B2(new_n1161), .ZN(G378));
  NAND3_X1  g0962(.A1(new_n1142), .A2(new_n1144), .A3(new_n1155), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1157), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n441), .A2(new_n673), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n440), .B2(new_n445), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n643), .A2(new_n444), .A3(new_n1167), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1166), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n643), .B2(new_n444), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n440), .A2(new_n445), .A3(new_n1168), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1165), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  AND4_X1   g0975(.A1(G330), .A2(new_n929), .A3(new_n934), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n668), .B1(new_n927), .B2(new_n928), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1177), .B2(new_n934), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n916), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n929), .A2(new_n934), .A3(G330), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1175), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n898), .A2(new_n899), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n915), .B1(new_n910), .B2(new_n912), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1177), .A2(new_n934), .A3(new_n1175), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1179), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1164), .A2(new_n1188), .A3(KEYINPUT57), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n695), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT57), .B1(new_n1164), .B2(new_n1188), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1181), .A2(new_n795), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n743), .B1(new_n201), .B2(new_n1110), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n789), .B2(new_n779), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n754), .A2(G128), .B1(G125), .B2(new_n771), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n769), .A2(G137), .B1(G150), .B2(new_n765), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1118), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n757), .A2(new_n1199), .B1(G132), .B2(new_n773), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1196), .B1(new_n1201), .B2(KEYINPUT59), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(KEYINPUT59), .B2(new_n1201), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n754), .A2(G107), .B1(new_n627), .B2(new_n769), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n274), .A2(new_n282), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n760), .A2(new_n778), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G68), .C2(new_n765), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n779), .A2(new_n317), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G116), .B2(new_n771), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n757), .A2(G77), .B1(G97), .B2(new_n773), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1204), .A2(new_n1207), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(G50), .B1(new_n250), .B2(new_n282), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1211), .A2(new_n1212), .B1(new_n1205), .B2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1203), .B(new_n1214), .C1(new_n1212), .C2(new_n1211), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1194), .B1(new_n1215), .B2(new_n750), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1188), .A2(new_n742), .B1(new_n1193), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1192), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT123), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1192), .A2(new_n1220), .A3(new_n1217), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1219), .A2(new_n1221), .ZN(G375));
  NAND2_X1  g1022(.A1(new_n866), .A2(new_n795), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n743), .B1(G68), .B2(new_n1110), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n274), .B(new_n1208), .C1(G128), .C2(new_n761), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n246), .B2(new_n766), .C1(new_n1090), .C2(new_n756), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n769), .A2(G150), .B1(new_n771), .B2(G132), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n843), .B2(new_n753), .C1(new_n836), .C2(new_n1118), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n769), .A2(G107), .B1(new_n771), .B2(G294), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n533), .B2(new_n836), .C1(new_n778), .C2(new_n753), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n757), .A2(G97), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n312), .B1(new_n761), .B2(G303), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n963), .A2(new_n1231), .A3(new_n1232), .A4(new_n1043), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1226), .A2(new_n1228), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1224), .B1(new_n1234), .B2(new_n750), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1155), .A2(new_n742), .B1(new_n1223), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1005), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1236), .B1(new_n1238), .B2(new_n1239), .ZN(G381));
  NAND2_X1  g1040(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n741), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1243), .A2(new_n1244), .B1(new_n949), .B2(new_n970), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1106), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1067), .A2(new_n1069), .A3(new_n816), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(G378), .A2(G381), .A3(G384), .A4(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1241), .A2(new_n1245), .A3(new_n1246), .A4(new_n1248), .ZN(G407));
  INV_X1    g1049(.A(new_n1161), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1146), .B1(new_n1250), .B2(new_n1159), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n674), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1241), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G407), .A2(G213), .A3(new_n1254), .ZN(G409));
  NAND2_X1  g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1247), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1245), .A2(G390), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(new_n1246), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(G387), .A2(new_n1246), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1258), .A2(new_n1263), .A3(new_n1257), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(G387), .B2(new_n1246), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1261), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1067), .A2(new_n1069), .A3(new_n816), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n816), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1245), .B2(G390), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1259), .A2(KEYINPUT125), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(KEYINPUT126), .A4(new_n1263), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1260), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1217), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1164), .A2(new_n1188), .A3(new_n1005), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1217), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1251), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1239), .A2(KEYINPUT60), .A3(new_n1237), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n695), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1239), .B1(KEYINPUT60), .B2(new_n1237), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1236), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(G384), .ZN(new_n1283));
  AND4_X1   g1083(.A1(KEYINPUT62), .A2(new_n1278), .A3(new_n1252), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1274), .A2(new_n1277), .A3(KEYINPUT124), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1286), .A2(new_n1252), .A3(new_n1283), .A4(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1284), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1253), .A2(G2897), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1283), .B(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1253), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1291), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1273), .B1(new_n1290), .B2(new_n1295), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1294), .A2(new_n1283), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1297), .B2(KEYINPUT63), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1288), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1260), .ZN(new_n1301));
  AND3_X1   g1101(.A1(G387), .A2(new_n1246), .A3(new_n1262), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1257), .B1(G387), .B2(new_n1246), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT126), .B1(new_n1304), .B2(new_n1271), .ZN(new_n1305));
  AND4_X1   g1105(.A1(KEYINPUT126), .A2(new_n1270), .A3(new_n1271), .A4(new_n1263), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1301), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1286), .A2(new_n1252), .A3(new_n1287), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1292), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1283), .B(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1298), .A2(new_n1300), .A3(new_n1307), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1296), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1218), .A2(G378), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(G375), .B2(G378), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1283), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1317), .B2(new_n1301), .ZN(new_n1318));
  AOI211_X1 g1118(.A(new_n1283), .B(new_n1260), .C1(new_n1266), .C2(new_n1272), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1315), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1307), .A2(new_n1283), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1314), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1241), .B2(new_n1251), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1273), .A2(new_n1316), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1320), .A2(new_n1325), .ZN(G402));
endmodule


