//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963;
  XOR2_X1   g000(.A(G183gat), .B(G190gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT24), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT23), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n205), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(KEYINPUT25), .C1(G169gat), .C2(new_n214), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n213), .A2(KEYINPUT25), .B1(new_n205), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT27), .B(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n219), .B(KEYINPUT28), .Z(new_n220));
  OAI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  OR3_X1    g021(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n209), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n204), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(KEYINPUT66), .A3(new_n204), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n220), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n234), .B(new_n235), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G227gat), .ZN(new_n239));
  INV_X1    g038(.A(G233gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n236), .A3(new_n231), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT69), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT34), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT34), .B1(new_n244), .B2(KEYINPUT69), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT32), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n242), .B1(new_n238), .B2(new_n243), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT67), .B(KEYINPUT33), .ZN(new_n253));
  XNOR2_X1  g052(.A(G71gat), .B(G99gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT68), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G15gat), .ZN(new_n256));
  INV_X1    g055(.A(G43gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  AOI211_X1 g057(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n252), .B2(new_n253), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n252), .A2(new_n251), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n249), .B(new_n250), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n243), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n241), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT32), .ZN(new_n267));
  INV_X1    g066(.A(new_n253), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n269), .A3(new_n258), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n260), .A2(new_n261), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n249), .B1(new_n272), .B2(new_n250), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT36), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n247), .A2(new_n248), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n249), .A2(new_n279), .A3(new_n270), .A4(new_n271), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT36), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(KEYINPUT36), .C1(new_n264), .C2(new_n273), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288));
  XNOR2_X1  g087(.A(G141gat), .B(G148gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(G155gat), .B2(G162gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G155gat), .B(G162gat), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n236), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n295), .B1(new_n303), .B2(new_n236), .ZN(new_n304));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n287), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n295), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT79), .B(KEYINPUT3), .Z(new_n311));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n237), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n314), .A3(KEYINPUT80), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT80), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n299), .B2(new_n301), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n318), .B2(new_n313), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n309), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n307), .B1(new_n320), .B2(new_n305), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n319), .ZN(new_n322));
  INV_X1    g121(.A(new_n309), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(KEYINPUT5), .A3(new_n305), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327));
  XOR2_X1   g126(.A(G1gat), .B(G29gat), .Z(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G57gat), .B(G85gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT6), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n305), .A3(new_n323), .ZN(new_n334));
  INV_X1    g133(.A(new_n295), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n302), .B2(new_n237), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT5), .B1(new_n336), .B2(new_n305), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n338), .A2(KEYINPUT6), .A3(new_n332), .A4(new_n324), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n232), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n216), .B2(new_n231), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT73), .B(G211gat), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT22), .B1(new_n350), .B2(G218gat), .ZN(new_n351));
  XOR2_X1   g150(.A(G197gat), .B(G204gat), .Z(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OR3_X1    g157(.A1(new_n353), .A2(new_n356), .A3(new_n354), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n349), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n347), .B(new_n360), .C1(new_n346), .C2(new_n348), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n345), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT87), .B1(new_n365), .B2(KEYINPUT37), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT37), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n344), .B(KEYINPUT75), .Z(new_n372));
  AOI211_X1 g171(.A(KEYINPUT38), .B(new_n372), .C1(new_n365), .C2(KEYINPUT37), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n364), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n332), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n321), .B2(new_n325), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n377));
  AOI211_X1 g176(.A(new_n306), .B(new_n309), .C1(new_n315), .C2(new_n319), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n324), .B(new_n332), .C1(new_n378), .C2(new_n307), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n381));
  AOI211_X1 g180(.A(KEYINPUT87), .B(KEYINPUT37), .C1(new_n362), .C2(new_n363), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n345), .B1(new_n367), .B2(new_n369), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT38), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n341), .A2(new_n374), .A3(new_n380), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT31), .B(G50gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n358), .A2(KEYINPUT84), .A3(new_n391), .A4(new_n359), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n392), .A2(new_n317), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n358), .A2(new_n391), .A3(new_n359), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n303), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n312), .A2(new_n391), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n360), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT85), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n317), .A3(new_n392), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n302), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n400), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G22gat), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n355), .B2(new_n357), .ZN(new_n409));
  INV_X1    g208(.A(new_n311), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n298), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n411), .A2(new_n412), .B1(new_n360), .B2(new_n399), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n412), .B2(new_n411), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n398), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n407), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n408), .B1(new_n407), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n390), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n397), .A2(KEYINPUT85), .A3(new_n401), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n405), .B1(new_n404), .B2(new_n400), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(G22gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n408), .A3(new_n415), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n389), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT76), .B(new_n426), .C1(new_n365), .C2(new_n345), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n364), .B2(KEYINPUT30), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n372), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n365), .A2(new_n431), .B1(new_n364), .B2(KEYINPUT30), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n320), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n306), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n336), .B2(new_n305), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n320), .B2(new_n305), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n375), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT86), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT40), .A4(new_n375), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n445), .A2(new_n379), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n433), .A2(new_n442), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n386), .A2(new_n425), .A3(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n416), .A2(new_n417), .A3(new_n390), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n389), .B1(new_n422), .B2(new_n423), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n339), .A2(KEYINPUT82), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n380), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n433), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n286), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n433), .B1(new_n341), .B2(new_n380), .ZN(new_n459));
  INV_X1    g258(.A(new_n273), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n263), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n425), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n379), .A2(new_n377), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n333), .A2(new_n340), .B1(new_n463), .B2(new_n376), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n277), .A2(new_n465), .A3(new_n278), .A4(new_n280), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n464), .A2(new_n466), .A3(new_n433), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n462), .A2(KEYINPUT35), .B1(new_n467), .B2(new_n425), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470));
  INV_X1    g269(.A(G50gat), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT15), .B1(new_n471), .B2(G43gat), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(G43gat), .B2(new_n471), .ZN(new_n473));
  INV_X1    g272(.A(G29gat), .ZN(new_n474));
  INV_X1    g273(.A(G36gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT14), .ZN(new_n476));
  NAND2_X1  g275(.A1(G29gat), .A2(G36gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT91), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(G29gat), .B2(G36gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(G29gat), .A3(G36gat), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n476), .A2(new_n478), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT89), .B(KEYINPUT15), .Z(new_n485));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n471), .B2(G43gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n257), .B2(G50gat), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n486), .A2(new_n471), .A3(G43gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G1gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT16), .ZN(new_n496));
  INV_X1    g295(.A(G15gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G22gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n408), .A2(G15gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(G1gat), .B1(new_n498), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g301(.A(G8gat), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n502), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n494), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n503), .A2(new_n506), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n484), .A2(new_n490), .B1(new_n492), .B2(new_n473), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(KEYINPUT17), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n491), .A2(KEYINPUT17), .A3(new_n493), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n470), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT18), .A3(new_n470), .A4(new_n508), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n509), .A2(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n508), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n470), .B(KEYINPUT13), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n515), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G169gat), .B(G197gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n515), .A2(new_n520), .A3(new_n524), .A4(new_n531), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G155gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G57gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  AND2_X1   g341(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n545), .A2(new_n550), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G64gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(G57gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n541), .A2(G64gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n556), .A2(new_n557), .B1(KEYINPUT92), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT95), .B1(new_n554), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n553), .A2(new_n551), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n548), .B1(new_n546), .B2(new_n549), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n552), .B1(new_n560), .B2(new_n551), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(new_n563), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n580), .A2(G127gat), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n507), .B1(new_n577), .B2(KEYINPUT21), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(G127gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n581), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n540), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(new_n585), .A3(new_n539), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  OAI21_X1  g395(.A(G92gat), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n597), .A2(new_n599), .B1(new_n595), .B2(new_n596), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT8), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(KEYINPUT97), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(KEYINPUT97), .B2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n600), .A2(new_n608), .A3(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n517), .A2(new_n518), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n600), .A2(new_n608), .A3(new_n604), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n608), .B1(new_n600), .B2(new_n604), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n494), .A2(new_n614), .B1(KEYINPUT41), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n594), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n594), .A3(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G134gat), .B(G162gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT96), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n617), .B2(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n618), .A2(KEYINPUT98), .A3(new_n619), .A4(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n592), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G230gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n240), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n566), .A2(new_n576), .B1(new_n607), .B2(new_n609), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n554), .A2(new_n565), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n640), .A2(new_n612), .A3(new_n613), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n638), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n637), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n637), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n639), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n635), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n554), .A2(new_n565), .A3(KEYINPUT95), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n571), .B1(new_n570), .B2(new_n575), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n610), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n607), .B(new_n609), .C1(new_n554), .C2(new_n565), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT10), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n643), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n645), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n646), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n634), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n631), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n469), .A2(new_n535), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n454), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT99), .B(G1gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  INV_X1    g463(.A(new_n661), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n505), .B1(new_n665), .B2(new_n433), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n661), .A2(new_n455), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n661), .B2(new_n286), .ZN(new_n671));
  INV_X1    g470(.A(new_n281), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n497), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n661), .B2(new_n673), .ZN(G1326gat));
  OR3_X1    g473(.A1(new_n661), .A2(KEYINPUT100), .A3(new_n425), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT100), .B1(new_n661), .B2(new_n425), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NOR3_X1   g478(.A1(new_n591), .A2(new_n629), .A3(new_n657), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n469), .A2(new_n535), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n474), .A3(new_n464), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n630), .A2(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n458), .B2(new_n468), .ZN(new_n686));
  INV_X1    g485(.A(new_n535), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n591), .A2(new_n687), .A3(new_n657), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT102), .B1(new_n459), .B2(new_n425), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n451), .A2(new_n456), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n689), .A2(new_n691), .A3(new_n448), .A4(new_n286), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n461), .B1(new_n449), .B2(new_n450), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT35), .B1(new_n693), .B2(new_n456), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n467), .A2(new_n425), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n629), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n686), .B(new_n688), .C1(new_n697), .C2(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n454), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n699), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n475), .A3(new_n433), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n698), .A2(KEYINPUT103), .A3(new_n455), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n698), .B2(new_n455), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G36gat), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n698), .B2(new_n286), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT47), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n681), .A2(new_n257), .A3(new_n672), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n708), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n710), .B(new_n712), .ZN(G1330gat));
  NOR2_X1   g512(.A1(new_n425), .A2(G50gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n681), .A2(new_n714), .B1(KEYINPUT105), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G50gat), .B1(new_n698), .B2(new_n425), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n715), .A2(KEYINPUT105), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1331gat));
  NAND2_X1  g519(.A1(new_n692), .A2(new_n696), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n592), .A2(new_n535), .A3(new_n630), .A4(new_n658), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n464), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT107), .B(G57gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1332gat));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n723), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n455), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n729), .A2(G71gat), .A3(new_n281), .ZN(new_n736));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n286), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n724), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G71gat), .B1(new_n729), .B2(new_n286), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n737), .A3(new_n672), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(KEYINPUT50), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n451), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n591), .A2(new_n535), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n721), .A2(KEYINPUT51), .A3(new_n630), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n721), .A2(new_n630), .A3(new_n747), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n697), .A2(new_n753), .A3(KEYINPUT51), .A4(new_n747), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n749), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n755), .A2(new_n596), .A3(new_n464), .A4(new_n657), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n591), .A2(new_n535), .A3(new_n658), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n686), .B(new_n757), .C1(new_n697), .C2(KEYINPUT44), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n454), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1336gat));
  OAI21_X1  g559(.A(G92gat), .B1(new_n758), .B2(new_n455), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT109), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(G92gat), .C1(new_n758), .C2(new_n455), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n455), .A2(G92gat), .A3(new_n658), .ZN(new_n765));
  INV_X1    g564(.A(new_n748), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT51), .B1(new_n697), .B2(new_n747), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n762), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT52), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n765), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(new_n761), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1337gat));
  NOR3_X1   g573(.A1(new_n281), .A2(G99gat), .A3(new_n658), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G99gat), .B1(new_n758), .B2(new_n286), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1338gat));
  NOR3_X1   g577(.A1(new_n425), .A2(G106gat), .A3(new_n658), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n755), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n755), .A2(KEYINPUT111), .A3(new_n779), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n758), .B2(new_n425), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n779), .B(KEYINPUT110), .Z(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n766), .B2(new_n767), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(G1339gat));
  NAND4_X1  g591(.A1(new_n591), .A2(new_n687), .A3(new_n629), .A4(new_n658), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n470), .B1(new_n519), .B2(new_n508), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n522), .A2(new_n523), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n530), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n627), .A2(new_n534), .A3(new_n628), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n798));
  AOI21_X1  g597(.A(new_n634), .B1(new_n644), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n642), .A2(new_n643), .A3(new_n637), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n656), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n797), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n807));
  INV_X1    g606(.A(new_n798), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n635), .B1(new_n654), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n535), .A3(new_n656), .A4(new_n802), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n534), .A2(new_n796), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n658), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(KEYINPUT113), .A3(new_n657), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n805), .B1(new_n817), .B2(new_n629), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n592), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g619(.A(KEYINPUT114), .B(new_n805), .C1(new_n817), .C2(new_n629), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n793), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n451), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n464), .A3(new_n455), .A4(new_n672), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n687), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  AND2_X1   g626(.A1(new_n822), .A2(new_n464), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT116), .B1(new_n829), .B2(new_n693), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(new_n693), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n433), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(G113gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n535), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n827), .A2(new_n836), .ZN(G1340gat));
  INV_X1    g636(.A(G120gat), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n825), .A2(new_n838), .A3(new_n658), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n657), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n834), .A2(new_n842), .A3(new_n591), .ZN(new_n843));
  OAI21_X1  g642(.A(G127gat), .B1(new_n825), .B2(new_n592), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1342gat));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n833), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n455), .A2(new_n630), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT117), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(G134gat), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n846), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n825), .B2(new_n629), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n852), .A2(KEYINPUT118), .A3(new_n854), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n738), .A2(new_n425), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n829), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n455), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G141gat), .A3(new_n687), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n464), .A2(new_n455), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n738), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n822), .B2(new_n451), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n451), .A2(KEYINPUT57), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n803), .B2(new_n804), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n810), .A2(new_n872), .A3(new_n656), .A4(new_n802), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n535), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n815), .A2(new_n657), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n630), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n592), .B1(new_n876), .B2(new_n805), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n870), .B1(new_n793), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n868), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n687), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n866), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT120), .B(new_n868), .C1(new_n869), .C2(new_n878), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n535), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(KEYINPUT121), .A3(G141gat), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n885), .B2(G141gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n865), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n881), .B1(new_n888), .B2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(new_n864), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n657), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n868), .A2(new_n657), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n793), .B(KEYINPUT122), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n425), .B1(new_n896), .B2(new_n877), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n870), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n822), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n895), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n892), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n894), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n883), .A2(new_n884), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n892), .C1(new_n907), .C2(new_n657), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n893), .B1(new_n906), .B2(new_n908), .ZN(G1345gat));
  AOI21_X1  g708(.A(G155gat), .B1(new_n891), .B2(new_n591), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n591), .A2(G155gat), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT124), .Z(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n907), .B2(new_n912), .ZN(G1346gat));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n630), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G162gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n848), .A2(G162gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n863), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n464), .A2(new_n455), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n672), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT125), .Z(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n824), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n687), .ZN(new_n923));
  NOR4_X1   g722(.A1(new_n823), .A2(new_n464), .A3(new_n455), .A4(new_n693), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n206), .A3(new_n535), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n922), .B2(new_n658), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n207), .A3(new_n657), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n922), .B2(new_n592), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n924), .A2(new_n217), .A3(new_n591), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n924), .A2(new_n218), .A3(new_n630), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n921), .A2(new_n630), .A3(new_n824), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(G190gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G190gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  NAND4_X1  g738(.A1(new_n861), .A2(new_n454), .A3(new_n433), .A4(new_n822), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n535), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n899), .A2(new_n901), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n286), .A2(new_n919), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n535), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n942), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  OAI21_X1  g749(.A(G204gat), .B1(new_n947), .B2(new_n658), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n940), .A2(G204gat), .A3(new_n658), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1353gat));
  OR3_X1    g753(.A1(new_n940), .A2(new_n350), .A3(new_n592), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n943), .A2(new_n591), .A3(new_n945), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  INV_X1    g758(.A(G218gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n940), .B2(new_n629), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n629), .A2(new_n960), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n948), .B2(new_n963), .ZN(G1355gat));
endmodule


