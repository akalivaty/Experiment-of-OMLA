//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(G137), .A3(new_n479), .A4(new_n465), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n465), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT71), .Z(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n483), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(new_n479), .A3(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n468), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n479), .A2(G138), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n478), .A2(new_n465), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n478), .A2(G126), .A3(G2105), .A4(new_n465), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n500), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT72), .B1(new_n500), .B2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(G2104), .B(new_n499), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n497), .A2(new_n504), .ZN(G164));
  XOR2_X1   g080(.A(KEYINPUT5), .B(G543), .Z(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(G88), .B1(new_n512), .B2(G50), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n513), .B1(KEYINPUT73), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n518), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n507), .A2(new_n508), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n506), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n526), .A2(new_n515), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n534), .A2(new_n527), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n514), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n537), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n527), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n506), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n514), .B1(new_n547), .B2(KEYINPUT74), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n510), .A2(G91), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT78), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT79), .B(G65), .Z(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(new_n515), .B1(G78), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n514), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT77), .B1(new_n563), .B2(KEYINPUT76), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n564), .B1(KEYINPUT77), .B2(new_n563), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n527), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n564), .B1(new_n512), .B2(G53), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n558), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND2_X1  g146(.A1(new_n510), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n512), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n535), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n514), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n506), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n514), .B1(new_n585), .B2(KEYINPUT80), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(KEYINPUT80), .B2(new_n585), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n510), .A2(G85), .B1(new_n512), .B2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n526), .A2(G92), .A3(new_n515), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n506), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n512), .B2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n598), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g185(.A1(new_n475), .A2(new_n465), .A3(new_n467), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n489), .A2(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n484), .A2(G123), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n479), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  AND3_X1   g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT82), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  MUX2_X1   g237(.A(new_n662), .B(new_n661), .S(new_n654), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  NOR2_X1   g245(.A1(G6), .A2(G16), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n581), .B2(G16), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT85), .Z(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  NAND2_X1  g249(.A1(G166), .A2(G16), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G16), .B2(G22), .ZN(new_n676));
  INV_X1    g251(.A(G1971), .ZN(new_n677));
  AOI22_X1  g252(.A1(new_n673), .A2(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G23), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT33), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n673), .B2(new_n674), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n679), .A2(KEYINPUT34), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(KEYINPUT34), .B1(new_n679), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(G24), .ZN(new_n689));
  INV_X1    g264(.A(G290), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n680), .ZN(new_n691));
  INV_X1    g266(.A(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT84), .B(G29), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n489), .A2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n484), .A2(G119), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(new_n695), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n687), .A2(new_n688), .A3(new_n693), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT36), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT93), .B(KEYINPUT23), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n680), .A2(G20), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n602), .B2(new_n680), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(G1956), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n694), .A2(G35), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT91), .Z(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n694), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2090), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT94), .Z(new_n720));
  NAND2_X1  g295(.A1(G301), .A2(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n680), .A2(G5), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1961), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G11), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT90), .B(G28), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n725), .B(new_n726), .C1(new_n728), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n680), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n680), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n736), .B1(new_n619), .B2(new_n694), .C1(new_n724), .C2(new_n723), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G34), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n694), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n481), .B2(new_n730), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n732), .B(new_n737), .C1(new_n738), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n717), .A2(new_n718), .ZN(new_n745));
  NOR2_X1   g320(.A1(G164), .A2(new_n694), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G27), .B2(new_n694), .ZN(new_n747));
  INV_X1    g322(.A(G2078), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G19), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n550), .B2(G16), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(new_n750), .B2(G1341), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n743), .A2(new_n738), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT89), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G140), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n484), .A2(G128), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n479), .A2(G116), .ZN(new_n756));
  OAI21_X1  g331(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n754), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n694), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n744), .A2(new_n745), .A3(new_n751), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n730), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n489), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n484), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT26), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AOI22_X1  g347(.A1(G105), .A2(new_n475), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n766), .B1(new_n775), .B2(new_n730), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT27), .Z(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G1996), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n680), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n598), .B2(new_n680), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT86), .B(G1348), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n780), .B(new_n781), .Z(new_n782));
  OAI22_X1  g357(.A1(new_n747), .A2(new_n748), .B1(new_n750), .B2(G1341), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G1996), .B2(new_n777), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n730), .A2(G33), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  AND2_X1   g363(.A1(new_n465), .A2(new_n467), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n789), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n489), .A2(KEYINPUT87), .A3(G139), .ZN(new_n791));
  AOI21_X1  g366(.A(KEYINPUT87), .B1(new_n489), .B2(G139), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n788), .B1(new_n479), .B2(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  OAI21_X1  g369(.A(new_n786), .B1(new_n794), .B2(new_n730), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2072), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n765), .A2(new_n785), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n707), .A2(new_n720), .A3(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  NAND2_X1  g374(.A1(new_n598), .A2(G559), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT38), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(new_n514), .ZN(new_n803));
  INV_X1    g378(.A(G55), .ZN(new_n804));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n804), .A2(new_n527), .B1(new_n535), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT95), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(KEYINPUT95), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n550), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n550), .B(new_n803), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n801), .B(new_n813), .Z(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT96), .B(G860), .Z(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n809), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n817), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n818), .A2(new_n821), .ZN(G145));
  NAND2_X1  g397(.A1(new_n489), .A2(G142), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n484), .A2(G130), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n479), .A2(G118), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n612), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n504), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n498), .A2(KEYINPUT97), .A3(new_n503), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n497), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n758), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n774), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n836));
  INV_X1    g411(.A(new_n494), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n498), .A2(KEYINPUT97), .A3(new_n503), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT97), .B1(new_n498), .B2(new_n503), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n758), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n775), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n794), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n835), .A2(new_n843), .A3(new_n846), .A4(new_n793), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n835), .A2(new_n843), .A3(new_n793), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT98), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n701), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n845), .A2(new_n847), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n849), .A2(KEYINPUT98), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(new_n702), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n829), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n848), .A2(new_n701), .A3(new_n850), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n702), .B1(new_n852), .B2(new_n853), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n856), .A2(new_n857), .A3(new_n828), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n619), .B(new_n481), .ZN(new_n860));
  XOR2_X1   g435(.A(G162), .B(new_n860), .Z(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n855), .A2(new_n863), .A3(new_n858), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT40), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n856), .A2(new_n828), .A3(new_n857), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n828), .B1(new_n856), .B2(new_n857), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n861), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  AND4_X1   g444(.A1(KEYINPUT40), .A2(new_n868), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n865), .A2(new_n870), .ZN(G395));
  XNOR2_X1  g446(.A(new_n813), .B(new_n607), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n602), .A2(new_n598), .ZN(new_n873));
  NAND2_X1  g448(.A1(G299), .A2(new_n597), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n873), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n873), .B2(new_n874), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n876), .B(new_n877), .C1(new_n881), .C2(new_n872), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n877), .B2(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n682), .A2(KEYINPUT100), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g460(.A1(G288), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n884), .B(new_n886), .C1(new_n522), .C2(new_n519), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(G288), .A2(new_n885), .ZN(new_n889));
  OAI21_X1  g464(.A(G166), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(G290), .A2(new_n581), .ZN(new_n892));
  NAND3_X1  g467(.A1(G305), .A2(new_n587), .A3(new_n588), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n887), .A2(new_n890), .A3(new_n892), .A4(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT101), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(KEYINPUT101), .A3(new_n896), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n902), .B2(KEYINPUT42), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n883), .B(new_n903), .Z(new_n904));
  MUX2_X1   g479(.A(new_n809), .B(new_n904), .S(G868), .Z(G295));
  MUX2_X1   g480(.A(new_n809), .B(new_n904), .S(G868), .Z(G331));
  AND3_X1   g481(.A1(new_n811), .A2(new_n812), .A3(G301), .ZN(new_n907));
  AOI21_X1  g482(.A(G301), .B1(new_n811), .B2(new_n812), .ZN(new_n908));
  OAI21_X1  g483(.A(G286), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n813), .A2(G171), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n811), .A2(new_n812), .A3(G301), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(G168), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n875), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n880), .A2(new_n909), .A3(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n902), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(new_n869), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n915), .A2(KEYINPUT103), .B1(new_n913), .B2(new_n875), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n880), .A2(new_n909), .A3(new_n912), .A4(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n901), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n923), .B2(new_n899), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n900), .A2(new_n925), .A3(new_n901), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n917), .B(new_n918), .C1(new_n922), .C2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n914), .A2(new_n915), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n927), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n916), .A2(new_n869), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n928), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n919), .B2(new_n921), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n935), .B2(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT104), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(KEYINPUT43), .C1(new_n935), .C2(new_n931), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n917), .B(new_n918), .C1(new_n929), .C2(new_n927), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n934), .B1(new_n941), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g517(.A(KEYINPUT116), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n841), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n471), .A2(G40), .A3(new_n480), .A4(new_n476), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n945), .B1(new_n497), .B2(new_n504), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n949), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT109), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n946), .B(new_n948), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n841), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n947), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G1971), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n952), .A2(G2090), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(G8), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G8), .ZN(new_n961));
  NOR2_X1   g536(.A1(G166), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT55), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n947), .A2(G2084), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n946), .B(new_n966), .C1(new_n950), .C2(new_n951), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n949), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(KEYINPUT115), .A3(new_n946), .A4(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n841), .B2(new_n945), .ZN(new_n976));
  INV_X1    g551(.A(new_n954), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n945), .B(new_n977), .C1(new_n497), .C2(new_n504), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n948), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n735), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n969), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G286), .A2(new_n961), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n981), .A2(KEYINPUT63), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(G8), .B(new_n963), .C1(new_n958), .C2(new_n959), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n572), .A2(new_n573), .A3(G1976), .A4(new_n574), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT110), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n841), .A2(new_n945), .A3(new_n948), .ZN(new_n988));
  INV_X1    g563(.A(G1976), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(G288), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n987), .A2(G8), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(G8), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n510), .A2(G86), .B1(new_n512), .B2(G48), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n995), .B(new_n996), .C1(new_n514), .C2(new_n579), .ZN(new_n997));
  OAI21_X1  g572(.A(G1981), .B1(new_n578), .B2(new_n580), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT49), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n994), .A2(KEYINPUT112), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n993), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n994), .A2(new_n987), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1003), .A2(new_n1006), .B1(new_n1007), .B2(KEYINPUT52), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n985), .A2(new_n992), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n943), .B1(new_n984), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n981), .A2(KEYINPUT63), .A3(new_n982), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n964), .B2(new_n960), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n985), .A2(new_n992), .A3(new_n1008), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT116), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT63), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n944), .B1(new_n841), .B2(new_n945), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n948), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(new_n1017), .A3(G2090), .ZN(new_n1018));
  OAI21_X1  g593(.A(G8), .B1(new_n1018), .B2(new_n956), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n964), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n985), .A2(new_n1020), .A3(new_n992), .A4(new_n1008), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n981), .A2(new_n982), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1010), .A2(new_n1014), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1008), .A2(new_n992), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n985), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n989), .A3(new_n682), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n997), .B(KEYINPUT113), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT114), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n993), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(KEYINPUT114), .A3(new_n1029), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1024), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT62), .ZN(new_n1035));
  INV_X1    g610(.A(new_n969), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n980), .B1(new_n967), .B2(new_n968), .ZN(new_n1037));
  OAI21_X1  g612(.A(G286), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n969), .A2(new_n975), .A3(G168), .A4(new_n980), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(KEYINPUT51), .A3(G8), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1035), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT124), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT62), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n953), .A2(new_n748), .A3(new_n955), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT126), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT126), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n833), .B2(G1384), .ZN(new_n1060));
  INV_X1    g635(.A(new_n979), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n748), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1060), .A2(new_n1061), .A3(KEYINPUT125), .A4(new_n748), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(KEYINPUT53), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n952), .A2(new_n724), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1058), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1021), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1047), .A2(new_n1051), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n988), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n841), .A2(new_n948), .A3(KEYINPUT120), .A4(new_n945), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G2067), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n952), .A2(new_n781), .ZN(new_n1079));
  AND4_X1   g654(.A1(KEYINPUT60), .A2(new_n1078), .A3(new_n597), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1077), .A2(new_n1076), .B1(new_n952), .B2(new_n781), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n597), .B1(new_n1084), .B2(KEYINPUT60), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1080), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n953), .A2(new_n955), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT119), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n953), .A2(new_n1090), .A3(new_n955), .A4(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(G299), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT118), .B(new_n1095), .C1(new_n558), .C2(new_n568), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT117), .B(G1956), .Z(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1097), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1092), .A2(new_n1097), .A3(KEYINPUT61), .A4(new_n1099), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND3_X1  g683(.A1(new_n1074), .A2(new_n1075), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT121), .B(G1996), .Z(new_n1111));
  NAND3_X1  g686(.A1(new_n953), .A2(new_n955), .A3(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT59), .B(new_n550), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n550), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1086), .A2(new_n1107), .A3(new_n1115), .A4(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1105), .B1(new_n597), .B2(new_n1084), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1100), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT105), .B1(new_n841), .B2(new_n945), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n977), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n841), .A2(KEYINPUT105), .A3(new_n945), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND4_X1   g701(.A1(KEYINPUT53), .A2(new_n953), .A3(new_n748), .A4(new_n948), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1067), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1052), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1056), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(G171), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1058), .A2(new_n1066), .A3(G301), .A4(new_n1067), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT54), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT127), .A4(KEYINPUT54), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1058), .A2(G301), .A3(new_n1067), .A4(new_n1128), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT54), .B1(new_n1069), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1021), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1072), .A2(new_n1122), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1034), .A2(new_n1071), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1126), .A2(new_n947), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n690), .A2(new_n692), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT107), .ZN(new_n1147));
  NAND2_X1  g722(.A1(G290), .A2(G1986), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n758), .B(new_n1077), .ZN(new_n1150));
  INV_X1    g725(.A(G1996), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n774), .B(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n702), .A2(new_n704), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n702), .A2(new_n704), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1145), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1144), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1150), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1145), .B1(new_n774), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1145), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1160), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT46), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1159), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT47), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1166), .A2(new_n1154), .B1(G2067), .B2(new_n758), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1145), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1160), .A2(new_n1146), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(KEYINPUT48), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1145), .A2(new_n1155), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1169), .B2(KEYINPUT48), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1168), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1165), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1157), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g750(.A1(new_n862), .A2(new_n864), .ZN(new_n1177));
  OR2_X1    g751(.A1(G401), .A2(new_n461), .ZN(new_n1178));
  OR3_X1    g752(.A1(G229), .A2(G227), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n1179), .B1(new_n928), .B2(new_n932), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1180), .ZN(G225));
  INV_X1    g755(.A(G225), .ZN(G308));
endmodule


