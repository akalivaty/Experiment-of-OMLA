

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757;

  AND2_X1 U378 ( .A1(n417), .A2(n416), .ZN(n376) );
  INV_X2 U379 ( .A(KEYINPUT71), .ZN(n374) );
  INV_X2 U380 ( .A(G953), .ZN(n749) );
  XNOR2_X2 U381 ( .A(n449), .B(n447), .ZN(n680) );
  NOR2_X2 U382 ( .A1(n756), .A2(n757), .ZN(n567) );
  XNOR2_X2 U383 ( .A(n379), .B(KEYINPUT40), .ZN(n756) );
  XNOR2_X2 U384 ( .A(n378), .B(n377), .ZN(n757) );
  XNOR2_X2 U385 ( .A(n374), .B(G110), .ZN(n373) );
  XNOR2_X2 U386 ( .A(G104), .B(G107), .ZN(n372) );
  XNOR2_X1 U387 ( .A(n432), .B(KEYINPUT22), .ZN(n591) );
  NAND2_X1 U388 ( .A1(n544), .A2(n670), .ZN(n545) );
  XNOR2_X1 U389 ( .A(n626), .B(n625), .ZN(n734) );
  XNOR2_X1 U390 ( .A(n445), .B(KEYINPUT35), .ZN(n754) );
  NAND2_X1 U391 ( .A1(n381), .A2(n384), .ZN(n445) );
  INV_X1 U392 ( .A(n591), .ZN(n396) );
  BUF_X1 U393 ( .A(n561), .Z(n575) );
  XNOR2_X1 U394 ( .A(n443), .B(G128), .ZN(n463) );
  XNOR2_X1 U395 ( .A(KEYINPUT75), .B(KEYINPUT18), .ZN(n406) );
  XNOR2_X1 U396 ( .A(KEYINPUT86), .B(KEYINPUT17), .ZN(n393) );
  INV_X1 U397 ( .A(G143), .ZN(n443) );
  OR2_X1 U398 ( .A1(n747), .A2(n734), .ZN(n660) );
  XNOR2_X2 U399 ( .A(n590), .B(n589), .ZN(n755) );
  XOR2_X2 U400 ( .A(KEYINPUT38), .B(n575), .Z(n683) );
  NOR2_X1 U401 ( .A1(n617), .A2(n616), .ZN(n618) );
  AND2_X1 U402 ( .A1(n620), .A2(KEYINPUT44), .ZN(n621) );
  XNOR2_X1 U403 ( .A(n518), .B(n454), .ZN(n522) );
  XNOR2_X1 U404 ( .A(KEYINPUT4), .B(G131), .ZN(n454) );
  XNOR2_X1 U405 ( .A(n463), .B(n442), .ZN(n518) );
  INV_X1 U406 ( .A(G134), .ZN(n442) );
  INV_X1 U407 ( .A(n611), .ZN(n667) );
  XOR2_X1 U408 ( .A(G140), .B(KEYINPUT11), .Z(n501) );
  XNOR2_X1 U409 ( .A(G131), .B(KEYINPUT98), .ZN(n500) );
  XNOR2_X1 U410 ( .A(G113), .B(G122), .ZN(n503) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(G146), .Z(n520) );
  XNOR2_X1 U412 ( .A(n470), .B(n469), .ZN(n523) );
  INV_X1 U413 ( .A(KEYINPUT88), .ZN(n467) );
  XNOR2_X1 U414 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n485) );
  XNOR2_X1 U415 ( .A(n563), .B(n448), .ZN(n447) );
  INV_X1 U416 ( .A(KEYINPUT108), .ZN(n448) );
  XNOR2_X1 U417 ( .A(n601), .B(n600), .ZN(n692) );
  XNOR2_X1 U418 ( .A(n472), .B(KEYINPUT89), .ZN(n473) );
  XNOR2_X1 U419 ( .A(n544), .B(n358), .ZN(n669) );
  INV_X1 U420 ( .A(KEYINPUT1), .ZN(n462) );
  XNOR2_X1 U421 ( .A(n496), .B(n495), .ZN(n664) );
  XNOR2_X1 U422 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U423 ( .A1(G902), .A2(n724), .ZN(n496) );
  NOR2_X1 U424 ( .A1(n658), .A2(n439), .ZN(n438) );
  INV_X1 U425 ( .A(n657), .ZN(n439) );
  NAND2_X1 U426 ( .A1(n623), .A2(n624), .ZN(n626) );
  NOR2_X1 U427 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U428 ( .A(n517), .B(KEYINPUT9), .ZN(n435) );
  XOR2_X1 U429 ( .A(G107), .B(KEYINPUT7), .Z(n517) );
  XNOR2_X1 U430 ( .A(n522), .B(n362), .ZN(n740) );
  INV_X1 U431 ( .A(KEYINPUT69), .ZN(n458) );
  XOR2_X1 U432 ( .A(G101), .B(G146), .Z(n456) );
  INV_X1 U433 ( .A(n680), .ZN(n371) );
  AND2_X1 U434 ( .A1(n566), .A2(n364), .ZN(n418) );
  AND2_X1 U435 ( .A1(n386), .A2(n385), .ZN(n383) );
  INV_X1 U436 ( .A(n602), .ZN(n385) );
  NAND2_X1 U437 ( .A1(n610), .A2(KEYINPUT34), .ZN(n386) );
  NOR2_X1 U438 ( .A1(n610), .A2(KEYINPUT34), .ZN(n387) );
  XNOR2_X1 U439 ( .A(n588), .B(KEYINPUT101), .ZN(n433) );
  BUF_X1 U440 ( .A(n669), .Z(n408) );
  XNOR2_X1 U441 ( .A(G472), .B(n525), .ZN(n611) );
  XNOR2_X1 U442 ( .A(n423), .B(n422), .ZN(n724) );
  XNOR2_X1 U443 ( .A(n425), .B(n741), .ZN(n423) );
  XNOR2_X1 U444 ( .A(n491), .B(n488), .ZN(n422) );
  XNOR2_X1 U445 ( .A(n487), .B(n426), .ZN(n425) );
  XNOR2_X1 U446 ( .A(KEYINPUT68), .B(G119), .ZN(n465) );
  XNOR2_X1 U447 ( .A(G113), .B(KEYINPUT3), .ZN(n468) );
  XNOR2_X1 U448 ( .A(n562), .B(n450), .ZN(n688) );
  INV_X1 U449 ( .A(KEYINPUT106), .ZN(n450) );
  INV_X1 U450 ( .A(KEYINPUT96), .ZN(n502) );
  XNOR2_X1 U451 ( .A(G143), .B(G104), .ZN(n507) );
  XNOR2_X1 U452 ( .A(n406), .B(n391), .ZN(n390) );
  AND2_X1 U453 ( .A1(n483), .A2(G224), .ZN(n391) );
  INV_X1 U454 ( .A(KEYINPUT104), .ZN(n546) );
  XNOR2_X1 U455 ( .A(n514), .B(n513), .ZN(n560) );
  NOR2_X1 U456 ( .A1(n560), .A2(n559), .ZN(n681) );
  XNOR2_X1 U457 ( .A(n522), .B(n451), .ZN(n632) );
  XNOR2_X1 U458 ( .A(n523), .B(n452), .ZN(n451) );
  XNOR2_X1 U459 ( .A(n521), .B(n363), .ZN(n452) );
  XOR2_X1 U460 ( .A(KEYINPUT16), .B(G122), .Z(n471) );
  XNOR2_X1 U461 ( .A(n490), .B(n424), .ZN(n741) );
  INV_X1 U462 ( .A(KEYINPUT10), .ZN(n424) );
  XNOR2_X1 U463 ( .A(G137), .B(G140), .ZN(n486) );
  XNOR2_X1 U464 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n426) );
  XNOR2_X1 U465 ( .A(G119), .B(G128), .ZN(n481) );
  XOR2_X1 U466 ( .A(KEYINPUT92), .B(G110), .Z(n482) );
  INV_X1 U467 ( .A(KEYINPUT19), .ZN(n431) );
  XNOR2_X1 U468 ( .A(n436), .B(n434), .ZN(n720) );
  XNOR2_X1 U469 ( .A(n518), .B(n359), .ZN(n436) );
  XNOR2_X1 U470 ( .A(n516), .B(n435), .ZN(n434) );
  XNOR2_X1 U471 ( .A(n397), .B(n740), .ZN(n713) );
  INV_X1 U472 ( .A(KEYINPUT42), .ZN(n377) );
  NAND2_X1 U473 ( .A1(n371), .A2(n370), .ZN(n378) );
  INV_X1 U474 ( .A(n564), .ZN(n370) );
  NAND2_X1 U475 ( .A1(n414), .A2(n380), .ZN(n576) );
  AND2_X1 U476 ( .A1(n415), .A2(n421), .ZN(n414) );
  NAND2_X1 U477 ( .A1(n418), .A2(n650), .ZN(n375) );
  AND2_X1 U478 ( .A1(n383), .A2(n382), .ZN(n381) );
  AND2_X1 U479 ( .A1(n356), .A2(n598), .ZN(n394) );
  NOR2_X2 U480 ( .A1(n593), .A2(n667), .ZN(n643) );
  NAND2_X1 U481 ( .A1(n428), .A2(n427), .ZN(n635) );
  INV_X1 U482 ( .A(n606), .ZN(n427) );
  INV_X1 U483 ( .A(KEYINPUT81), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n723), .B(n407), .ZN(n725) );
  XNOR2_X1 U485 ( .A(n724), .B(KEYINPUT122), .ZN(n407) );
  INV_X1 U486 ( .A(KEYINPUT60), .ZN(n401) );
  INV_X1 U487 ( .A(KEYINPUT56), .ZN(n399) );
  NOR2_X1 U488 ( .A1(n577), .A2(n664), .ZN(n356) );
  XOR2_X1 U489 ( .A(n717), .B(n368), .Z(n357) );
  XOR2_X1 U490 ( .A(n462), .B(KEYINPUT64), .Z(n358) );
  XOR2_X1 U491 ( .A(G122), .B(G116), .Z(n359) );
  XOR2_X1 U492 ( .A(n463), .B(KEYINPUT4), .Z(n360) );
  AND2_X1 U493 ( .A1(n419), .A2(n650), .ZN(n361) );
  XNOR2_X1 U494 ( .A(G137), .B(G140), .ZN(n362) );
  AND2_X1 U495 ( .A1(n524), .A2(G210), .ZN(n363) );
  INV_X1 U496 ( .A(n529), .ZN(n650) );
  XOR2_X1 U497 ( .A(KEYINPUT79), .B(KEYINPUT39), .Z(n364) );
  XOR2_X1 U498 ( .A(KEYINPUT48), .B(KEYINPUT66), .Z(n365) );
  XOR2_X1 U499 ( .A(n709), .B(n708), .Z(n366) );
  XOR2_X1 U500 ( .A(n633), .B(KEYINPUT87), .Z(n367) );
  XNOR2_X1 U501 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n368) );
  NOR2_X1 U502 ( .A1(G952), .A2(n749), .ZN(n726) );
  INV_X1 U503 ( .A(n726), .ZN(n403) );
  XOR2_X1 U504 ( .A(n634), .B(KEYINPUT84), .Z(n369) );
  NOR2_X1 U505 ( .A1(n591), .A2(n408), .ZN(n592) );
  NOR2_X1 U506 ( .A1(n605), .A2(n408), .ZN(n430) );
  NAND2_X1 U507 ( .A1(n396), .A2(n394), .ZN(n590) );
  XNOR2_X1 U508 ( .A(n430), .B(n429), .ZN(n428) );
  NOR2_X2 U509 ( .A1(n755), .A2(n643), .ZN(n619) );
  XNOR2_X2 U510 ( .A(n727), .B(n458), .ZN(n464) );
  XNOR2_X2 U511 ( .A(n373), .B(n372), .ZN(n727) );
  NAND2_X1 U512 ( .A1(n376), .A2(n375), .ZN(n379) );
  INV_X1 U513 ( .A(n669), .ZN(n577) );
  NAND2_X1 U514 ( .A1(n669), .A2(n670), .ZN(n607) );
  XNOR2_X2 U515 ( .A(n461), .B(n460), .ZN(n544) );
  INV_X1 U516 ( .A(n418), .ZN(n380) );
  NAND2_X1 U517 ( .A1(n692), .A2(KEYINPUT34), .ZN(n382) );
  NAND2_X1 U518 ( .A1(n388), .A2(n387), .ZN(n384) );
  INV_X1 U519 ( .A(n692), .ZN(n388) );
  XNOR2_X1 U520 ( .A(n389), .B(n360), .ZN(n446) );
  XNOR2_X1 U521 ( .A(n392), .B(n390), .ZN(n389) );
  XNOR2_X1 U522 ( .A(n489), .B(n393), .ZN(n392) );
  XNOR2_X2 U523 ( .A(G146), .B(G125), .ZN(n489) );
  NAND2_X1 U524 ( .A1(n396), .A2(n598), .ZN(n395) );
  XNOR2_X1 U525 ( .A(n395), .B(KEYINPUT80), .ZN(n605) );
  XNOR2_X1 U526 ( .A(n512), .B(n511), .ZN(n717) );
  XNOR2_X1 U527 ( .A(n464), .B(n446), .ZN(n410) );
  NOR2_X1 U528 ( .A1(n607), .A2(n598), .ZN(n601) );
  XNOR2_X1 U529 ( .A(n398), .B(n367), .ZN(n411) );
  XNOR2_X1 U530 ( .A(n413), .B(n459), .ZN(n397) );
  NAND2_X1 U531 ( .A1(n411), .A2(n403), .ZN(n409) );
  NAND2_X1 U532 ( .A1(n688), .A2(n681), .ZN(n449) );
  NAND2_X1 U533 ( .A1(n722), .A2(G472), .ZN(n398) );
  XNOR2_X1 U534 ( .A(n409), .B(n369), .ZN(G57) );
  XNOR2_X1 U535 ( .A(n400), .B(n399), .ZN(G51) );
  NAND2_X1 U536 ( .A1(n405), .A2(n403), .ZN(n400) );
  XNOR2_X1 U537 ( .A(n402), .B(n401), .ZN(G60) );
  NAND2_X1 U538 ( .A1(n404), .A2(n403), .ZN(n402) );
  XNOR2_X1 U539 ( .A(n718), .B(n357), .ZN(n404) );
  XNOR2_X1 U540 ( .A(n710), .B(n366), .ZN(n405) );
  NAND2_X1 U541 ( .A1(n420), .A2(n361), .ZN(n417) );
  XNOR2_X1 U542 ( .A(n536), .B(n431), .ZN(n585) );
  NOR2_X2 U543 ( .A1(n585), .A2(n584), .ZN(n412) );
  XNOR2_X1 U544 ( .A(n410), .B(n728), .ZN(n707) );
  XNOR2_X2 U545 ( .A(n412), .B(n587), .ZN(n608) );
  XNOR2_X1 U546 ( .A(n464), .B(KEYINPUT73), .ZN(n413) );
  NAND2_X1 U547 ( .A1(n420), .A2(n419), .ZN(n415) );
  OR2_X1 U548 ( .A1(n421), .A2(n529), .ZN(n416) );
  XNOR2_X2 U549 ( .A(n553), .B(KEYINPUT72), .ZN(n566) );
  NOR2_X1 U550 ( .A1(n565), .A2(n364), .ZN(n419) );
  INV_X1 U551 ( .A(n566), .ZN(n420) );
  NAND2_X1 U552 ( .A1(n565), .A2(n364), .ZN(n421) );
  NAND2_X1 U553 ( .A1(n635), .A2(n618), .ZN(n622) );
  NAND2_X1 U554 ( .A1(n608), .A2(n433), .ZN(n432) );
  NAND2_X1 U555 ( .A1(n754), .A2(KEYINPUT82), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n441), .B(n365), .ZN(n440) );
  INV_X1 U557 ( .A(n608), .ZN(n610) );
  NOR2_X1 U558 ( .A1(n610), .A2(n437), .ZN(n612) );
  XNOR2_X1 U559 ( .A(n437), .B(n546), .ZN(n552) );
  XNOR2_X2 U560 ( .A(n545), .B(KEYINPUT94), .ZN(n437) );
  NAND2_X1 U561 ( .A1(n440), .A2(n438), .ZN(n747) );
  NAND2_X1 U562 ( .A1(n568), .A2(n569), .ZN(n441) );
  NAND2_X1 U563 ( .A1(n619), .A2(n444), .ZN(n620) );
  XNOR2_X1 U564 ( .A(n713), .B(n453), .ZN(n714) );
  NOR2_X2 U565 ( .A1(G902), .A2(n713), .ZN(n461) );
  XOR2_X1 U566 ( .A(n712), .B(n711), .Z(n453) );
  XNOR2_X1 U567 ( .A(n520), .B(G137), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n599), .B(KEYINPUT102), .ZN(n600) );
  XNOR2_X1 U570 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U571 ( .A(KEYINPUT25), .ZN(n493) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n586), .B(KEYINPUT85), .ZN(n587) );
  INV_X1 U574 ( .A(KEYINPUT63), .ZN(n634) );
  NAND2_X1 U575 ( .A1(G227), .A2(n749), .ZN(n455) );
  XNOR2_X1 U576 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U577 ( .A(n457), .B(KEYINPUT74), .Z(n459) );
  XNOR2_X1 U578 ( .A(KEYINPUT67), .B(G469), .ZN(n460) );
  XOR2_X1 U579 ( .A(G116), .B(G101), .Z(n466) );
  XNOR2_X1 U580 ( .A(n466), .B(n465), .ZN(n470) );
  XNOR2_X1 U581 ( .A(n523), .B(n471), .ZN(n728) );
  XNOR2_X1 U582 ( .A(G902), .B(KEYINPUT15), .ZN(n628) );
  NAND2_X1 U583 ( .A1(n707), .A2(n628), .ZN(n474) );
  OR2_X1 U584 ( .A1(G237), .A2(G902), .ZN(n475) );
  NAND2_X1 U585 ( .A1(n475), .A2(G210), .ZN(n472) );
  XNOR2_X2 U586 ( .A(n474), .B(n473), .ZN(n561) );
  NAND2_X1 U587 ( .A1(G214), .A2(n475), .ZN(n682) );
  NAND2_X1 U588 ( .A1(n561), .A2(n682), .ZN(n536) );
  NOR2_X1 U589 ( .A1(G900), .A2(n749), .ZN(n476) );
  NAND2_X1 U590 ( .A1(n476), .A2(G902), .ZN(n477) );
  NAND2_X1 U591 ( .A1(G952), .A2(n749), .ZN(n578) );
  NAND2_X1 U592 ( .A1(n477), .A2(n578), .ZN(n480) );
  NAND2_X1 U593 ( .A1(G234), .A2(G237), .ZN(n478) );
  XOR2_X1 U594 ( .A(n478), .B(KEYINPUT14), .Z(n698) );
  INV_X1 U595 ( .A(n698), .ZN(n479) );
  NAND2_X1 U596 ( .A1(n480), .A2(n479), .ZN(n549) );
  XNOR2_X1 U597 ( .A(n482), .B(n481), .ZN(n491) );
  INV_X1 U598 ( .A(G953), .ZN(n483) );
  NAND2_X1 U599 ( .A1(n749), .A2(G234), .ZN(n484) );
  XNOR2_X1 U600 ( .A(n485), .B(n484), .ZN(n515) );
  NAND2_X1 U601 ( .A1(G221), .A2(n515), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n486), .B(KEYINPUT93), .ZN(n487) );
  INV_X1 U603 ( .A(n489), .ZN(n490) );
  NAND2_X1 U604 ( .A1(n628), .A2(G234), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n492), .B(KEYINPUT20), .ZN(n497) );
  AND2_X1 U606 ( .A1(G217), .A2(n497), .ZN(n494) );
  INV_X1 U607 ( .A(n664), .ZN(n606) );
  NAND2_X1 U608 ( .A1(G221), .A2(n497), .ZN(n498) );
  XOR2_X1 U609 ( .A(KEYINPUT21), .B(n498), .Z(n663) );
  NAND2_X1 U610 ( .A1(n606), .A2(n663), .ZN(n499) );
  NOR2_X1 U611 ( .A1(n549), .A2(n499), .ZN(n533) );
  XNOR2_X1 U612 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X1 U613 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U614 ( .A(n741), .B(n506), .Z(n512) );
  XOR2_X1 U615 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n508) );
  XNOR2_X1 U616 ( .A(n508), .B(n507), .ZN(n510) );
  NOR2_X1 U617 ( .A1(G953), .A2(G237), .ZN(n524) );
  NAND2_X1 U618 ( .A1(G214), .A2(n524), .ZN(n509) );
  NOR2_X1 U619 ( .A1(G902), .A2(n717), .ZN(n514) );
  XNOR2_X1 U620 ( .A(KEYINPUT13), .B(G475), .ZN(n513) );
  XOR2_X1 U621 ( .A(n560), .B(KEYINPUT99), .Z(n531) );
  NAND2_X1 U622 ( .A1(G217), .A2(n515), .ZN(n516) );
  NOR2_X1 U623 ( .A1(G902), .A2(n720), .ZN(n519) );
  XOR2_X1 U624 ( .A(G478), .B(n519), .Z(n559) );
  INV_X1 U625 ( .A(n559), .ZN(n530) );
  NAND2_X1 U626 ( .A1(n531), .A2(n530), .ZN(n529) );
  NOR2_X1 U627 ( .A1(n632), .A2(G902), .ZN(n525) );
  XOR2_X1 U628 ( .A(n611), .B(KEYINPUT6), .Z(n598) );
  NOR2_X1 U629 ( .A1(n529), .A2(n598), .ZN(n526) );
  NAND2_X1 U630 ( .A1(n533), .A2(n526), .ZN(n570) );
  NOR2_X1 U631 ( .A1(n536), .A2(n570), .ZN(n527) );
  XOR2_X1 U632 ( .A(KEYINPUT36), .B(n527), .Z(n528) );
  NOR2_X1 U633 ( .A1(n577), .A2(n528), .ZN(n655) );
  NOR2_X1 U634 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U635 ( .A(KEYINPUT100), .B(n532), .ZN(n653) );
  NOR2_X1 U636 ( .A1(n650), .A2(n653), .ZN(n615) );
  INV_X1 U637 ( .A(n615), .ZN(n687) );
  OR2_X1 U638 ( .A1(KEYINPUT77), .A2(n687), .ZN(n537) );
  AND2_X1 U639 ( .A1(n667), .A2(n533), .ZN(n534) );
  XNOR2_X1 U640 ( .A(KEYINPUT28), .B(n534), .ZN(n535) );
  NAND2_X1 U641 ( .A1(n535), .A2(n544), .ZN(n564) );
  NOR2_X1 U642 ( .A1(n564), .A2(n585), .ZN(n648) );
  NAND2_X1 U643 ( .A1(n537), .A2(n648), .ZN(n538) );
  NAND2_X1 U644 ( .A1(n538), .A2(KEYINPUT47), .ZN(n540) );
  NAND2_X1 U645 ( .A1(n687), .A2(KEYINPUT77), .ZN(n539) );
  NAND2_X1 U646 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U647 ( .A1(n655), .A2(n541), .ZN(n558) );
  AND2_X1 U648 ( .A1(n648), .A2(n687), .ZN(n542) );
  NOR2_X1 U649 ( .A1(KEYINPUT77), .A2(n542), .ZN(n543) );
  NOR2_X1 U650 ( .A1(KEYINPUT47), .A2(n543), .ZN(n556) );
  XOR2_X1 U651 ( .A(KEYINPUT30), .B(KEYINPUT105), .Z(n548) );
  NAND2_X1 U652 ( .A1(n667), .A2(n682), .ZN(n547) );
  XNOR2_X1 U653 ( .A(n548), .B(n547), .ZN(n550) );
  NOR2_X1 U654 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U655 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U656 ( .A1(n560), .A2(n559), .ZN(n602) );
  NOR2_X1 U657 ( .A1(n566), .A2(n602), .ZN(n554) );
  NAND2_X1 U658 ( .A1(n575), .A2(n554), .ZN(n646) );
  INV_X1 U659 ( .A(n646), .ZN(n555) );
  NOR2_X1 U660 ( .A1(n556), .A2(n555), .ZN(n557) );
  AND2_X1 U661 ( .A1(n558), .A2(n557), .ZN(n569) );
  XOR2_X1 U662 ( .A(KEYINPUT41), .B(KEYINPUT107), .Z(n563) );
  NAND2_X1 U663 ( .A1(n683), .A2(n682), .ZN(n562) );
  INV_X1 U664 ( .A(n683), .ZN(n565) );
  XNOR2_X1 U665 ( .A(n567), .B(KEYINPUT46), .ZN(n568) );
  NOR2_X1 U666 ( .A1(n408), .A2(n570), .ZN(n571) );
  NAND2_X1 U667 ( .A1(n682), .A2(n571), .ZN(n572) );
  XNOR2_X1 U668 ( .A(n572), .B(KEYINPUT103), .ZN(n573) );
  XNOR2_X1 U669 ( .A(n573), .B(KEYINPUT43), .ZN(n574) );
  NOR2_X1 U670 ( .A1(n575), .A2(n574), .ZN(n658) );
  NAND2_X1 U671 ( .A1(n576), .A2(n653), .ZN(n657) );
  NOR2_X1 U672 ( .A1(n578), .A2(n698), .ZN(n583) );
  NOR2_X1 U673 ( .A1(G898), .A2(n749), .ZN(n579) );
  XNOR2_X1 U674 ( .A(KEYINPUT90), .B(n579), .ZN(n730) );
  NAND2_X1 U675 ( .A1(G902), .A2(n730), .ZN(n580) );
  NOR2_X1 U676 ( .A1(n698), .A2(n580), .ZN(n581) );
  XOR2_X1 U677 ( .A(KEYINPUT91), .B(n581), .Z(n582) );
  NOR2_X1 U678 ( .A1(n583), .A2(n582), .ZN(n584) );
  INV_X1 U679 ( .A(KEYINPUT0), .ZN(n586) );
  NAND2_X1 U680 ( .A1(n681), .A2(n663), .ZN(n588) );
  INV_X1 U681 ( .A(KEYINPUT32), .ZN(n589) );
  NAND2_X1 U682 ( .A1(n606), .A2(n592), .ZN(n593) );
  INV_X1 U683 ( .A(KEYINPUT83), .ZN(n594) );
  XNOR2_X1 U684 ( .A(n619), .B(n594), .ZN(n596) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U686 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U687 ( .A1(n597), .A2(KEYINPUT82), .ZN(n604) );
  AND2_X1 U688 ( .A1(n664), .A2(n663), .ZN(n670) );
  XNOR2_X1 U689 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n599) );
  INV_X1 U690 ( .A(n754), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n624) );
  NOR2_X1 U692 ( .A1(n611), .A2(n607), .ZN(n676) );
  NAND2_X1 U693 ( .A1(n676), .A2(n608), .ZN(n609) );
  XNOR2_X1 U694 ( .A(KEYINPUT31), .B(n609), .ZN(n652) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U696 ( .A(KEYINPUT95), .B(n613), .ZN(n638) );
  NOR2_X1 U697 ( .A1(n652), .A2(n638), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n617) );
  NOR2_X1 U699 ( .A1(KEYINPUT44), .A2(KEYINPUT82), .ZN(n616) );
  INV_X1 U700 ( .A(KEYINPUT45), .ZN(n625) );
  NOR2_X1 U701 ( .A1(n747), .A2(n734), .ZN(n627) );
  NOR2_X2 U702 ( .A1(n627), .A2(KEYINPUT78), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n660), .B(KEYINPUT2), .ZN(n630) );
  AND2_X2 U705 ( .A1(n631), .A2(n630), .ZN(n722) );
  XOR2_X1 U706 ( .A(n632), .B(KEYINPUT62), .Z(n633) );
  INV_X1 U707 ( .A(n635), .ZN(n636) );
  XOR2_X1 U708 ( .A(G101), .B(n636), .Z(G3) );
  NAND2_X1 U709 ( .A1(n638), .A2(n650), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(G104), .ZN(G6) );
  XOR2_X1 U711 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  NAND2_X1 U712 ( .A1(n638), .A2(n653), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n642) );
  XOR2_X1 U714 ( .A(G107), .B(KEYINPUT109), .Z(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(G9) );
  XOR2_X1 U716 ( .A(n643), .B(G110), .Z(G12) );
  XOR2_X1 U717 ( .A(G128), .B(KEYINPUT29), .Z(n645) );
  NAND2_X1 U718 ( .A1(n648), .A2(n653), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(G30) );
  XNOR2_X1 U720 ( .A(G143), .B(KEYINPUT110), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(G45) );
  NAND2_X1 U722 ( .A1(n648), .A2(n650), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(G146), .ZN(G48) );
  NAND2_X1 U724 ( .A1(n652), .A2(n650), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(G113), .ZN(G15) );
  NAND2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n654), .B(G116), .ZN(G18) );
  XNOR2_X1 U728 ( .A(G125), .B(n655), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U730 ( .A(G134), .B(n657), .ZN(G36) );
  XNOR2_X1 U731 ( .A(G140), .B(n658), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT111), .ZN(G42) );
  NAND2_X1 U733 ( .A1(KEYINPUT76), .A2(n660), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT2), .ZN(n704) );
  NOR2_X1 U735 ( .A1(n680), .A2(n692), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(KEYINPUT117), .ZN(n701) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U738 ( .A(KEYINPUT49), .B(n665), .Z(n666) );
  NOR2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U740 ( .A(KEYINPUT112), .B(n668), .Z(n673) );
  NOR2_X1 U741 ( .A1(n670), .A2(n408), .ZN(n671) );
  XNOR2_X1 U742 ( .A(KEYINPUT50), .B(n671), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U744 ( .A(KEYINPUT113), .B(n674), .Z(n675) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U746 ( .A(n677), .B(KEYINPUT114), .Z(n678) );
  XNOR2_X1 U747 ( .A(KEYINPUT51), .B(n678), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n695) );
  INV_X1 U749 ( .A(n681), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U751 ( .A(KEYINPUT115), .B(n684), .Z(n685) );
  NOR2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U754 ( .A(KEYINPUT116), .B(n689), .Z(n690) );
  NOR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n693) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U758 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n699), .A2(G952), .ZN(n700) );
  NAND2_X1 U761 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U762 ( .A(KEYINPUT118), .B(n702), .Z(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U764 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U765 ( .A(n706), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U766 ( .A1(n722), .A2(G210), .ZN(n710) );
  INV_X1 U767 ( .A(n707), .ZN(n709) );
  XOR2_X1 U768 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n708) );
  NAND2_X1 U769 ( .A1(n722), .A2(G469), .ZN(n715) );
  XOR2_X1 U770 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n712) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n711) );
  XNOR2_X1 U772 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n726), .A2(n716), .ZN(G54) );
  NAND2_X1 U774 ( .A1(n722), .A2(G475), .ZN(n718) );
  NAND2_X1 U775 ( .A1(G478), .A2(n722), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n726), .A2(n721), .ZN(G63) );
  NAND2_X1 U778 ( .A1(n722), .A2(G217), .ZN(n723) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(G66) );
  XOR2_X1 U780 ( .A(n728), .B(n727), .Z(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n738) );
  XOR2_X1 U782 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n732) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n733), .A2(G898), .ZN(n736) );
  OR2_X1 U786 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(KEYINPUT124), .B(n739), .ZN(G69) );
  XNOR2_X1 U790 ( .A(n740), .B(n741), .ZN(n742) );
  XOR2_X1 U791 ( .A(n742), .B(KEYINPUT125), .Z(n748) );
  INV_X1 U792 ( .A(n748), .ZN(n743) );
  XOR2_X1 U793 ( .A(KEYINPUT127), .B(n743), .Z(n744) );
  XNOR2_X1 U794 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G953), .ZN(n753) );
  XOR2_X1 U797 ( .A(n748), .B(n747), .Z(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U799 ( .A(KEYINPUT126), .B(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U801 ( .A(n754), .B(G122), .Z(G24) );
  XOR2_X1 U802 ( .A(G119), .B(n755), .Z(G21) );
  XOR2_X1 U803 ( .A(n756), .B(G131), .Z(G33) );
  XOR2_X1 U804 ( .A(G137), .B(n757), .Z(G39) );
endmodule

