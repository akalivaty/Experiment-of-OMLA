

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770;

  BUF_X1 U373 ( .A(n716), .Z(n358) );
  AND2_X1 U374 ( .A1(n429), .A2(n646), .ZN(n428) );
  INV_X1 U375 ( .A(n628), .ZN(n354) );
  INV_X1 U376 ( .A(n352), .ZN(n351) );
  AND2_X1 U377 ( .A1(n437), .A2(n436), .ZN(n435) );
  INV_X1 U378 ( .A(KEYINPUT44), .ZN(n353) );
  XNOR2_X1 U379 ( .A(n356), .B(n355), .ZN(n767) );
  NAND2_X1 U380 ( .A1(n412), .A2(n411), .ZN(n356) );
  INV_X1 U381 ( .A(n624), .ZN(n355) );
  XNOR2_X1 U382 ( .A(n478), .B(n610), .ZN(n616) );
  XNOR2_X1 U383 ( .A(n541), .B(n386), .ZN(n357) );
  XNOR2_X1 U384 ( .A(n479), .B(n532), .ZN(n423) );
  XNOR2_X1 U385 ( .A(n550), .B(KEYINPUT4), .ZN(n522) );
  XNOR2_X1 U386 ( .A(KEYINPUT93), .B(G104), .ZN(n487) );
  XNOR2_X1 U387 ( .A(n423), .B(n460), .ZN(n654) );
  NAND2_X1 U388 ( .A1(n354), .A2(n351), .ZN(n627) );
  NAND2_X1 U389 ( .A1(n768), .A2(n353), .ZN(n352) );
  NAND2_X1 U390 ( .A1(n619), .A2(n696), .ZN(n635) );
  XNOR2_X1 U391 ( .A(n575), .B(KEYINPUT1), .ZN(n619) );
  XNOR2_X2 U392 ( .A(n522), .B(n357), .ZN(n753) );
  INV_X2 U393 ( .A(KEYINPUT69), .ZN(n388) );
  XOR2_X1 U394 ( .A(n362), .B(KEYINPUT19), .Z(n359) );
  XNOR2_X2 U395 ( .A(n593), .B(n447), .ZN(n446) );
  NOR2_X2 U396 ( .A1(n670), .A2(n559), .ZN(n560) );
  INV_X2 U397 ( .A(G953), .ZN(n757) );
  XNOR2_X1 U398 ( .A(n627), .B(KEYINPUT76), .ZN(n427) );
  XNOR2_X1 U399 ( .A(n582), .B(n419), .ZN(n769) );
  NAND2_X1 U400 ( .A1(n441), .A2(n439), .ZN(n394) );
  AND2_X1 U401 ( .A1(n431), .A2(n442), .ZN(n441) );
  NAND2_X1 U402 ( .A1(n471), .A2(n466), .ZN(n580) );
  XNOR2_X1 U403 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U404 ( .A(n546), .B(n547), .ZN(n584) );
  NOR2_X1 U405 ( .A1(G902), .A2(n732), .ZN(n546) );
  BUF_X1 U406 ( .A(n674), .Z(n360) );
  XNOR2_X1 U407 ( .A(n581), .B(KEYINPUT108), .ZN(n674) );
  XNOR2_X1 U408 ( .A(KEYINPUT30), .B(n361), .ZN(n578) );
  AND2_X1 U409 ( .A1(n706), .A2(n614), .ZN(n361) );
  NAND2_X1 U410 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U411 ( .A1(n416), .A2(n706), .ZN(n362) );
  NAND2_X1 U412 ( .A1(n425), .A2(n706), .ZN(n574) );
  XNOR2_X1 U413 ( .A(n544), .B(n545), .ZN(n732) );
  XNOR2_X1 U414 ( .A(n574), .B(KEYINPUT19), .ZN(n607) );
  XNOR2_X1 U415 ( .A(n387), .B(G134), .ZN(n386) );
  INV_X1 U416 ( .A(KEYINPUT70), .ZN(n387) );
  XNOR2_X1 U417 ( .A(G140), .B(G137), .ZN(n496) );
  OR2_X1 U418 ( .A1(n740), .A2(G902), .ZN(n464) );
  XOR2_X1 U419 ( .A(G116), .B(G107), .Z(n552) );
  XNOR2_X1 U420 ( .A(n481), .B(G110), .ZN(n530) );
  INV_X1 U421 ( .A(G119), .ZN(n481) );
  XNOR2_X1 U422 ( .A(n543), .B(n496), .ZN(n755) );
  NOR2_X1 U423 ( .A1(G902), .A2(n737), .ZN(n556) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n534) );
  XOR2_X1 U425 ( .A(KEYINPUT5), .B(G137), .Z(n514) );
  XNOR2_X1 U426 ( .A(G116), .B(G119), .ZN(n513) );
  INV_X1 U427 ( .A(G146), .ZN(n420) );
  XNOR2_X1 U428 ( .A(n453), .B(n413), .ZN(n412) );
  INV_X1 U429 ( .A(KEYINPUT34), .ZN(n413) );
  NAND2_X1 U430 ( .A1(n613), .A2(n375), .ZN(n442) );
  NAND2_X1 U431 ( .A1(n363), .A2(KEYINPUT109), .ZN(n469) );
  NAND2_X1 U432 ( .A1(n476), .A2(n475), .ZN(n474) );
  NAND2_X1 U433 ( .A1(n567), .A2(n566), .ZN(n472) );
  AND2_X1 U434 ( .A1(n618), .A2(n408), .ZN(n696) );
  XNOR2_X1 U435 ( .A(n542), .B(n531), .ZN(n482) );
  XNOR2_X1 U436 ( .A(KEYINPUT16), .B(KEYINPUT93), .ZN(n531) );
  XNOR2_X1 U437 ( .A(n543), .B(n368), .ZN(n544) );
  XNOR2_X1 U438 ( .A(n686), .B(n407), .ZN(n650) );
  INV_X1 U439 ( .A(KEYINPUT2), .ZN(n407) );
  XNOR2_X1 U440 ( .A(n409), .B(KEYINPUT39), .ZN(n597) );
  NAND2_X1 U441 ( .A1(n580), .A2(n579), .ZN(n409) );
  XNOR2_X1 U442 ( .A(KEYINPUT22), .B(KEYINPUT67), .ZN(n610) );
  XNOR2_X1 U443 ( .A(n465), .B(n755), .ZN(n740) );
  XNOR2_X1 U444 ( .A(n452), .B(n450), .ZN(n737) );
  XNOR2_X1 U445 ( .A(n451), .B(n367), .ZN(n450) );
  NOR2_X1 U446 ( .A1(n689), .A2(n372), .ZN(n397) );
  INV_X1 U447 ( .A(KEYINPUT91), .ZN(n443) );
  XNOR2_X1 U448 ( .A(n571), .B(KEYINPUT84), .ZN(n391) );
  INV_X1 U449 ( .A(KEYINPUT72), .ZN(n444) );
  XNOR2_X1 U450 ( .A(KEYINPUT48), .B(KEYINPUT71), .ZN(n592) );
  INV_X1 U451 ( .A(KEYINPUT8), .ZN(n462) );
  NAND2_X1 U452 ( .A1(n757), .A2(G234), .ZN(n463) );
  XOR2_X1 U453 ( .A(G140), .B(KEYINPUT12), .Z(n538) );
  XNOR2_X1 U454 ( .A(G113), .B(G143), .ZN(n537) );
  XNOR2_X1 U455 ( .A(n495), .B(KEYINPUT10), .ZN(n543) );
  XOR2_X1 U456 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n535) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT15), .ZN(n648) );
  INV_X1 U458 ( .A(n683), .ZN(n686) );
  XNOR2_X1 U459 ( .A(n524), .B(n523), .ZN(n526) );
  INV_X1 U460 ( .A(KEYINPUT81), .ZN(n523) );
  XOR2_X1 U461 ( .A(G125), .B(G146), .Z(n521) );
  XNOR2_X1 U462 ( .A(n406), .B(n376), .ZN(n716) );
  NOR2_X1 U463 ( .A1(n635), .A2(n620), .ZN(n406) );
  NAND2_X1 U464 ( .A1(G234), .A2(G237), .ZN(n505) );
  OR2_X1 U465 ( .A1(G237), .A2(G902), .ZN(n533) );
  INV_X1 U466 ( .A(KEYINPUT38), .ZN(n424) );
  INV_X1 U467 ( .A(n622), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n515), .B(n366), .ZN(n516) );
  XOR2_X1 U469 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n501) );
  XNOR2_X1 U470 ( .A(n549), .B(n548), .ZN(n451) );
  XNOR2_X1 U471 ( .A(G122), .B(KEYINPUT7), .ZN(n548) );
  XOR2_X1 U472 ( .A(G134), .B(KEYINPUT104), .Z(n549) );
  XNOR2_X1 U473 ( .A(n373), .B(n485), .ZN(n454) );
  NAND2_X1 U474 ( .A1(n440), .A2(n365), .ZN(n439) );
  NAND2_X1 U475 ( .A1(n470), .A2(n467), .ZN(n466) );
  AND2_X1 U476 ( .A1(n473), .A2(n472), .ZN(n471) );
  NAND2_X1 U477 ( .A1(n469), .A2(n468), .ZN(n467) );
  INV_X1 U478 ( .A(KEYINPUT100), .ZN(n563) );
  INV_X1 U479 ( .A(KEYINPUT0), .ZN(n430) );
  XNOR2_X1 U480 ( .A(n482), .B(n480), .ZN(n479) );
  INV_X1 U481 ( .A(n530), .ZN(n480) );
  INV_X1 U482 ( .A(KEYINPUT40), .ZN(n419) );
  AND2_X1 U483 ( .A1(n597), .A2(n581), .ZN(n582) );
  INV_X1 U484 ( .A(KEYINPUT82), .ZN(n456) );
  XNOR2_X1 U485 ( .A(n739), .B(n740), .ZN(n395) );
  XNOR2_X1 U486 ( .A(n736), .B(n737), .ZN(n398) );
  INV_X1 U487 ( .A(KEYINPUT60), .ZN(n421) );
  INV_X1 U488 ( .A(KEYINPUT56), .ZN(n401) );
  NOR2_X1 U489 ( .A1(n723), .A2(G953), .ZN(n724) );
  AND2_X1 U490 ( .A1(n565), .A2(KEYINPUT78), .ZN(n363) );
  XOR2_X1 U491 ( .A(n504), .B(KEYINPUT25), .Z(n364) );
  NOR2_X1 U492 ( .A1(n613), .A2(n375), .ZN(n365) );
  INV_X1 U493 ( .A(n690), .ZN(n408) );
  XOR2_X1 U494 ( .A(n514), .B(n513), .Z(n366) );
  XNOR2_X1 U495 ( .A(KEYINPUT103), .B(KEYINPUT9), .ZN(n367) );
  XOR2_X1 U496 ( .A(n542), .B(n541), .Z(n368) );
  AND2_X1 U497 ( .A1(G210), .A2(n533), .ZN(n369) );
  OR2_X1 U498 ( .A1(KEYINPUT2), .A2(n684), .ZN(n370) );
  NOR2_X1 U499 ( .A1(n596), .A2(n416), .ZN(n371) );
  AND2_X1 U500 ( .A1(n722), .A2(n721), .ZN(n372) );
  AND2_X1 U501 ( .A1(G227), .A2(n757), .ZN(n373) );
  AND2_X1 U502 ( .A1(n609), .A2(n408), .ZN(n374) );
  XNOR2_X1 U503 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n375) );
  XNOR2_X1 U504 ( .A(KEYINPUT75), .B(n621), .ZN(n376) );
  XOR2_X1 U505 ( .A(KEYINPUT36), .B(KEYINPUT112), .Z(n377) );
  XOR2_X1 U506 ( .A(n651), .B(KEYINPUT62), .Z(n378) );
  XNOR2_X1 U507 ( .A(n732), .B(KEYINPUT59), .ZN(n379) );
  XOR2_X1 U508 ( .A(n656), .B(n655), .Z(n380) );
  AND2_X1 U509 ( .A1(n399), .A2(KEYINPUT2), .ZN(n381) );
  NOR2_X1 U510 ( .A1(G952), .A2(n757), .ZN(n741) );
  XOR2_X1 U511 ( .A(n653), .B(KEYINPUT114), .Z(n382) );
  INV_X1 U512 ( .A(KEYINPUT83), .ZN(n399) );
  XNOR2_X1 U513 ( .A(n405), .B(n486), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n487), .B(KEYINPUT96), .ZN(n405) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n488) );
  XNOR2_X1 U516 ( .A(n414), .B(n377), .ZN(n576) );
  NAND2_X1 U517 ( .A1(n435), .A2(n432), .ZN(n383) );
  NAND2_X1 U518 ( .A1(n435), .A2(n432), .ZN(n628) );
  XNOR2_X1 U519 ( .A(n555), .B(n553), .ZN(n452) );
  XOR2_X1 U520 ( .A(G478), .B(n556), .Z(n583) );
  BUF_X1 U521 ( .A(n654), .Z(n384) );
  BUF_X1 U522 ( .A(n425), .Z(n416) );
  NAND2_X1 U523 ( .A1(n394), .A2(n443), .ZN(n437) );
  NAND2_X1 U524 ( .A1(n385), .A2(n374), .ZN(n478) );
  XNOR2_X2 U525 ( .A(n608), .B(n430), .ZN(n385) );
  NAND2_X1 U526 ( .A1(n702), .A2(n385), .ZN(n636) );
  NAND2_X1 U527 ( .A1(n385), .A2(n638), .ZN(n639) );
  NAND2_X1 U528 ( .A1(n716), .A2(n385), .ZN(n453) );
  XNOR2_X2 U529 ( .A(n388), .B(G131), .ZN(n541) );
  XNOR2_X1 U530 ( .A(n389), .B(n444), .ZN(n591) );
  NAND2_X1 U531 ( .A1(n393), .A2(n390), .ZN(n389) );
  NOR2_X1 U532 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U533 ( .A1(n562), .A2(n561), .ZN(n392) );
  XNOR2_X1 U534 ( .A(n764), .B(KEYINPUT89), .ZN(n393) );
  XNOR2_X2 U535 ( .A(n577), .B(KEYINPUT113), .ZN(n764) );
  INV_X1 U536 ( .A(n394), .ZN(n433) );
  XNOR2_X1 U537 ( .A(n433), .B(G119), .ZN(G21) );
  XNOR2_X1 U538 ( .A(n649), .B(n648), .ZN(n396) );
  NOR2_X1 U539 ( .A1(n395), .A2(n741), .ZN(G66) );
  AND2_X2 U540 ( .A1(n396), .A2(n650), .ZN(n731) );
  NAND2_X1 U541 ( .A1(n370), .A2(n397), .ZN(n410) );
  NAND2_X1 U542 ( .A1(n683), .A2(n381), .ZN(n687) );
  XNOR2_X1 U543 ( .A(n519), .B(n520), .ZN(n458) );
  XNOR2_X1 U544 ( .A(n629), .B(KEYINPUT64), .ZN(n429) );
  NOR2_X1 U545 ( .A1(n664), .A2(n443), .ZN(n434) );
  NOR2_X1 U546 ( .A1(n398), .A2(n741), .ZN(G63) );
  INV_X1 U547 ( .A(n584), .ZN(n557) );
  XNOR2_X1 U548 ( .A(n400), .B(n382), .ZN(G57) );
  NAND2_X1 U549 ( .A1(n403), .A2(n734), .ZN(n400) );
  XNOR2_X1 U550 ( .A(n402), .B(n401), .ZN(G51) );
  NAND2_X1 U551 ( .A1(n404), .A2(n734), .ZN(n402) );
  NAND2_X1 U552 ( .A1(n383), .A2(KEYINPUT44), .ZN(n629) );
  XNOR2_X1 U553 ( .A(n652), .B(n378), .ZN(n403) );
  XNOR2_X1 U554 ( .A(n657), .B(n380), .ZN(n404) );
  NAND2_X1 U555 ( .A1(n554), .A2(G217), .ZN(n555) );
  XNOR2_X2 U556 ( .A(n463), .B(n462), .ZN(n554) );
  NOR2_X2 U557 ( .A1(n557), .A2(n583), .ZN(n581) );
  NAND2_X1 U558 ( .A1(n664), .A2(n443), .ZN(n436) );
  XNOR2_X2 U559 ( .A(n464), .B(n364), .ZN(n618) );
  NAND2_X1 U560 ( .A1(n769), .A2(n770), .ZN(n589) );
  NAND2_X1 U561 ( .A1(n731), .A2(G472), .ZN(n652) );
  XNOR2_X1 U562 ( .A(n410), .B(KEYINPUT124), .ZN(n723) );
  XNOR2_X1 U563 ( .A(n683), .B(n399), .ZN(n684) );
  NAND2_X1 U564 ( .A1(n654), .A2(n648), .ZN(n459) );
  INV_X4 U565 ( .A(G122), .ZN(n483) );
  AND2_X2 U566 ( .A1(n438), .A2(n691), .ZN(n664) );
  NAND2_X1 U567 ( .A1(n446), .A2(n445), .ZN(n414) );
  NAND2_X1 U568 ( .A1(n434), .A2(n433), .ZN(n432) );
  XNOR2_X1 U569 ( .A(n502), .B(n417), .ZN(n465) );
  XNOR2_X1 U570 ( .A(n500), .B(n501), .ZN(n417) );
  XNOR2_X1 U571 ( .A(n418), .B(n592), .ZN(n600) );
  NAND2_X1 U572 ( .A1(n590), .A2(n591), .ZN(n418) );
  XNOR2_X2 U573 ( .A(n753), .B(n420), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n614), .A2(n573), .ZN(n519) );
  XNOR2_X2 U575 ( .A(n640), .B(KEYINPUT106), .ZN(n614) );
  XNOR2_X1 U576 ( .A(n422), .B(n421), .ZN(G60) );
  NAND2_X1 U577 ( .A1(n735), .A2(n734), .ZN(n422) );
  AND2_X2 U578 ( .A1(n683), .A2(n647), .ZN(n649) );
  NAND2_X2 U579 ( .A1(n748), .A2(n756), .ZN(n683) );
  XNOR2_X1 U580 ( .A(n423), .B(KEYINPUT127), .ZN(n742) );
  XNOR2_X1 U581 ( .A(n416), .B(n424), .ZN(n707) );
  NAND2_X1 U582 ( .A1(n569), .A2(n416), .ZN(n669) );
  XNOR2_X2 U583 ( .A(n459), .B(n369), .ZN(n425) );
  XNOR2_X2 U584 ( .A(n426), .B(KEYINPUT45), .ZN(n748) );
  XNOR2_X1 U585 ( .A(n461), .B(n617), .ZN(n438) );
  NAND2_X1 U586 ( .A1(n632), .A2(n375), .ZN(n431) );
  INV_X1 U587 ( .A(n632), .ZN(n440) );
  INV_X1 U588 ( .A(n362), .ZN(n445) );
  INV_X1 U589 ( .A(KEYINPUT111), .ZN(n447) );
  AND2_X2 U590 ( .A1(n448), .A2(n674), .ZN(n593) );
  AND2_X1 U591 ( .A1(n449), .A2(n573), .ZN(n448) );
  INV_X1 U592 ( .A(n620), .ZN(n449) );
  XNOR2_X2 U593 ( .A(n457), .B(n456), .ZN(n670) );
  NOR2_X2 U594 ( .A1(n586), .A2(n359), .ZN(n457) );
  NAND2_X1 U595 ( .A1(n458), .A2(n575), .ZN(n586) );
  XNOR2_X1 U596 ( .A(n527), .B(n528), .ZN(n460) );
  NAND2_X1 U597 ( .A1(n616), .A2(n615), .ZN(n461) );
  XNOR2_X1 U598 ( .A(n488), .B(n496), .ZN(n489) );
  NAND2_X1 U599 ( .A1(n477), .A2(n566), .ZN(n468) );
  INV_X1 U600 ( .A(n638), .ZN(n470) );
  NAND2_X1 U601 ( .A1(n638), .A2(n474), .ZN(n473) );
  NAND2_X1 U602 ( .A1(KEYINPUT109), .A2(n566), .ZN(n475) );
  NAND2_X1 U603 ( .A1(n363), .A2(n477), .ZN(n476) );
  INV_X1 U604 ( .A(KEYINPUT109), .ZN(n477) );
  XNOR2_X2 U605 ( .A(n483), .B(G104), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X2 U607 ( .A1(n651), .A2(G902), .ZN(n518) );
  XNOR2_X2 U608 ( .A(n491), .B(n490), .ZN(n575) );
  NOR2_X2 U609 ( .A1(G902), .A2(n725), .ZN(n491) );
  XOR2_X1 U610 ( .A(n498), .B(n497), .Z(n484) );
  XNOR2_X1 U611 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U612 ( .A(n499), .B(n484), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n517), .B(n489), .ZN(n725) );
  INV_X1 U614 ( .A(KEYINPUT35), .ZN(n623) );
  XNOR2_X1 U615 ( .A(n623), .B(KEYINPUT87), .ZN(n624) );
  INV_X1 U616 ( .A(n741), .ZN(n734) );
  XOR2_X1 U617 ( .A(KEYINPUT80), .B(G110), .Z(n486) );
  XNOR2_X1 U618 ( .A(G101), .B(G107), .ZN(n485) );
  XNOR2_X2 U619 ( .A(G143), .B(G128), .ZN(n550) );
  XNOR2_X1 U620 ( .A(KEYINPUT73), .B(G469), .ZN(n490) );
  XOR2_X1 U621 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n520) );
  XOR2_X1 U622 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n493) );
  NAND2_X1 U623 ( .A1(G234), .A2(n648), .ZN(n492) );
  XNOR2_X1 U624 ( .A(n493), .B(n492), .ZN(n503) );
  NAND2_X1 U625 ( .A1(n503), .A2(G221), .ZN(n494) );
  XNOR2_X1 U626 ( .A(n494), .B(KEYINPUT21), .ZN(n690) );
  INV_X1 U627 ( .A(n521), .ZN(n495) );
  NAND2_X1 U628 ( .A1(G221), .A2(n554), .ZN(n499) );
  XOR2_X1 U629 ( .A(KEYINPUT23), .B(KEYINPUT79), .Z(n498) );
  XNOR2_X1 U630 ( .A(G128), .B(KEYINPUT24), .ZN(n497) );
  XNOR2_X1 U631 ( .A(n530), .B(KEYINPUT74), .ZN(n500) );
  NAND2_X1 U632 ( .A1(n503), .A2(G217), .ZN(n504) );
  NOR2_X1 U633 ( .A1(n690), .A2(n618), .ZN(n510) );
  XNOR2_X1 U634 ( .A(n505), .B(KEYINPUT14), .ZN(n507) );
  NAND2_X1 U635 ( .A1(G902), .A2(n507), .ZN(n601) );
  NOR2_X1 U636 ( .A1(G900), .A2(n601), .ZN(n506) );
  NAND2_X1 U637 ( .A1(G953), .A2(n506), .ZN(n509) );
  NAND2_X1 U638 ( .A1(n507), .A2(G952), .ZN(n508) );
  XOR2_X1 U639 ( .A(KEYINPUT94), .B(n508), .Z(n721) );
  NAND2_X1 U640 ( .A1(n757), .A2(n721), .ZN(n604) );
  NAND2_X1 U641 ( .A1(n509), .A2(n604), .ZN(n565) );
  AND2_X1 U642 ( .A1(n510), .A2(n565), .ZN(n573) );
  XNOR2_X1 U643 ( .A(G101), .B(KEYINPUT3), .ZN(n511) );
  XNOR2_X1 U644 ( .A(n511), .B(G113), .ZN(n529) );
  NAND2_X1 U645 ( .A1(n534), .A2(G210), .ZN(n512) );
  XNOR2_X1 U646 ( .A(n529), .B(n512), .ZN(n515) );
  XNOR2_X2 U647 ( .A(n517), .B(n516), .ZN(n651) );
  XNOR2_X2 U648 ( .A(n518), .B(G472), .ZN(n694) );
  INV_X1 U649 ( .A(n694), .ZN(n640) );
  XNOR2_X1 U650 ( .A(n522), .B(n521), .ZN(n528) );
  XOR2_X1 U651 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n524) );
  NAND2_X1 U652 ( .A1(G224), .A2(n757), .ZN(n525) );
  XNOR2_X1 U653 ( .A(n529), .B(n552), .ZN(n532) );
  NAND2_X1 U654 ( .A1(G214), .A2(n533), .ZN(n706) );
  XOR2_X1 U655 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n558) );
  XNOR2_X1 U656 ( .A(KEYINPUT13), .B(G475), .ZN(n547) );
  NAND2_X1 U657 ( .A1(n534), .A2(G214), .ZN(n536) );
  XNOR2_X1 U658 ( .A(n536), .B(n535), .ZN(n540) );
  XNOR2_X1 U659 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U660 ( .A(n540), .B(n539), .Z(n545) );
  INV_X1 U661 ( .A(n550), .ZN(n551) );
  XNOR2_X1 U662 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U663 ( .A1(n557), .A2(n583), .ZN(n665) );
  INV_X1 U664 ( .A(n665), .ZN(n677) );
  NOR2_X1 U665 ( .A1(n581), .A2(n677), .ZN(n711) );
  XNOR2_X1 U666 ( .A(KEYINPUT85), .B(n711), .ZN(n634) );
  NAND2_X1 U667 ( .A1(n558), .A2(n634), .ZN(n559) );
  XNOR2_X1 U668 ( .A(n560), .B(KEYINPUT77), .ZN(n562) );
  NAND2_X1 U669 ( .A1(n670), .A2(KEYINPUT47), .ZN(n561) );
  INV_X1 U670 ( .A(n618), .ZN(n691) );
  NAND2_X1 U671 ( .A1(n696), .A2(n575), .ZN(n564) );
  XNOR2_X2 U672 ( .A(n564), .B(n563), .ZN(n638) );
  INV_X1 U673 ( .A(n565), .ZN(n567) );
  INV_X1 U674 ( .A(KEYINPUT78), .ZN(n566) );
  NAND2_X1 U675 ( .A1(n580), .A2(n578), .ZN(n568) );
  NAND2_X1 U676 ( .A1(n584), .A2(n583), .ZN(n622) );
  NOR2_X1 U677 ( .A1(n568), .A2(n622), .ZN(n569) );
  NAND2_X1 U678 ( .A1(KEYINPUT47), .A2(n711), .ZN(n570) );
  NAND2_X1 U679 ( .A1(n669), .A2(n570), .ZN(n571) );
  INV_X1 U680 ( .A(KEYINPUT6), .ZN(n572) );
  XNOR2_X1 U681 ( .A(n572), .B(n694), .ZN(n620) );
  INV_X1 U682 ( .A(n619), .ZN(n611) );
  INV_X1 U683 ( .A(n611), .ZN(n695) );
  NAND2_X1 U684 ( .A1(n576), .A2(n695), .ZN(n577) );
  AND2_X1 U685 ( .A1(n578), .A2(n707), .ZN(n579) );
  NOR2_X1 U686 ( .A1(n584), .A2(n583), .ZN(n609) );
  INV_X1 U687 ( .A(n609), .ZN(n709) );
  NAND2_X1 U688 ( .A1(n707), .A2(n706), .ZN(n712) );
  NOR2_X1 U689 ( .A1(n709), .A2(n712), .ZN(n585) );
  XNOR2_X1 U690 ( .A(n585), .B(KEYINPUT41), .ZN(n685) );
  NOR2_X1 U691 ( .A1(n685), .A2(n586), .ZN(n587) );
  XOR2_X1 U692 ( .A(KEYINPUT42), .B(n587), .Z(n770) );
  XOR2_X1 U693 ( .A(KEYINPUT46), .B(KEYINPUT88), .Z(n588) );
  XNOR2_X1 U694 ( .A(n589), .B(n588), .ZN(n590) );
  NAND2_X1 U695 ( .A1(n593), .A2(n706), .ZN(n594) );
  NOR2_X1 U696 ( .A1(n695), .A2(n594), .ZN(n595) );
  XNOR2_X1 U697 ( .A(n595), .B(KEYINPUT43), .ZN(n596) );
  NAND2_X1 U698 ( .A1(n597), .A2(n677), .ZN(n681) );
  INV_X1 U699 ( .A(n681), .ZN(n598) );
  NOR2_X1 U700 ( .A1(n371), .A2(n598), .ZN(n599) );
  AND2_X2 U701 ( .A1(n600), .A2(n599), .ZN(n756) );
  INV_X1 U702 ( .A(n601), .ZN(n602) );
  NOR2_X1 U703 ( .A1(G898), .A2(n757), .ZN(n743) );
  NAND2_X1 U704 ( .A1(n602), .A2(n743), .ZN(n603) );
  NAND2_X1 U705 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U706 ( .A(KEYINPUT95), .B(n605), .Z(n606) );
  NAND2_X1 U707 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U708 ( .A1(n620), .A2(n616), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n611), .A2(n618), .ZN(n612) );
  XNOR2_X1 U710 ( .A(n612), .B(KEYINPUT105), .ZN(n613) );
  INV_X1 U711 ( .A(KEYINPUT66), .ZN(n617) );
  NOR2_X1 U712 ( .A1(n695), .A2(n614), .ZN(n615) );
  XOR2_X1 U713 ( .A(KEYINPUT107), .B(KEYINPUT33), .Z(n621) );
  INV_X1 U714 ( .A(n767), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n630), .A2(KEYINPUT44), .ZN(n631) );
  XNOR2_X1 U716 ( .A(n631), .B(KEYINPUT90), .ZN(n645) );
  OR2_X1 U717 ( .A1(n632), .A2(n695), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n691), .A2(n633), .ZN(n658) );
  INV_X1 U719 ( .A(n634), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT31), .B(KEYINPUT101), .Z(n637) );
  NOR2_X1 U721 ( .A1(n694), .A2(n635), .ZN(n702) );
  XNOR2_X1 U722 ( .A(n637), .B(n636), .ZN(n678) );
  NOR2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n660) );
  NOR2_X1 U724 ( .A1(n678), .A2(n660), .ZN(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U726 ( .A1(n658), .A2(n643), .ZN(n644) );
  AND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  INV_X1 U728 ( .A(KEYINPUT86), .ZN(n647) );
  INV_X1 U729 ( .A(KEYINPUT63), .ZN(n653) );
  XNOR2_X1 U730 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n384), .B(KEYINPUT92), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n731), .A2(G210), .ZN(n657) );
  XOR2_X1 U733 ( .A(G101), .B(n658), .Z(G3) );
  NAND2_X1 U734 ( .A1(n360), .A2(n660), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(G104), .ZN(G6) );
  XOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n662) );
  NAND2_X1 U737 ( .A1(n660), .A2(n677), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(G107), .B(n663), .ZN(G9) );
  XOR2_X1 U740 ( .A(n664), .B(G110), .Z(G12) );
  NOR2_X1 U741 ( .A1(n670), .A2(n665), .ZN(n667) );
  XNOR2_X1 U742 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n666) );
  XNOR2_X1 U743 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U744 ( .A(G128), .B(n668), .Z(G30) );
  XNOR2_X1 U745 ( .A(G143), .B(n669), .ZN(G45) );
  INV_X1 U746 ( .A(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n360), .A2(n671), .ZN(n672) );
  XNOR2_X1 U748 ( .A(n672), .B(KEYINPUT116), .ZN(n673) );
  XNOR2_X1 U749 ( .A(G146), .B(n673), .ZN(G48) );
  XOR2_X1 U750 ( .A(G113), .B(KEYINPUT117), .Z(n676) );
  NAND2_X1 U751 ( .A1(n678), .A2(n360), .ZN(n675) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(G15) );
  NAND2_X1 U753 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n679), .B(KEYINPUT118), .ZN(n680) );
  XNOR2_X1 U755 ( .A(G116), .B(n680), .ZN(G18) );
  XNOR2_X1 U756 ( .A(G134), .B(KEYINPUT120), .ZN(n682) );
  XNOR2_X1 U757 ( .A(n682), .B(n681), .ZN(G36) );
  XOR2_X1 U758 ( .A(G140), .B(n371), .Z(G42) );
  INV_X1 U759 ( .A(n685), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n358), .A2(n704), .ZN(n688) );
  NAND2_X1 U761 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n692), .B(KEYINPUT49), .ZN(n693) );
  NAND2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n699) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(KEYINPUT50), .ZN(n698) );
  NOR2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U768 ( .A(KEYINPUT121), .B(n700), .Z(n701) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT51), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n710), .B(KEYINPUT122), .ZN(n714) );
  NOR2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U777 ( .A(KEYINPUT123), .B(n715), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n717), .A2(n358), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U780 ( .A(n720), .B(KEYINPUT52), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n724), .B(KEYINPUT53), .ZN(G75) );
  BUF_X2 U782 ( .A(n731), .Z(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(G469), .ZN(n729) );
  BUF_X1 U784 ( .A(n725), .Z(n727) );
  XOR2_X1 U785 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n726) );
  NOR2_X1 U786 ( .A1(n741), .A2(n730), .ZN(G54) );
  NAND2_X1 U787 ( .A1(n731), .A2(G475), .ZN(n733) );
  XNOR2_X1 U788 ( .A(n733), .B(n379), .ZN(n735) );
  NAND2_X1 U789 ( .A1(G478), .A2(n738), .ZN(n736) );
  NAND2_X1 U790 ( .A1(G217), .A2(n738), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n752) );
  XOR2_X1 U792 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n745) );
  NAND2_X1 U793 ( .A1(G224), .A2(G953), .ZN(n744) );
  XNOR2_X1 U794 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U795 ( .A(KEYINPUT61), .B(n746), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n747), .A2(G898), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n748), .A2(n757), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(G69) );
  XOR2_X1 U800 ( .A(n753), .B(KEYINPUT96), .Z(n754) );
  XOR2_X1 U801 ( .A(n755), .B(n754), .Z(n759) );
  XOR2_X1 U802 ( .A(n759), .B(n756), .Z(n758) );
  NAND2_X1 U803 ( .A1(n758), .A2(n757), .ZN(n763) );
  XNOR2_X1 U804 ( .A(G227), .B(n759), .ZN(n760) );
  NAND2_X1 U805 ( .A1(n760), .A2(G900), .ZN(n761) );
  NAND2_X1 U806 ( .A1(n761), .A2(G953), .ZN(n762) );
  NAND2_X1 U807 ( .A1(n763), .A2(n762), .ZN(G72) );
  XOR2_X1 U808 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n766) );
  XNOR2_X1 U809 ( .A(n764), .B(G125), .ZN(n765) );
  XNOR2_X1 U810 ( .A(n766), .B(n765), .ZN(G27) );
  BUF_X1 U811 ( .A(n767), .Z(n768) );
  XNOR2_X1 U812 ( .A(G122), .B(n768), .ZN(G24) );
  XNOR2_X1 U813 ( .A(G131), .B(n769), .ZN(G33) );
  XNOR2_X1 U814 ( .A(G137), .B(n770), .ZN(G39) );
endmodule

