

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n675, n676, n677, n678, n680, n681, n682, n683, n684, n685,
         n686, n688, n689, n690, n691, n692, n693, n694, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805;

  BUF_X1 U371 ( .A(n769), .Z(n351) );
  INV_X1 U372 ( .A(n772), .ZN(n356) );
  INV_X1 U373 ( .A(n772), .ZN(n359) );
  INV_X1 U374 ( .A(n772), .ZN(n363) );
  INV_X1 U375 ( .A(n772), .ZN(n366) );
  INV_X1 U376 ( .A(n481), .ZN(n353) );
  NAND2_X1 U377 ( .A1(n779), .A2(n792), .ZN(n717) );
  NOR2_X1 U378 ( .A1(n608), .A2(n607), .ZN(n697) );
  NOR2_X1 U379 ( .A1(n805), .A2(n352), .ZN(n381) );
  NOR2_X1 U380 ( .A1(n440), .A2(n438), .ZN(n655) );
  INV_X1 U381 ( .A(n593), .ZN(n352) );
  AND2_X1 U382 ( .A1(n654), .A2(n380), .ZN(n436) );
  OR2_X1 U383 ( .A1(n670), .A2(G902), .ZN(n550) );
  XNOR2_X1 U384 ( .A(n565), .B(n371), .ZN(n718) );
  XNOR2_X1 U385 ( .A(n575), .B(n492), .ZN(n547) );
  BUF_X1 U386 ( .A(G104), .Z(n699) );
  XNOR2_X1 U387 ( .A(G128), .B(G119), .ZN(n551) );
  XNOR2_X1 U388 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n454) );
  INV_X1 U389 ( .A(G146), .ZN(n463) );
  AND2_X2 U390 ( .A1(n624), .A2(n623), .ZN(n652) );
  AND2_X1 U391 ( .A1(n357), .A2(n356), .ZN(n688) );
  AND2_X1 U392 ( .A1(n360), .A2(n359), .ZN(n681) );
  AND2_X1 U393 ( .A1(n364), .A2(n363), .ZN(n675) );
  AND2_X1 U394 ( .A1(n367), .A2(n366), .ZN(n696) );
  XNOR2_X1 U395 ( .A(n413), .B(n547), .ZN(n689) );
  XNOR2_X2 U396 ( .A(n597), .B(KEYINPUT31), .ZN(n710) );
  XNOR2_X2 U397 ( .A(KEYINPUT79), .B(n494), .ZN(n495) );
  XNOR2_X2 U398 ( .A(n425), .B(n424), .ZN(n805) );
  XNOR2_X2 U399 ( .A(n541), .B(KEYINPUT22), .ZN(n608) );
  XNOR2_X2 U400 ( .A(n621), .B(KEYINPUT1), .ZN(n581) );
  NAND2_X1 U401 ( .A1(n354), .A2(n353), .ZN(n485) );
  INV_X1 U402 ( .A(n717), .ZN(n354) );
  NAND2_X2 U403 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X2 U404 ( .A(KEYINPUT98), .B(n596), .Z(n734) );
  XNOR2_X2 U405 ( .A(n531), .B(KEYINPUT4), .ZN(n788) );
  NAND2_X1 U406 ( .A1(n355), .A2(n388), .ZN(n450) );
  AND2_X1 U407 ( .A1(n393), .A2(n392), .ZN(n355) );
  AND2_X2 U408 ( .A1(n600), .A2(n599), .ZN(n700) );
  XNOR2_X1 U409 ( .A(n686), .B(n358), .ZN(n357) );
  INV_X1 U410 ( .A(n685), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n678), .B(n361), .ZN(n360) );
  INV_X1 U412 ( .A(n677), .ZN(n361) );
  NAND2_X1 U413 ( .A1(n362), .A2(n374), .ZN(n773) );
  NAND2_X1 U414 ( .A1(n372), .A2(n373), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n672), .B(n365), .ZN(n364) );
  INV_X1 U416 ( .A(n671), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n694), .B(n368), .ZN(n367) );
  INV_X1 U418 ( .A(n693), .ZN(n368) );
  NOR2_X2 U419 ( .A1(n644), .A2(n643), .ZN(n484) );
  NAND2_X2 U420 ( .A1(n431), .A2(n383), .ZN(n666) );
  BUF_X2 U421 ( .A(n609), .Z(n649) );
  INV_X1 U422 ( .A(G119), .ZN(n429) );
  XNOR2_X1 U423 ( .A(G116), .B(G113), .ZN(n572) );
  INV_X1 U424 ( .A(G146), .ZN(n451) );
  INV_X2 U425 ( .A(G953), .ZN(n673) );
  XNOR2_X1 U426 ( .A(n396), .B(n377), .ZN(n376) );
  NAND2_X1 U427 ( .A1(n407), .A2(n408), .ZN(n721) );
  OR2_X1 U428 ( .A1(n676), .A2(n471), .ZN(n408) );
  XNOR2_X1 U429 ( .A(n626), .B(n625), .ZN(n657) );
  BUF_X1 U430 ( .A(n581), .Z(n728) );
  AND2_X1 U431 ( .A1(n603), .A2(n602), .ZN(n711) );
  INV_X1 U432 ( .A(KEYINPUT41), .ZN(n377) );
  NAND2_X1 U433 ( .A1(n707), .A2(n648), .ZN(n435) );
  BUF_X1 U434 ( .A(n700), .Z(n370) );
  NAND2_X1 U435 ( .A1(n657), .A2(n711), .ZN(n627) );
  XNOR2_X1 U436 ( .A(n581), .B(n423), .ZN(n640) );
  XNOR2_X1 U437 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U438 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U439 ( .A1(n614), .A2(n504), .ZN(n505) );
  AND2_X1 U440 ( .A1(n470), .A2(n472), .ZN(n407) );
  XNOR2_X1 U441 ( .A(n684), .B(KEYINPUT59), .ZN(n685) );
  XNOR2_X1 U442 ( .A(n676), .B(KEYINPUT62), .ZN(n677) );
  XNOR2_X1 U443 ( .A(n434), .B(n432), .ZN(n676) );
  XNOR2_X1 U444 ( .A(n486), .B(n566), .ZN(n371) );
  XNOR2_X1 U445 ( .A(n573), .B(n433), .ZN(n432) );
  XNOR2_X1 U446 ( .A(n789), .B(n463), .ZN(n574) );
  XNOR2_X1 U447 ( .A(n530), .B(n460), .ZN(n459) );
  NAND2_X1 U448 ( .A1(n497), .A2(G214), .ZN(n738) );
  XNOR2_X1 U449 ( .A(n451), .B(G125), .ZN(n508) );
  XNOR2_X1 U450 ( .A(n429), .B(KEYINPUT3), .ZN(n569) );
  XNOR2_X1 U451 ( .A(n464), .B(G134), .ZN(n789) );
  INV_X1 U452 ( .A(G116), .ZN(n461) );
  XNOR2_X1 U453 ( .A(G131), .B(KEYINPUT66), .ZN(n464) );
  XNOR2_X1 U454 ( .A(KEYINPUT97), .B(KEYINPUT23), .ZN(n553) );
  XNOR2_X1 U455 ( .A(G110), .B(KEYINPUT24), .ZN(n554) );
  NAND2_X1 U456 ( .A1(n369), .A2(n389), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n391), .A2(n381), .ZN(n369) );
  NAND2_X1 U458 ( .A1(n683), .A2(n802), .ZN(n629) );
  XNOR2_X2 U459 ( .A(n627), .B(KEYINPUT40), .ZN(n683) );
  NAND2_X1 U460 ( .A1(n462), .A2(n459), .ZN(n374) );
  INV_X1 U461 ( .A(n462), .ZN(n372) );
  INV_X1 U462 ( .A(n459), .ZN(n373) );
  XNOR2_X1 U463 ( .A(n490), .B(G122), .ZN(n507) );
  NOR2_X2 U464 ( .A1(G953), .A2(n760), .ZN(n761) );
  INV_X1 U465 ( .A(n376), .ZN(n754) );
  NOR2_X1 U466 ( .A1(n387), .A2(n697), .ZN(n393) );
  XNOR2_X2 U467 ( .A(n588), .B(KEYINPUT35), .ZN(n409) );
  NAND2_X1 U468 ( .A1(n405), .A2(n399), .ZN(n402) );
  AND2_X1 U469 ( .A1(n407), .A2(n631), .ZN(n399) );
  NAND2_X1 U470 ( .A1(n409), .A2(n449), .ZN(n391) );
  NAND2_X1 U471 ( .A1(n394), .A2(KEYINPUT83), .ZN(n392) );
  XNOR2_X1 U472 ( .A(n605), .B(KEYINPUT105), .ZN(n387) );
  XNOR2_X1 U473 ( .A(n422), .B(KEYINPUT106), .ZN(n577) );
  NAND2_X1 U474 ( .A1(n640), .A2(n567), .ZN(n422) );
  AND2_X1 U475 ( .A1(n408), .A2(n406), .ZN(n405) );
  NAND2_X1 U476 ( .A1(n407), .A2(n408), .ZN(n403) );
  XNOR2_X1 U477 ( .A(n417), .B(KEYINPUT99), .ZN(n604) );
  NAND2_X1 U478 ( .A1(n384), .A2(n457), .ZN(n389) );
  NAND2_X1 U479 ( .A1(n589), .A2(n385), .ZN(n384) );
  XNOR2_X1 U480 ( .A(n588), .B(n386), .ZN(n385) );
  NAND2_X1 U481 ( .A1(n403), .A2(n379), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n569), .B(n568), .ZN(n433) );
  XNOR2_X1 U483 ( .A(n461), .B(G107), .ZN(n530) );
  NOR2_X1 U484 ( .A1(G953), .A2(G237), .ZN(n570) );
  XOR2_X1 U485 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n512) );
  XNOR2_X1 U486 ( .A(n452), .B(n508), .ZN(n458) );
  XNOR2_X1 U487 ( .A(n454), .B(n453), .ZN(n452) );
  INV_X1 U488 ( .A(n664), .ZN(n480) );
  NAND2_X1 U489 ( .A1(G902), .A2(n474), .ZN(n472) );
  NAND2_X1 U490 ( .A1(n676), .A2(n474), .ZN(n470) );
  NAND2_X1 U491 ( .A1(n473), .A2(G472), .ZN(n471) );
  XNOR2_X1 U492 ( .A(n507), .B(n569), .ZN(n462) );
  INV_X1 U493 ( .A(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U494 ( .A(G134), .B(G122), .ZN(n526) );
  XOR2_X1 U495 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n527) );
  INV_X1 U496 ( .A(KEYINPUT77), .ZN(n428) );
  INV_X1 U497 ( .A(KEYINPUT30), .ZN(n415) );
  XNOR2_X1 U498 ( .A(n466), .B(n465), .ZN(n647) );
  INV_X1 U499 ( .A(KEYINPUT111), .ZN(n465) );
  INV_X1 U500 ( .A(n621), .ZN(n467) );
  AND2_X1 U501 ( .A1(n397), .A2(n719), .ZN(n539) );
  INV_X1 U502 ( .A(KEYINPUT47), .ZN(n445) );
  NOR2_X1 U503 ( .A1(n445), .A2(n648), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n803), .B(n418), .ZN(n643) );
  INV_X1 U505 ( .A(KEYINPUT82), .ZN(n418) );
  XNOR2_X1 U506 ( .A(KEYINPUT35), .B(KEYINPUT65), .ZN(n386) );
  INV_X1 U507 ( .A(KEYINPUT83), .ZN(n449) );
  INV_X1 U508 ( .A(G237), .ZN(n493) );
  XNOR2_X1 U509 ( .A(G902), .B(KEYINPUT15), .ZN(n664) );
  XNOR2_X1 U510 ( .A(n482), .B(n656), .ZN(n431) );
  INV_X1 U511 ( .A(KEYINPUT45), .ZN(n456) );
  INV_X1 U512 ( .A(G137), .ZN(n545) );
  NAND2_X1 U513 ( .A1(G234), .A2(G237), .ZN(n498) );
  XNOR2_X1 U514 ( .A(n618), .B(n469), .ZN(n468) );
  INV_X1 U515 ( .A(KEYINPUT28), .ZN(n469) );
  NAND2_X1 U516 ( .A1(n402), .A2(n401), .ZN(n617) );
  INV_X1 U517 ( .A(KEYINPUT88), .ZN(n491) );
  XOR2_X1 U518 ( .A(KEYINPUT102), .B(G140), .Z(n516) );
  XNOR2_X1 U519 ( .A(G143), .B(G131), .ZN(n515) );
  XNOR2_X1 U520 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n511) );
  XNOR2_X1 U521 ( .A(n773), .B(n414), .ZN(n413) );
  INV_X1 U522 ( .A(KEYINPUT64), .ZN(n479) );
  INV_X1 U523 ( .A(KEYINPUT86), .ZN(n423) );
  NAND2_X1 U524 ( .A1(n405), .A2(n407), .ZN(n404) );
  INV_X1 U525 ( .A(KEYINPUT95), .ZN(n448) );
  BUF_X1 U526 ( .A(n673), .Z(n793) );
  XNOR2_X1 U527 ( .A(n529), .B(n382), .ZN(n764) );
  XOR2_X1 U528 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n525) );
  NOR2_X1 U529 ( .A1(n793), .A2(G952), .ZN(n772) );
  OR2_X2 U530 ( .A1(n647), .A2(n376), .ZN(n395) );
  INV_X1 U531 ( .A(KEYINPUT32), .ZN(n424) );
  BUF_X1 U532 ( .A(n710), .Z(n713) );
  NOR2_X1 U533 ( .A1(n603), .A2(n602), .ZN(n378) );
  AND2_X1 U534 ( .A1(n631), .A2(KEYINPUT107), .ZN(n379) );
  INV_X1 U535 ( .A(G472), .ZN(n474) );
  AND2_X1 U536 ( .A1(n437), .A2(n439), .ZN(n380) );
  INV_X1 U537 ( .A(n743), .ZN(n447) );
  XOR2_X1 U538 ( .A(n532), .B(n528), .Z(n382) );
  INV_X1 U539 ( .A(n741), .ZN(n397) );
  AND2_X1 U540 ( .A1(n682), .A2(n715), .ZN(n383) );
  INV_X1 U541 ( .A(KEYINPUT107), .ZN(n406) );
  INV_X1 U542 ( .A(KEYINPUT2), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n409), .A2(KEYINPUT44), .ZN(n394) );
  XNOR2_X1 U544 ( .A(n575), .B(n574), .ZN(n434) );
  XNOR2_X2 U545 ( .A(n788), .B(G101), .ZN(n575) );
  XNOR2_X2 U546 ( .A(G143), .B(G128), .ZN(n531) );
  XNOR2_X2 U547 ( .A(n395), .B(KEYINPUT42), .ZN(n802) );
  NAND2_X1 U548 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U549 ( .A(n742), .ZN(n398) );
  NAND2_X1 U550 ( .A1(n400), .A2(n404), .ZN(n619) );
  NAND2_X1 U551 ( .A1(n403), .A2(KEYINPUT107), .ZN(n400) );
  BUF_X1 U552 ( .A(n773), .Z(n410) );
  NAND2_X1 U553 ( .A1(n739), .A2(n652), .ZN(n626) );
  NAND2_X2 U554 ( .A1(n411), .A2(n587), .ZN(n588) );
  XNOR2_X2 U555 ( .A(n412), .B(n586), .ZN(n411) );
  NAND2_X1 U556 ( .A1(n600), .A2(n753), .ZN(n412) );
  XNOR2_X1 U557 ( .A(n540), .B(n448), .ZN(n600) );
  NAND2_X1 U558 ( .A1(n689), .A2(n664), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n458), .B(n489), .ZN(n414) );
  INV_X1 U560 ( .A(KEYINPUT44), .ZN(n457) );
  XNOR2_X1 U561 ( .A(n416), .B(n415), .ZN(n624) );
  NAND2_X1 U562 ( .A1(n619), .A2(n738), .ZN(n416) );
  NOR2_X2 U563 ( .A1(n710), .A2(n700), .ZN(n417) );
  XNOR2_X1 U564 ( .A(n547), .B(n419), .ZN(n670) );
  XNOR2_X1 U565 ( .A(n420), .B(n574), .ZN(n419) );
  XNOR2_X1 U566 ( .A(n546), .B(n421), .ZN(n420) );
  INV_X1 U567 ( .A(n562), .ZN(n421) );
  NAND2_X1 U568 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U569 ( .A(n608), .ZN(n426) );
  XNOR2_X1 U570 ( .A(n578), .B(n428), .ZN(n427) );
  NAND2_X1 U571 ( .A1(n430), .A2(n481), .ZN(n478) );
  XNOR2_X1 U572 ( .A(n666), .B(KEYINPUT74), .ZN(n430) );
  NAND2_X1 U573 ( .A1(n436), .A2(n435), .ZN(n438) );
  NAND2_X1 U574 ( .A1(n743), .A2(n648), .ZN(n437) );
  NAND2_X1 U575 ( .A1(n445), .A2(n648), .ZN(n439) );
  NAND2_X1 U576 ( .A1(n443), .A2(n441), .ZN(n440) );
  NAND2_X1 U577 ( .A1(n446), .A2(n442), .ZN(n441) );
  NAND2_X1 U578 ( .A1(n444), .A2(n445), .ZN(n443) );
  INV_X1 U579 ( .A(n446), .ZN(n444) );
  NAND2_X1 U580 ( .A1(n707), .A2(n447), .ZN(n446) );
  XNOR2_X2 U581 ( .A(n506), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X2 U582 ( .A(n450), .B(n456), .ZN(n665) );
  XNOR2_X2 U583 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n453) );
  NAND2_X1 U584 ( .A1(n609), .A2(n738), .ZN(n455) );
  XNOR2_X2 U585 ( .A(n635), .B(KEYINPUT19), .ZN(n645) );
  XNOR2_X2 U586 ( .A(n455), .B(KEYINPUT85), .ZN(n635) );
  XNOR2_X2 U587 ( .A(n496), .B(n495), .ZN(n609) );
  NOR2_X1 U588 ( .A1(n704), .A2(n805), .ZN(n589) );
  NOR2_X2 U589 ( .A1(n647), .A2(n646), .ZN(n707) );
  NAND2_X1 U590 ( .A1(n468), .A2(n467), .ZN(n466) );
  INV_X1 U591 ( .A(G902), .ZN(n473) );
  XNOR2_X1 U592 ( .A(n475), .B(n479), .ZN(n667) );
  NAND2_X1 U593 ( .A1(n477), .A2(n476), .ZN(n475) );
  NAND2_X1 U594 ( .A1(n665), .A2(n481), .ZN(n476) );
  AND2_X1 U595 ( .A1(n478), .A2(n480), .ZN(n477) );
  NAND2_X1 U596 ( .A1(n484), .A2(n483), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n655), .B(KEYINPUT72), .ZN(n483) );
  BUF_X1 U598 ( .A(n763), .Z(n768) );
  AND2_X1 U599 ( .A1(n564), .A2(G217), .ZN(n486) );
  BUF_X1 U600 ( .A(n689), .Z(n692) );
  INV_X1 U601 ( .A(n666), .ZN(n792) );
  XOR2_X1 U602 ( .A(KEYINPUT89), .B(KEYINPUT76), .Z(n488) );
  NAND2_X1 U603 ( .A1(G224), .A2(n673), .ZN(n487) );
  XNOR2_X1 U604 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X2 U605 ( .A(G113), .B(G104), .ZN(n490) );
  XNOR2_X1 U606 ( .A(n491), .B(G110), .ZN(n774) );
  XNOR2_X1 U607 ( .A(n774), .B(KEYINPUT69), .ZN(n492) );
  NAND2_X1 U608 ( .A1(n473), .A2(n493), .ZN(n497) );
  NAND2_X1 U609 ( .A1(G210), .A2(n497), .ZN(n494) );
  XNOR2_X1 U610 ( .A(n498), .B(KEYINPUT14), .ZN(n500) );
  NAND2_X1 U611 ( .A1(n500), .A2(G952), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n499), .B(KEYINPUT92), .ZN(n752) );
  NOR2_X1 U613 ( .A1(n752), .A2(G953), .ZN(n614) );
  NAND2_X1 U614 ( .A1(G902), .A2(n500), .ZN(n501) );
  XNOR2_X1 U615 ( .A(KEYINPUT93), .B(n501), .ZN(n502) );
  NAND2_X1 U616 ( .A1(n502), .A2(G953), .ZN(n611) );
  NOR2_X1 U617 ( .A1(G898), .A2(n611), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n503), .B(KEYINPUT94), .ZN(n504) );
  NOR2_X2 U619 ( .A1(n645), .A2(n505), .ZN(n506) );
  BUF_X1 U620 ( .A(n507), .Z(n510) );
  XNOR2_X1 U621 ( .A(n508), .B(KEYINPUT10), .ZN(n561) );
  INV_X1 U622 ( .A(n561), .ZN(n509) );
  XOR2_X1 U623 ( .A(n510), .B(n509), .Z(n520) );
  XNOR2_X1 U624 ( .A(n512), .B(n511), .ZN(n514) );
  NAND2_X1 U625 ( .A1(G214), .A2(n570), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U627 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U628 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n520), .B(n519), .ZN(n684) );
  NAND2_X1 U630 ( .A1(n684), .A2(n473), .ZN(n522) );
  XNOR2_X1 U631 ( .A(KEYINPUT13), .B(G475), .ZN(n521) );
  XNOR2_X1 U632 ( .A(n522), .B(n521), .ZN(n601) );
  NAND2_X1 U633 ( .A1(G234), .A2(n673), .ZN(n523) );
  XOR2_X1 U634 ( .A(KEYINPUT8), .B(n523), .Z(n558) );
  NAND2_X1 U635 ( .A1(G217), .A2(n558), .ZN(n524) );
  XNOR2_X1 U636 ( .A(n525), .B(n524), .ZN(n529) );
  XNOR2_X1 U637 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U639 ( .A1(n764), .A2(n473), .ZN(n534) );
  INV_X1 U640 ( .A(G478), .ZN(n533) );
  XNOR2_X1 U641 ( .A(n534), .B(n533), .ZN(n602) );
  NAND2_X1 U642 ( .A1(n601), .A2(n602), .ZN(n741) );
  NAND2_X1 U643 ( .A1(G234), .A2(n664), .ZN(n535) );
  XNOR2_X1 U644 ( .A(KEYINPUT20), .B(n535), .ZN(n564) );
  NAND2_X1 U645 ( .A1(n564), .A2(G221), .ZN(n537) );
  INV_X1 U646 ( .A(KEYINPUT21), .ZN(n536) );
  XNOR2_X1 U647 ( .A(n537), .B(n536), .ZN(n719) );
  INV_X1 U648 ( .A(n719), .ZN(n538) );
  NAND2_X1 U649 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U650 ( .A1(n673), .A2(G227), .ZN(n542) );
  XNOR2_X1 U651 ( .A(n542), .B(KEYINPUT96), .ZN(n544) );
  XNOR2_X1 U652 ( .A(G107), .B(n699), .ZN(n543) );
  XNOR2_X1 U653 ( .A(n544), .B(n543), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n545), .B(G140), .ZN(n562) );
  INV_X1 U655 ( .A(KEYINPUT68), .ZN(n548) );
  XNOR2_X1 U656 ( .A(n548), .B(G469), .ZN(n549) );
  XNOR2_X2 U657 ( .A(n550), .B(n549), .ZN(n621) );
  XNOR2_X1 U658 ( .A(n551), .B(KEYINPUT75), .ZN(n552) );
  INV_X1 U659 ( .A(n552), .ZN(n557) );
  INV_X1 U660 ( .A(n553), .ZN(n555) );
  XNOR2_X1 U661 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U662 ( .A(n556), .B(n557), .ZN(n560) );
  NAND2_X1 U663 ( .A1(G221), .A2(n558), .ZN(n559) );
  XNOR2_X1 U664 ( .A(n560), .B(n559), .ZN(n563) );
  XNOR2_X1 U665 ( .A(n562), .B(n561), .ZN(n787) );
  XNOR2_X1 U666 ( .A(n563), .B(n787), .ZN(n769) );
  NOR2_X1 U667 ( .A1(n769), .A2(G902), .ZN(n565) );
  INV_X1 U668 ( .A(KEYINPUT25), .ZN(n566) );
  INV_X1 U669 ( .A(n718), .ZN(n567) );
  XNOR2_X1 U670 ( .A(KEYINPUT5), .B(G137), .ZN(n568) );
  NAND2_X1 U671 ( .A1(G210), .A2(n570), .ZN(n571) );
  XNOR2_X1 U672 ( .A(n572), .B(n571), .ZN(n573) );
  INV_X1 U673 ( .A(n721), .ZN(n594) );
  XNOR2_X1 U674 ( .A(n594), .B(KEYINPUT6), .ZN(n633) );
  XOR2_X1 U675 ( .A(KEYINPUT78), .B(n633), .Z(n576) );
  NOR2_X1 U676 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U677 ( .A1(n619), .A2(n718), .ZN(n579) );
  NAND2_X1 U678 ( .A1(n728), .A2(n579), .ZN(n580) );
  NOR2_X1 U679 ( .A1(n608), .A2(n580), .ZN(n704) );
  INV_X1 U680 ( .A(n581), .ZN(n582) );
  AND2_X1 U681 ( .A1(n718), .A2(n719), .ZN(n726) );
  AND2_X1 U682 ( .A1(n582), .A2(n726), .ZN(n595) );
  INV_X1 U683 ( .A(n633), .ZN(n583) );
  NAND2_X1 U684 ( .A1(n595), .A2(n583), .ZN(n585) );
  XNOR2_X1 U685 ( .A(KEYINPUT70), .B(KEYINPUT33), .ZN(n584) );
  XNOR2_X1 U686 ( .A(n585), .B(n584), .ZN(n753) );
  INV_X1 U687 ( .A(KEYINPUT34), .ZN(n586) );
  OR2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n650) );
  INV_X1 U689 ( .A(n650), .ZN(n587) );
  INV_X1 U690 ( .A(KEYINPUT65), .ZN(n590) );
  NAND2_X1 U691 ( .A1(n590), .A2(KEYINPUT44), .ZN(n591) );
  NOR2_X1 U692 ( .A1(n704), .A2(n591), .ZN(n593) );
  NAND2_X1 U693 ( .A1(n540), .A2(n734), .ZN(n597) );
  NAND2_X1 U694 ( .A1(n726), .A2(n721), .ZN(n598) );
  NOR2_X1 U695 ( .A1(n598), .A2(n621), .ZN(n599) );
  INV_X1 U696 ( .A(n601), .ZN(n603) );
  NOR2_X1 U697 ( .A1(n711), .A2(n378), .ZN(n743) );
  NAND2_X1 U698 ( .A1(n604), .A2(n447), .ZN(n605) );
  AND2_X1 U699 ( .A1(n633), .A2(n718), .ZN(n606) );
  NAND2_X1 U700 ( .A1(n728), .A2(n606), .ZN(n607) );
  XNOR2_X1 U701 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n610) );
  XNOR2_X2 U702 ( .A(n649), .B(n610), .ZN(n739) );
  NAND2_X1 U703 ( .A1(n739), .A2(n738), .ZN(n742) );
  NOR2_X1 U704 ( .A1(n718), .A2(n538), .ZN(n630) );
  XNOR2_X1 U705 ( .A(KEYINPUT108), .B(n611), .ZN(n612) );
  NOR2_X1 U706 ( .A1(G900), .A2(n612), .ZN(n613) );
  XNOR2_X1 U707 ( .A(n613), .B(KEYINPUT109), .ZN(n616) );
  INV_X1 U708 ( .A(n614), .ZN(n615) );
  NAND2_X1 U709 ( .A1(n616), .A2(n615), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n630), .A2(n617), .ZN(n618) );
  INV_X1 U711 ( .A(n631), .ZN(n620) );
  NOR2_X1 U712 ( .A1(n621), .A2(n620), .ZN(n622) );
  AND2_X1 U713 ( .A1(n726), .A2(n622), .ZN(n623) );
  XOR2_X1 U714 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n625) );
  XOR2_X1 U715 ( .A(KEYINPUT81), .B(KEYINPUT46), .Z(n628) );
  XNOR2_X1 U716 ( .A(n629), .B(n628), .ZN(n644) );
  AND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n711), .A2(n632), .ZN(n634) );
  OR2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n659) );
  INV_X1 U720 ( .A(n659), .ZN(n637) );
  BUF_X1 U721 ( .A(n635), .Z(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT36), .B(KEYINPUT84), .Z(n638) );
  XNOR2_X1 U724 ( .A(n639), .B(n638), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U726 ( .A(n642), .B(KEYINPUT112), .ZN(n803) );
  BUF_X1 U727 ( .A(n645), .Z(n646) );
  INV_X1 U728 ( .A(KEYINPUT80), .ZN(n648) );
  INV_X1 U729 ( .A(n649), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n662), .A2(n650), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U732 ( .A(KEYINPUT110), .B(n653), .Z(n801) );
  INV_X1 U733 ( .A(n801), .ZN(n654) );
  XNOR2_X1 U734 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n657), .A2(n378), .ZN(n682) );
  INV_X1 U736 ( .A(n738), .ZN(n658) );
  NOR2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n660), .A2(n728), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT43), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n715) );
  INV_X1 U741 ( .A(n665), .ZN(n779) );
  AND2_X2 U742 ( .A1(n667), .A2(n485), .ZN(n763) );
  NAND2_X1 U743 ( .A1(n763), .A2(G469), .ZN(n672) );
  XNOR2_X1 U744 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(KEYINPUT57), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n763), .A2(G472), .ZN(n678) );
  XNOR2_X1 U748 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(G57) );
  XNOR2_X1 U750 ( .A(n682), .B(G134), .ZN(G36) );
  XNOR2_X1 U751 ( .A(n683), .B(G131), .ZN(G33) );
  NAND2_X1 U752 ( .A1(n763), .A2(G475), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n688), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U754 ( .A1(n763), .A2(G210), .ZN(n694) );
  XNOR2_X1 U755 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT55), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U758 ( .A(n409), .B(G122), .Z(G24) );
  XOR2_X1 U759 ( .A(G101), .B(n697), .Z(G3) );
  NAND2_X1 U760 ( .A1(n370), .A2(n711), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n699), .B(n698), .ZN(G6) );
  XOR2_X1 U762 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U763 ( .A1(n370), .A2(n378), .ZN(n701) );
  XNOR2_X1 U764 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(G107), .B(n703), .ZN(G9) );
  XOR2_X1 U766 ( .A(G110), .B(n704), .Z(G12) );
  XOR2_X1 U767 ( .A(G128), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U768 ( .A1(n378), .A2(n707), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n706), .B(n705), .ZN(G30) );
  XOR2_X1 U770 ( .A(G146), .B(KEYINPUT113), .Z(n709) );
  NAND2_X1 U771 ( .A1(n707), .A2(n711), .ZN(n708) );
  XNOR2_X1 U772 ( .A(n709), .B(n708), .ZN(G48) );
  NAND2_X1 U773 ( .A1(n713), .A2(n711), .ZN(n712) );
  XNOR2_X1 U774 ( .A(n712), .B(G113), .ZN(G15) );
  NAND2_X1 U775 ( .A1(n713), .A2(n378), .ZN(n714) );
  XNOR2_X1 U776 ( .A(n714), .B(G116), .ZN(G18) );
  XNOR2_X1 U777 ( .A(G140), .B(KEYINPUT114), .ZN(n716) );
  XNOR2_X1 U778 ( .A(n716), .B(n715), .ZN(G42) );
  XNOR2_X1 U779 ( .A(n717), .B(n481), .ZN(n759) );
  NOR2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U781 ( .A(KEYINPUT49), .B(n720), .ZN(n722) );
  AND2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n732) );
  INV_X1 U783 ( .A(n726), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n728), .A2(n723), .ZN(n724) );
  XOR2_X1 U785 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n725) );
  NAND2_X1 U786 ( .A1(n724), .A2(n725), .ZN(n730) );
  NOR2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n735), .B(KEYINPUT116), .ZN(n736) );
  XNOR2_X1 U793 ( .A(n736), .B(KEYINPUT51), .ZN(n737) );
  NAND2_X1 U794 ( .A1(n737), .A2(n754), .ZN(n749) );
  NOR2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U796 ( .A1(n741), .A2(n740), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U798 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U799 ( .A(KEYINPUT117), .B(n746), .ZN(n747) );
  NAND2_X1 U800 ( .A1(n747), .A2(n753), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U802 ( .A(KEYINPUT52), .B(n750), .Z(n751) );
  NOR2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U805 ( .A(n755), .B(KEYINPUT118), .Z(n756) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U808 ( .A(KEYINPUT53), .B(n761), .Z(n762) );
  XNOR2_X1 U809 ( .A(KEYINPUT119), .B(n762), .ZN(G75) );
  NAND2_X1 U810 ( .A1(n768), .A2(G478), .ZN(n766) );
  XNOR2_X1 U811 ( .A(n764), .B(KEYINPUT123), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U813 ( .A1(n772), .A2(n767), .ZN(G63) );
  NAND2_X1 U814 ( .A1(n768), .A2(G217), .ZN(n770) );
  XNOR2_X1 U815 ( .A(n351), .B(n770), .ZN(n771) );
  NOR2_X1 U816 ( .A1(n772), .A2(n771), .ZN(G66) );
  XOR2_X1 U817 ( .A(KEYINPUT125), .B(n410), .Z(n776) );
  XNOR2_X1 U818 ( .A(G101), .B(n774), .ZN(n775) );
  XNOR2_X1 U819 ( .A(n776), .B(n775), .ZN(n778) );
  NOR2_X1 U820 ( .A1(G898), .A2(n793), .ZN(n777) );
  NOR2_X1 U821 ( .A1(n778), .A2(n777), .ZN(n786) );
  NAND2_X1 U822 ( .A1(n779), .A2(n793), .ZN(n784) );
  NAND2_X1 U823 ( .A1(G224), .A2(G953), .ZN(n780) );
  XNOR2_X1 U824 ( .A(n780), .B(KEYINPUT124), .ZN(n781) );
  XNOR2_X1 U825 ( .A(KEYINPUT61), .B(n781), .ZN(n782) );
  NAND2_X1 U826 ( .A1(G898), .A2(n782), .ZN(n783) );
  NAND2_X1 U827 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U828 ( .A(n786), .B(n785), .ZN(G69) );
  XOR2_X1 U829 ( .A(n787), .B(KEYINPUT126), .Z(n791) );
  XOR2_X1 U830 ( .A(n789), .B(n788), .Z(n790) );
  XNOR2_X1 U831 ( .A(n791), .B(n790), .ZN(n795) );
  XNOR2_X1 U832 ( .A(n792), .B(n795), .ZN(n794) );
  NAND2_X1 U833 ( .A1(n794), .A2(n793), .ZN(n800) );
  XNOR2_X1 U834 ( .A(n795), .B(G227), .ZN(n796) );
  XNOR2_X1 U835 ( .A(n796), .B(KEYINPUT127), .ZN(n797) );
  NAND2_X1 U836 ( .A1(n797), .A2(G900), .ZN(n798) );
  NAND2_X1 U837 ( .A1(n798), .A2(G953), .ZN(n799) );
  NAND2_X1 U838 ( .A1(n800), .A2(n799), .ZN(G72) );
  XOR2_X1 U839 ( .A(n801), .B(G143), .Z(G45) );
  XNOR2_X1 U840 ( .A(n802), .B(G137), .ZN(G39) );
  XOR2_X1 U841 ( .A(G125), .B(n803), .Z(n804) );
  XNOR2_X1 U842 ( .A(KEYINPUT37), .B(n804), .ZN(G27) );
  XOR2_X1 U843 ( .A(n805), .B(G119), .Z(G21) );
endmodule

