

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U547 ( .A1(n673), .A2(n671), .ZN(n655) );
  NOR2_X1 U548 ( .A1(n657), .A2(n654), .ZN(n592) );
  NOR2_X2 U549 ( .A1(n596), .A2(G168), .ZN(n597) );
  AND2_X1 U550 ( .A1(n743), .A2(n510), .ZN(n745) );
  XNOR2_X2 U551 ( .A(n585), .B(KEYINPUT85), .ZN(n711) );
  XNOR2_X2 U552 ( .A(n528), .B(KEYINPUT65), .ZN(n577) );
  XNOR2_X1 U553 ( .A(KEYINPUT31), .B(n604), .ZN(n673) );
  XNOR2_X1 U554 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n679) );
  INV_X1 U555 ( .A(KEYINPUT23), .ZN(n578) );
  AND2_X1 U556 ( .A1(n751), .A2(n742), .ZN(n510) );
  AND2_X1 U557 ( .A1(n626), .A2(n625), .ZN(n511) );
  XOR2_X1 U558 ( .A(KEYINPUT67), .B(n575), .Z(n512) );
  XOR2_X1 U559 ( .A(KEYINPUT29), .B(n652), .Z(n513) );
  INV_X1 U560 ( .A(n1007), .ZN(n625) );
  AND2_X1 U561 ( .A1(n627), .A2(n511), .ZN(n628) );
  INV_X1 U562 ( .A(KEYINPUT95), .ZN(n591) );
  INV_X1 U563 ( .A(KEYINPUT91), .ZN(n587) );
  XNOR2_X1 U564 ( .A(n588), .B(n587), .ZN(n657) );
  INV_X1 U565 ( .A(KEYINPUT89), .ZN(n589) );
  XNOR2_X1 U566 ( .A(n680), .B(n679), .ZN(n697) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n530) );
  INV_X1 U568 ( .A(KEYINPUT102), .ZN(n744) );
  NOR2_X2 U569 ( .A1(G2104), .A2(n534), .ZN(n903) );
  AND2_X2 U570 ( .A1(G2105), .A2(G2104), .ZN(n904) );
  NOR2_X1 U571 ( .A1(G651), .A2(n551), .ZN(n800) );
  XNOR2_X1 U572 ( .A(n759), .B(KEYINPUT40), .ZN(n760) );
  NOR2_X2 U573 ( .A1(G651), .A2(G543), .ZN(n807) );
  NAND2_X1 U574 ( .A1(G89), .A2(n807), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n514), .B(KEYINPUT72), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n515), .B(KEYINPUT4), .ZN(n517) );
  XOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .Z(n551) );
  INV_X1 U578 ( .A(G651), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n551), .A2(n519), .ZN(n802) );
  NAND2_X1 U580 ( .A1(G76), .A2(n802), .ZN(n516) );
  NAND2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT5), .ZN(n525) );
  NOR2_X1 U583 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n520), .Z(n806) );
  NAND2_X1 U585 ( .A1(G63), .A2(n806), .ZN(n522) );
  NAND2_X1 U586 ( .A1(G51), .A2(n800), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(n523), .Z(n524) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U591 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U592 ( .A1(n527), .A2(G2104), .ZN(n528) );
  INV_X1 U593 ( .A(n577), .ZN(n529) );
  INV_X1 U594 ( .A(n529), .ZN(n898) );
  NAND2_X1 U595 ( .A1(G102), .A2(n898), .ZN(n533) );
  NOR2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XNOR2_X2 U597 ( .A(n531), .B(n530), .ZN(n899) );
  NAND2_X1 U598 ( .A1(G138), .A2(n899), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n538) );
  INV_X1 U600 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U601 ( .A1(G126), .A2(n903), .ZN(n536) );
  NAND2_X1 U602 ( .A1(G114), .A2(n904), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G64), .A2(n806), .ZN(n540) );
  NAND2_X1 U606 ( .A1(G52), .A2(n800), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U608 ( .A1(G77), .A2(n802), .ZN(n542) );
  NAND2_X1 U609 ( .A1(G90), .A2(n807), .ZN(n541) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT70), .B(n546), .ZN(G171) );
  NAND2_X1 U614 ( .A1(G49), .A2(n800), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G74), .A2(G651), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U617 ( .A1(n806), .A2(n549), .ZN(n550) );
  XOR2_X1 U618 ( .A(KEYINPUT79), .B(n550), .Z(n553) );
  NAND2_X1 U619 ( .A1(n551), .A2(G87), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(G288) );
  NAND2_X1 U621 ( .A1(G75), .A2(n802), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G88), .A2(n807), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G62), .A2(n806), .ZN(n557) );
  NAND2_X1 U625 ( .A1(G50), .A2(n800), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(G166) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G61), .A2(n806), .ZN(n561) );
  NAND2_X1 U631 ( .A1(G86), .A2(n807), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n802), .A2(G73), .ZN(n562) );
  XOR2_X1 U634 ( .A(KEYINPUT2), .B(n562), .Z(n563) );
  NOR2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n800), .A2(G48), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n566), .A2(n565), .ZN(G305) );
  NAND2_X1 U638 ( .A1(G60), .A2(n806), .ZN(n568) );
  NAND2_X1 U639 ( .A1(G47), .A2(n800), .ZN(n567) );
  NAND2_X1 U640 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U641 ( .A(KEYINPUT69), .B(n569), .Z(n572) );
  NAND2_X1 U642 ( .A1(G72), .A2(n802), .ZN(n570) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(n570), .Z(n571) );
  NOR2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n807), .A2(G85), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(G290) );
  NAND2_X1 U647 ( .A1(G113), .A2(n904), .ZN(n575) );
  AND2_X1 U648 ( .A1(G40), .A2(n512), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n899), .A2(G137), .ZN(n762) );
  AND2_X1 U650 ( .A1(n576), .A2(n762), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n577), .A2(G101), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n579), .B(n578), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n903), .A2(G125), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U655 ( .A(KEYINPUT66), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n583), .B(n582), .ZN(n763) );
  NAND2_X1 U657 ( .A1(n584), .A2(n763), .ZN(n585) );
  NOR2_X1 U658 ( .A1(G164), .A2(G1384), .ZN(n710) );
  NAND2_X1 U659 ( .A1(n711), .A2(n710), .ZN(n586) );
  XNOR2_X2 U660 ( .A(n586), .B(KEYINPUT64), .ZN(n598) );
  BUF_X2 U661 ( .A(n598), .Z(n665) );
  NOR2_X1 U662 ( .A1(n665), .A2(G2084), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n598), .A2(G8), .ZN(n590) );
  XNOR2_X2 U664 ( .A(n590), .B(n589), .ZN(n660) );
  NOR2_X2 U665 ( .A1(G1966), .A2(n660), .ZN(n654) );
  XNOR2_X1 U666 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n593), .A2(G8), .ZN(n595) );
  XNOR2_X1 U668 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n597), .B(KEYINPUT97), .ZN(n603) );
  INV_X1 U671 ( .A(n598), .ZN(n613) );
  NOR2_X1 U672 ( .A1(G1961), .A2(n613), .ZN(n600) );
  XOR2_X1 U673 ( .A(G2078), .B(KEYINPUT25), .Z(n954) );
  NOR2_X1 U674 ( .A1(n665), .A2(n954), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U676 ( .A(KEYINPUT92), .B(n601), .Z(n605) );
  OR2_X1 U677 ( .A1(G171), .A2(n605), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G171), .A2(n605), .ZN(n653) );
  NAND2_X1 U680 ( .A1(G66), .A2(n806), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G92), .A2(n807), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G54), .A2(n800), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G79), .A2(n802), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U687 ( .A(KEYINPUT15), .B(n612), .Z(n849) );
  AND2_X1 U688 ( .A1(n613), .A2(G1996), .ZN(n614) );
  XOR2_X1 U689 ( .A(n614), .B(KEYINPUT26), .Z(n627) );
  NAND2_X1 U690 ( .A1(n665), .A2(G1341), .ZN(n626) );
  NAND2_X1 U691 ( .A1(G56), .A2(n806), .ZN(n615) );
  XOR2_X1 U692 ( .A(KEYINPUT14), .B(n615), .Z(n622) );
  NAND2_X1 U693 ( .A1(G81), .A2(n807), .ZN(n616) );
  XOR2_X1 U694 ( .A(KEYINPUT12), .B(n616), .Z(n617) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT71), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G68), .A2(n802), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT13), .B(n620), .Z(n621) );
  NOR2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n800), .A2(G43), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n1007) );
  OR2_X1 U702 ( .A1(n849), .A2(n628), .ZN(n635) );
  NAND2_X1 U703 ( .A1(n849), .A2(n628), .ZN(n633) );
  AND2_X1 U704 ( .A1(n613), .A2(G2067), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n629), .B(KEYINPUT93), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n665), .A2(G1348), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT94), .ZN(n647) );
  NAND2_X1 U711 ( .A1(G2072), .A2(n613), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n637), .B(KEYINPUT27), .ZN(n639) );
  INV_X1 U713 ( .A(G1956), .ZN(n1002) );
  NOR2_X1 U714 ( .A1(n613), .A2(n1002), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n648) );
  NAND2_X1 U716 ( .A1(G65), .A2(n806), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G53), .A2(n800), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G78), .A2(n802), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G91), .A2(n807), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n1003) );
  NAND2_X1 U723 ( .A1(n648), .A2(n1003), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n648), .A2(n1003), .ZN(n649) );
  XOR2_X1 U726 ( .A(n649), .B(KEYINPUT28), .Z(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n513), .ZN(n671) );
  NOR2_X2 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT98), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n657), .A2(G8), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n696) );
  NAND2_X1 U733 ( .A1(G1976), .A2(G288), .ZN(n1010) );
  INV_X1 U734 ( .A(n1010), .ZN(n662) );
  BUF_X1 U735 ( .A(n660), .Z(n661) );
  OR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n687) );
  INV_X1 U737 ( .A(n687), .ZN(n663) );
  AND2_X1 U738 ( .A1(n696), .A2(n663), .ZN(n684) );
  INV_X1 U739 ( .A(G8), .ZN(n670) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n661), .ZN(n664) );
  XNOR2_X1 U741 ( .A(KEYINPUT99), .B(n664), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n665), .A2(G2090), .ZN(n666) );
  NOR2_X1 U743 ( .A1(G166), .A2(n666), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n668), .A2(n667), .ZN(n669) );
  OR2_X1 U745 ( .A1(n670), .A2(n669), .ZN(n674) );
  AND2_X1 U746 ( .A1(n671), .A2(n674), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n678) );
  INV_X1 U748 ( .A(n674), .ZN(n676) );
  AND2_X1 U749 ( .A1(G286), .A2(G8), .ZN(n675) );
  OR2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n680) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n686), .A2(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U754 ( .A1(n661), .A2(n681), .ZN(n691) );
  INV_X1 U755 ( .A(n691), .ZN(n682) );
  AND2_X1 U756 ( .A1(n697), .A2(n682), .ZN(n683) );
  NAND2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n693) );
  INV_X1 U758 ( .A(KEYINPUT33), .ZN(n689) );
  NOR2_X1 U759 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U760 ( .A1(n686), .A2(n685), .ZN(n1017) );
  OR2_X1 U761 ( .A1(n687), .A2(n1017), .ZN(n688) );
  AND2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  OR2_X1 U763 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U765 ( .A(G1981), .B(G305), .Z(n1020) );
  NAND2_X1 U766 ( .A1(n694), .A2(n1020), .ZN(n702) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U768 ( .A1(G8), .A2(n695), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n700), .A2(n661), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U773 ( .A(n703), .B(KEYINPUT101), .ZN(n709) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XNOR2_X1 U775 ( .A(n704), .B(KEYINPUT24), .ZN(n705) );
  XNOR2_X1 U776 ( .A(n705), .B(KEYINPUT90), .ZN(n707) );
  INV_X1 U777 ( .A(n661), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n743) );
  INV_X1 U780 ( .A(n710), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n739) );
  INV_X1 U782 ( .A(n739), .ZN(n755) );
  NAND2_X1 U783 ( .A1(G104), .A2(n898), .ZN(n714) );
  NAND2_X1 U784 ( .A1(G140), .A2(n899), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U786 ( .A(KEYINPUT34), .B(n715), .ZN(n720) );
  NAND2_X1 U787 ( .A1(G128), .A2(n903), .ZN(n717) );
  NAND2_X1 U788 ( .A1(G116), .A2(n904), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U790 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U792 ( .A(KEYINPUT36), .B(n721), .ZN(n913) );
  XNOR2_X1 U793 ( .A(KEYINPUT37), .B(G2067), .ZN(n753) );
  NOR2_X1 U794 ( .A1(n913), .A2(n753), .ZN(n923) );
  NAND2_X1 U795 ( .A1(n755), .A2(n923), .ZN(n751) );
  NAND2_X1 U796 ( .A1(G119), .A2(n903), .ZN(n723) );
  NAND2_X1 U797 ( .A1(G107), .A2(n904), .ZN(n722) );
  NAND2_X1 U798 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G95), .A2(n898), .ZN(n725) );
  NAND2_X1 U800 ( .A1(G131), .A2(n899), .ZN(n724) );
  NAND2_X1 U801 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n910) );
  INV_X1 U803 ( .A(G1991), .ZN(n952) );
  NOR2_X1 U804 ( .A1(n910), .A2(n952), .ZN(n738) );
  NAND2_X1 U805 ( .A1(G105), .A2(n898), .ZN(n728) );
  XNOR2_X1 U806 ( .A(n728), .B(KEYINPUT38), .ZN(n736) );
  NAND2_X1 U807 ( .A1(n903), .A2(G129), .ZN(n729) );
  XNOR2_X1 U808 ( .A(n729), .B(KEYINPUT86), .ZN(n731) );
  NAND2_X1 U809 ( .A1(G117), .A2(n904), .ZN(n730) );
  NAND2_X1 U810 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U811 ( .A1(G141), .A2(n899), .ZN(n732) );
  XNOR2_X1 U812 ( .A(KEYINPUT87), .B(n732), .ZN(n733) );
  NOR2_X1 U813 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U814 ( .A1(n736), .A2(n735), .ZN(n894) );
  AND2_X1 U815 ( .A1(G1996), .A2(n894), .ZN(n737) );
  NOR2_X1 U816 ( .A1(n738), .A2(n737), .ZN(n934) );
  NOR2_X1 U817 ( .A1(n934), .A2(n739), .ZN(n748) );
  XOR2_X1 U818 ( .A(n748), .B(KEYINPUT88), .Z(n741) );
  XNOR2_X1 U819 ( .A(G1986), .B(G290), .ZN(n1019) );
  NAND2_X1 U820 ( .A1(n1019), .A2(n755), .ZN(n740) );
  AND2_X1 U821 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U822 ( .A(n745), .B(n744), .ZN(n758) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n894), .ZN(n927) );
  AND2_X1 U824 ( .A1(n952), .A2(n910), .ZN(n932) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n746) );
  NOR2_X1 U826 ( .A1(n932), .A2(n746), .ZN(n747) );
  NOR2_X1 U827 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U828 ( .A1(n927), .A2(n749), .ZN(n750) );
  XNOR2_X1 U829 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U830 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U831 ( .A1(n913), .A2(n753), .ZN(n925) );
  NAND2_X1 U832 ( .A1(n754), .A2(n925), .ZN(n756) );
  NAND2_X1 U833 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U834 ( .A1(n758), .A2(n757), .ZN(n761) );
  XOR2_X1 U835 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n759) );
  XNOR2_X1 U836 ( .A(n761), .B(n760), .ZN(G329) );
  AND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n764) );
  AND2_X1 U838 ( .A1(n764), .A2(n512), .ZN(G160) );
  XOR2_X1 U839 ( .A(KEYINPUT105), .B(G2435), .Z(n766) );
  XNOR2_X1 U840 ( .A(G2430), .B(G2438), .ZN(n765) );
  XNOR2_X1 U841 ( .A(n766), .B(n765), .ZN(n773) );
  XOR2_X1 U842 ( .A(G2446), .B(G2454), .Z(n768) );
  XNOR2_X1 U843 ( .A(G2451), .B(G2443), .ZN(n767) );
  XNOR2_X1 U844 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U845 ( .A(n769), .B(G2427), .Z(n771) );
  XNOR2_X1 U846 ( .A(G1341), .B(G1348), .ZN(n770) );
  XNOR2_X1 U847 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U848 ( .A(n773), .B(n772), .ZN(n774) );
  AND2_X1 U849 ( .A1(n774), .A2(G14), .ZN(G401) );
  AND2_X1 U850 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U851 ( .A1(G123), .A2(n903), .ZN(n775) );
  XNOR2_X1 U852 ( .A(n775), .B(KEYINPUT74), .ZN(n776) );
  XNOR2_X1 U853 ( .A(n776), .B(KEYINPUT18), .ZN(n778) );
  NAND2_X1 U854 ( .A1(G111), .A2(n904), .ZN(n777) );
  NAND2_X1 U855 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U856 ( .A1(G99), .A2(n898), .ZN(n780) );
  NAND2_X1 U857 ( .A1(G135), .A2(n899), .ZN(n779) );
  NAND2_X1 U858 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U859 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U860 ( .A(KEYINPUT75), .B(n783), .ZN(n929) );
  XNOR2_X1 U861 ( .A(G2096), .B(n929), .ZN(n784) );
  OR2_X1 U862 ( .A1(G2100), .A2(n784), .ZN(G156) );
  INV_X1 U863 ( .A(G132), .ZN(G219) );
  INV_X1 U864 ( .A(G82), .ZN(G220) );
  INV_X1 U865 ( .A(G120), .ZN(G236) );
  NAND2_X1 U866 ( .A1(G7), .A2(G661), .ZN(n785) );
  XNOR2_X1 U867 ( .A(n785), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U868 ( .A(G223), .ZN(n842) );
  NAND2_X1 U869 ( .A1(n842), .A2(G567), .ZN(n786) );
  XOR2_X1 U870 ( .A(KEYINPUT11), .B(n786), .Z(G234) );
  INV_X1 U871 ( .A(G860), .ZN(n791) );
  OR2_X1 U872 ( .A1(n1007), .A2(n791), .ZN(G153) );
  INV_X1 U873 ( .A(G171), .ZN(G301) );
  NAND2_X1 U874 ( .A1(G301), .A2(G868), .ZN(n788) );
  INV_X1 U875 ( .A(n849), .ZN(n1012) );
  INV_X1 U876 ( .A(G868), .ZN(n823) );
  NAND2_X1 U877 ( .A1(n1012), .A2(n823), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(G284) );
  INV_X1 U879 ( .A(n1003), .ZN(G299) );
  NOR2_X1 U880 ( .A1(G868), .A2(G299), .ZN(n790) );
  NOR2_X1 U881 ( .A1(G286), .A2(n823), .ZN(n789) );
  NOR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(G297) );
  NAND2_X1 U883 ( .A1(n791), .A2(G559), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n792), .A2(n849), .ZN(n793) );
  XNOR2_X1 U885 ( .A(n793), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U886 ( .A1(n1012), .A2(n823), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n794), .B(KEYINPUT73), .ZN(n795) );
  NOR2_X1 U888 ( .A1(G559), .A2(n795), .ZN(n797) );
  NOR2_X1 U889 ( .A1(G868), .A2(n1007), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(G282) );
  NAND2_X1 U891 ( .A1(G559), .A2(n849), .ZN(n798) );
  XNOR2_X1 U892 ( .A(n798), .B(KEYINPUT76), .ZN(n820) );
  XNOR2_X1 U893 ( .A(n820), .B(n1007), .ZN(n799) );
  NOR2_X1 U894 ( .A1(n799), .A2(G860), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G55), .A2(n800), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n801), .B(KEYINPUT78), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G80), .A2(n802), .ZN(n803) );
  XOR2_X1 U898 ( .A(KEYINPUT77), .B(n803), .Z(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n811) );
  NAND2_X1 U900 ( .A1(G67), .A2(n806), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G93), .A2(n807), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  OR2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n822) );
  XOR2_X1 U904 ( .A(n812), .B(n822), .Z(G145) );
  XNOR2_X1 U905 ( .A(n822), .B(KEYINPUT80), .ZN(n814) );
  XNOR2_X1 U906 ( .A(G166), .B(KEYINPUT19), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n814), .B(n813), .ZN(n817) );
  XOR2_X1 U908 ( .A(G290), .B(n1007), .Z(n815) );
  XNOR2_X1 U909 ( .A(G288), .B(n815), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n817), .B(n816), .ZN(n819) );
  XNOR2_X1 U911 ( .A(G305), .B(n1003), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n819), .B(n818), .ZN(n850) );
  XNOR2_X1 U913 ( .A(n820), .B(n850), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(G868), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U917 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT20), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n827), .B(KEYINPUT81), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n828), .A2(G2090), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U923 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U924 ( .A1(G69), .A2(G57), .ZN(n831) );
  NOR2_X1 U925 ( .A1(G236), .A2(n831), .ZN(n832) );
  XNOR2_X1 U926 ( .A(KEYINPUT82), .B(n832), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(G108), .ZN(n847) );
  NAND2_X1 U928 ( .A1(n847), .A2(G567), .ZN(n838) );
  NOR2_X1 U929 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U930 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U931 ( .A1(G218), .A2(n835), .ZN(n836) );
  NAND2_X1 U932 ( .A1(G96), .A2(n836), .ZN(n848) );
  NAND2_X1 U933 ( .A1(n848), .A2(G2106), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n922) );
  NAND2_X1 U935 ( .A1(G661), .A2(G483), .ZN(n839) );
  XOR2_X1 U936 ( .A(KEYINPUT83), .B(n839), .Z(n840) );
  NOR2_X1 U937 ( .A1(n922), .A2(n840), .ZN(n841) );
  XNOR2_X1 U938 ( .A(KEYINPUT84), .B(n841), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G36), .A2(n845), .ZN(G176) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U942 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U944 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT106), .B(n846), .ZN(G188) );
  XNOR2_X1 U946 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  XOR2_X1 U947 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NOR2_X1 U948 ( .A1(n848), .A2(n847), .ZN(G325) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  XNOR2_X1 U950 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U952 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U953 ( .A(G286), .B(n849), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(G171), .B(n852), .Z(n853) );
  NOR2_X1 U956 ( .A1(G37), .A2(n853), .ZN(n854) );
  XOR2_X1 U957 ( .A(KEYINPUT115), .B(n854), .Z(G397) );
  XOR2_X1 U958 ( .A(G2096), .B(KEYINPUT43), .Z(n856) );
  XNOR2_X1 U959 ( .A(G2067), .B(KEYINPUT110), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U961 ( .A(n857), .B(G2678), .Z(n859) );
  XNOR2_X1 U962 ( .A(G2090), .B(G2072), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U964 ( .A(KEYINPUT42), .B(G2100), .Z(n861) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(G227) );
  XOR2_X1 U968 ( .A(G1976), .B(G1961), .Z(n865) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1971), .ZN(n864) );
  XNOR2_X1 U970 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U971 ( .A(n866), .B(KEYINPUT41), .Z(n868) );
  XNOR2_X1 U972 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U973 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U974 ( .A(G2474), .B(G1966), .Z(n870) );
  XNOR2_X1 U975 ( .A(G1981), .B(G1956), .ZN(n869) );
  XNOR2_X1 U976 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n872), .B(n871), .ZN(G229) );
  NAND2_X1 U978 ( .A1(n903), .A2(G124), .ZN(n873) );
  XNOR2_X1 U979 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G112), .A2(n904), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G100), .A2(n898), .ZN(n877) );
  NAND2_X1 U983 ( .A1(G136), .A2(n899), .ZN(n876) );
  NAND2_X1 U984 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U985 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G130), .A2(n903), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n904), .A2(G118), .ZN(n880) );
  XNOR2_X1 U988 ( .A(KEYINPUT111), .B(n880), .ZN(n886) );
  NAND2_X1 U989 ( .A1(G106), .A2(n898), .ZN(n882) );
  NAND2_X1 U990 ( .A1(G142), .A2(n899), .ZN(n881) );
  NAND2_X1 U991 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  XNOR2_X1 U993 ( .A(KEYINPUT112), .B(n884), .ZN(n885) );
  NOR2_X1 U994 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U995 ( .A1(n888), .A2(n887), .ZN(n892) );
  XOR2_X1 U996 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n890) );
  XNOR2_X1 U997 ( .A(G164), .B(KEYINPUT114), .ZN(n889) );
  XNOR2_X1 U998 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U999 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U1000 ( .A(n929), .B(n893), .ZN(n896) );
  XOR2_X1 U1001 ( .A(G160), .B(n894), .Z(n895) );
  XNOR2_X1 U1002 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U1003 ( .A(n897), .B(G162), .Z(n912) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n898), .ZN(n901) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n899), .ZN(n900) );
  NAND2_X1 U1006 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1007 ( .A(KEYINPUT113), .B(n902), .Z(n909) );
  NAND2_X1 U1008 ( .A1(G127), .A2(n903), .ZN(n906) );
  NAND2_X1 U1009 ( .A1(G115), .A2(n904), .ZN(n905) );
  NAND2_X1 U1010 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1011 ( .A(KEYINPUT47), .B(n907), .Z(n908) );
  NOR2_X1 U1012 ( .A1(n909), .A2(n908), .ZN(n935) );
  XNOR2_X1 U1013 ( .A(n910), .B(n935), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n915), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n922), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(G397), .A2(n917), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n920), .A2(G395), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(n921), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1024 ( .A(G308), .ZN(G225) );
  INV_X1 U1025 ( .A(n922), .ZN(G319) );
  INV_X1 U1026 ( .A(n923), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n945) );
  XNOR2_X1 U1028 ( .A(G160), .B(G2084), .ZN(n943) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n928), .Z(n930) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n941) );
  XOR2_X1 U1035 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT118), .B(n938), .Z(n939) );
  XNOR2_X1 U1039 ( .A(KEYINPUT50), .B(n939), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1043 ( .A(KEYINPUT52), .B(n946), .Z(n947) );
  NOR2_X1 U1044 ( .A1(KEYINPUT55), .A2(n947), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT119), .B(n948), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(G29), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(n950), .ZN(n1001) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(G2090), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(n951), .B(G35), .ZN(n967) );
  XNOR2_X1 U1050 ( .A(G25), .B(n952), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n953), .A2(G28), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(G1996), .B(G32), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n954), .B(G27), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(KEYINPUT122), .B(n957), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G2067), .B(G26), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(n965), .B(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G34), .B(G2084), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1067 ( .A(KEYINPUT55), .B(n971), .Z(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT124), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(G29), .A2(n973), .ZN(n999) );
  XOR2_X1 U1070 ( .A(G16), .B(KEYINPUT126), .Z(n996) );
  XNOR2_X1 U1071 ( .A(G1961), .B(G5), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G21), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n986) );
  XOR2_X1 U1074 ( .A(G1981), .B(G6), .Z(n977) );
  XNOR2_X1 U1075 ( .A(n1002), .B(G20), .ZN(n976) );
  NAND2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n983) );
  XOR2_X1 U1077 ( .A(G1341), .B(G19), .Z(n981) );
  XOR2_X1 U1078 ( .A(KEYINPUT59), .B(G4), .Z(n978) );
  XNOR2_X1 U1079 ( .A(KEYINPUT127), .B(n978), .ZN(n979) );
  XNOR2_X1 U1080 ( .A(n979), .B(G1348), .ZN(n980) );
  NAND2_X1 U1081 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1082 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1083 ( .A(n984), .B(KEYINPUT60), .ZN(n985) );
  NAND2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1086 ( .A(G23), .B(G1976), .ZN(n987) );
  NOR2_X1 U1087 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1088 ( .A(G1986), .B(G24), .Z(n989) );
  NAND2_X1 U1089 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1090 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1092 ( .A(n994), .B(KEYINPUT61), .ZN(n995) );
  NAND2_X1 U1093 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1094 ( .A1(G11), .A2(n997), .ZN(n998) );
  NOR2_X1 U1095 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1096 ( .A1(n1001), .A2(n1000), .ZN(n1030) );
  XOR2_X1 U1097 ( .A(KEYINPUT56), .B(G16), .Z(n1028) );
  XNOR2_X1 U1098 ( .A(G1961), .B(G171), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(KEYINPUT125), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1100 ( .A(n1004), .B(n1003), .ZN(n1006) );
  NAND2_X1 U1101 ( .A1(G1971), .A2(G303), .ZN(n1005) );
  NAND2_X1 U1102 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1103 ( .A(G1341), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1104 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1105 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1106 ( .A(G1348), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1026) );
  INV_X1 U1109 ( .A(n1017), .ZN(n1018) );
  NOR2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(G168), .B(G1966), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT57), .ZN(n1023) );
  NAND2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1118 ( .A(n1031), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

