

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U326 ( .A(n355), .B(n354), .ZN(n357) );
  XOR2_X1 U327 ( .A(KEYINPUT36), .B(n567), .Z(n584) );
  NOR2_X1 U328 ( .A1(n539), .A2(n454), .ZN(n566) );
  XNOR2_X1 U329 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G204GAT), .B(KEYINPUT72), .Z(n294) );
  XNOR2_X1 U332 ( .A(G92GAT), .B(G64GAT), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n417) );
  XNOR2_X1 U334 ( .A(G148GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n295), .B(G78GAT), .ZN(n337) );
  XOR2_X1 U336 ( .A(n417), .B(n337), .Z(n300) );
  XOR2_X1 U337 ( .A(G120GAT), .B(G176GAT), .Z(n297) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G71GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n317) );
  XNOR2_X1 U340 ( .A(G85GAT), .B(KEYINPUT70), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n298), .B(KEYINPUT71), .ZN(n356) );
  XNOR2_X1 U342 ( .A(n317), .B(n356), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n307) );
  XOR2_X1 U344 ( .A(G57GAT), .B(KEYINPUT13), .Z(n368) );
  XOR2_X1 U345 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n302) );
  XNOR2_X1 U346 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U348 ( .A(n368), .B(n303), .Z(n305) );
  NAND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U351 ( .A(n307), .B(n306), .Z(n577) );
  XNOR2_X1 U352 ( .A(n577), .B(KEYINPUT41), .ZN(n555) );
  XNOR2_X1 U353 ( .A(KEYINPUT108), .B(n555), .ZN(n541) );
  XOR2_X1 U354 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n309) );
  XNOR2_X1 U355 ( .A(G190GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U357 ( .A(n310), .B(KEYINPUT17), .Z(n312) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(KEYINPUT86), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n425) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n313), .B(KEYINPUT83), .ZN(n437) );
  XOR2_X1 U362 ( .A(G43GAT), .B(G134GAT), .Z(n352) );
  XOR2_X1 U363 ( .A(n437), .B(n352), .Z(n315) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(n316), .B(KEYINPUT84), .Z(n319) );
  XNOR2_X1 U367 ( .A(n317), .B(KEYINPUT20), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n320), .B(KEYINPUT85), .Z(n322) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G127GAT), .Z(n370) );
  XNOR2_X1 U371 ( .A(n370), .B(KEYINPUT87), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n425), .B(n323), .ZN(n525) );
  INV_X1 U374 ( .A(n525), .ZN(n539) );
  XOR2_X1 U375 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n325) );
  XNOR2_X1 U376 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(KEYINPUT95), .B(n326), .Z(n328) );
  NAND2_X1 U379 ( .A1(G228GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U381 ( .A(n329), .B(KEYINPUT89), .Z(n335) );
  XNOR2_X1 U382 ( .A(G218GAT), .B(G211GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n330), .B(KEYINPUT21), .ZN(n331) );
  XOR2_X1 U384 ( .A(n331), .B(KEYINPUT92), .Z(n333) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(KEYINPUT91), .ZN(n332) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n426) );
  XOR2_X1 U387 ( .A(G204GAT), .B(n426), .Z(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G155GAT), .Z(n369) );
  XOR2_X1 U390 ( .A(n336), .B(n369), .Z(n339) );
  XOR2_X1 U391 ( .A(G50GAT), .B(G162GAT), .Z(n350) );
  XNOR2_X1 U392 ( .A(n337), .B(n350), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U394 ( .A(KEYINPUT93), .B(KEYINPUT2), .Z(n341) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT94), .B(n342), .Z(n436) );
  XOR2_X1 U398 ( .A(n343), .B(n436), .Z(n469) );
  XOR2_X1 U399 ( .A(G36GAT), .B(KEYINPUT78), .Z(n420) );
  XOR2_X1 U400 ( .A(G29GAT), .B(KEYINPUT8), .Z(n345) );
  XNOR2_X1 U401 ( .A(KEYINPUT7), .B(KEYINPUT68), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n392) );
  XOR2_X1 U403 ( .A(n420), .B(n392), .Z(n347) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT79), .B(KEYINPUT74), .Z(n349) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U409 ( .A(n351), .B(n350), .Z(n353) );
  XOR2_X1 U410 ( .A(n357), .B(n356), .Z(n359) );
  XNOR2_X1 U411 ( .A(G190GAT), .B(KEYINPUT77), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n367) );
  XOR2_X1 U413 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n361) );
  XNOR2_X1 U414 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U416 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n363) );
  XNOR2_X1 U417 ( .A(G99GAT), .B(KEYINPUT76), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U419 ( .A(n365), .B(n364), .Z(n366) );
  XOR2_X2 U420 ( .A(n367), .B(n366), .Z(n567) );
  INV_X1 U421 ( .A(n567), .ZN(n408) );
  XOR2_X1 U422 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U423 ( .A(G8GAT), .B(G1GAT), .Z(n389) );
  XNOR2_X1 U424 ( .A(n389), .B(n370), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n385) );
  XOR2_X1 U426 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n374) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U429 ( .A(n375), .B(KEYINPUT82), .Z(n383) );
  XOR2_X1 U430 ( .A(G211GAT), .B(KEYINPUT15), .Z(n377) );
  XNOR2_X1 U431 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U433 ( .A(G64GAT), .B(G78GAT), .Z(n379) );
  XNOR2_X1 U434 ( .A(G183GAT), .B(G71GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n487) );
  INV_X1 U439 ( .A(n487), .ZN(n580) );
  XOR2_X1 U440 ( .A(KEYINPUT69), .B(G22GAT), .Z(n387) );
  XNOR2_X1 U441 ( .A(G50GAT), .B(G15GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U443 ( .A(n388), .B(G43GAT), .Z(n391) );
  XNOR2_X1 U444 ( .A(n389), .B(G36GAT), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n396) );
  XOR2_X1 U446 ( .A(G169GAT), .B(n392), .Z(n394) );
  NAND2_X1 U447 ( .A1(G229GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U449 ( .A(n396), .B(n395), .Z(n404) );
  XOR2_X1 U450 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n398) );
  XNOR2_X1 U451 ( .A(KEYINPUT65), .B(KEYINPUT30), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U453 ( .A(G197GAT), .B(G141GAT), .Z(n400) );
  XNOR2_X1 U454 ( .A(KEYINPUT29), .B(G113GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U457 ( .A(n404), .B(n403), .Z(n504) );
  INV_X1 U458 ( .A(n504), .ZN(n573) );
  NAND2_X1 U459 ( .A1(n573), .A2(n555), .ZN(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT46), .B(n405), .Z(n406) );
  NOR2_X1 U461 ( .A1(n580), .A2(n406), .ZN(n407) );
  NAND2_X1 U462 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n409), .B(KEYINPUT47), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n410), .B(KEYINPUT118), .ZN(n415) );
  NOR2_X1 U465 ( .A1(n584), .A2(n487), .ZN(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT45), .B(n411), .ZN(n412) );
  NAND2_X1 U467 ( .A1(n412), .A2(n577), .ZN(n413) );
  NOR2_X1 U468 ( .A1(n413), .A2(n573), .ZN(n414) );
  NOR2_X1 U469 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(KEYINPUT48), .B(n416), .ZN(n535) );
  XOR2_X1 U471 ( .A(n417), .B(KEYINPUT98), .Z(n419) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U474 ( .A(n421), .B(n420), .Z(n423) );
  XNOR2_X1 U475 ( .A(G8GAT), .B(G176GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n428) );
  INV_X1 U478 ( .A(n426), .ZN(n427) );
  XOR2_X1 U479 ( .A(n428), .B(n427), .Z(n495) );
  NOR2_X1 U480 ( .A1(n535), .A2(n495), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT54), .ZN(n452) );
  XOR2_X1 U482 ( .A(KEYINPUT4), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U483 ( .A(G120GAT), .B(G155GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U485 ( .A(KEYINPUT6), .B(KEYINPUT97), .Z(n433) );
  XNOR2_X1 U486 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n443) );
  INV_X1 U489 ( .A(n436), .ZN(n441) );
  XOR2_X1 U490 ( .A(n437), .B(KEYINPUT1), .Z(n439) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U493 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n451) );
  XOR2_X1 U495 ( .A(G57GAT), .B(KEYINPUT77), .Z(n445) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(G127GAT), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U498 ( .A(G162GAT), .B(G85GAT), .Z(n447) );
  XNOR2_X1 U499 ( .A(G29GAT), .B(G134GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U501 ( .A(n449), .B(n448), .Z(n450) );
  XOR2_X1 U502 ( .A(n451), .B(n450), .Z(n520) );
  INV_X1 U503 ( .A(n520), .ZN(n492) );
  NAND2_X1 U504 ( .A1(n452), .A2(n492), .ZN(n572) );
  NOR2_X1 U505 ( .A1(n469), .A2(n572), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  NAND2_X1 U507 ( .A1(n541), .A2(n566), .ZN(n458) );
  XOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT56), .Z(n456) );
  XNOR2_X1 U509 ( .A(KEYINPUT57), .B(KEYINPUT126), .ZN(n455) );
  XNOR2_X1 U510 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n477) );
  NAND2_X1 U511 ( .A1(n573), .A2(n577), .ZN(n490) );
  NOR2_X1 U512 ( .A1(n567), .A2(n487), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT16), .ZN(n475) );
  XOR2_X1 U514 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n462) );
  NOR2_X1 U515 ( .A1(n539), .A2(n495), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n469), .A2(n460), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U518 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n464) );
  NAND2_X1 U519 ( .A1(n469), .A2(n539), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n570) );
  INV_X1 U521 ( .A(n495), .ZN(n522) );
  XNOR2_X1 U522 ( .A(KEYINPUT27), .B(n522), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n570), .A2(n468), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n492), .A2(n467), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n520), .A2(n468), .ZN(n534) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT28), .ZN(n530) );
  NOR2_X1 U528 ( .A1(n534), .A2(n530), .ZN(n470) );
  XOR2_X1 U529 ( .A(KEYINPUT99), .B(n470), .Z(n472) );
  XOR2_X1 U530 ( .A(n525), .B(KEYINPUT88), .Z(n471) );
  NAND2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n475), .A2(n486), .ZN(n505) );
  NOR2_X1 U534 ( .A1(n490), .A2(n505), .ZN(n483) );
  NAND2_X1 U535 ( .A1(n520), .A2(n483), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n483), .A2(n522), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U541 ( .A1(n483), .A2(n525), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U543 ( .A(G15GAT), .B(n482), .Z(G1326GAT) );
  NAND2_X1 U544 ( .A1(n530), .A2(n483), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(KEYINPUT104), .ZN(n485) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n488), .A2(n584), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT37), .ZN(n518) );
  NOR2_X1 U550 ( .A1(n518), .A2(n490), .ZN(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n491), .Z(n501) );
  NOR2_X1 U552 ( .A1(n501), .A2(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n501), .A2(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n539), .A2(n501), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U561 ( .A(G43GAT), .B(n500), .Z(G1330GAT) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n503) );
  INV_X1 U563 ( .A(n530), .ZN(n537) );
  NOR2_X1 U564 ( .A1(n537), .A2(n501), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n508) );
  NAND2_X1 U567 ( .A1(n541), .A2(n504), .ZN(n517) );
  NOR2_X1 U568 ( .A1(n517), .A2(n505), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT109), .B(n506), .Z(n513) );
  NAND2_X1 U570 ( .A1(n513), .A2(n520), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n509), .Z(G1332GAT) );
  NAND2_X1 U573 ( .A1(n513), .A2(n522), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT111), .Z(n512) );
  NAND2_X1 U576 ( .A1(n513), .A2(n525), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n530), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT113), .B(n519), .Z(n531) );
  NAND2_X1 U584 ( .A1(n531), .A2(n520), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G85GAT), .ZN(G1336GAT) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT114), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n531), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT117), .B(KEYINPUT44), .Z(n528) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(n529), .Z(n533) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT119), .B(n536), .Z(n552) );
  NAND2_X1 U599 ( .A1(n552), .A2(n537), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n547), .A2(n573), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U604 ( .A1(n547), .A2(n541), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n545) );
  NAND2_X1 U607 ( .A1(n547), .A2(n580), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U609 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U611 ( .A1(n547), .A2(n567), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT121), .Z(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n570), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n553), .B(KEYINPUT123), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n561), .A2(n573), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT124), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U621 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n580), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n567), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n573), .A2(n566), .ZN(n564) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT125), .Z(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n580), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  INV_X1 U637 ( .A(n570), .ZN(n571) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U643 ( .A(n581), .ZN(n583) );
  OR2_X1 U644 ( .A1(n583), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

