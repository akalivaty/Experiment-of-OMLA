

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U320 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U321 ( .A(n421), .B(n420), .ZN(n425) );
  NOR2_X1 U322 ( .A1(n540), .A2(n522), .ZN(n526) );
  XNOR2_X1 U323 ( .A(n358), .B(n357), .ZN(n362) );
  XNOR2_X1 U324 ( .A(KEYINPUT97), .B(n405), .ZN(n516) );
  NOR2_X1 U325 ( .A1(n487), .A2(n503), .ZN(n495) );
  XOR2_X1 U326 ( .A(KEYINPUT95), .B(n342), .Z(n288) );
  XNOR2_X1 U327 ( .A(n463), .B(KEYINPUT47), .ZN(n464) );
  INV_X1 U328 ( .A(n436), .ZN(n355) );
  INV_X1 U329 ( .A(KEYINPUT64), .ZN(n468) );
  XNOR2_X1 U330 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U331 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U332 ( .A(n468), .B(KEYINPUT48), .ZN(n469) );
  NOR2_X1 U333 ( .A1(n581), .A2(n409), .ZN(n411) );
  XNOR2_X1 U334 ( .A(n470), .B(n469), .ZN(n541) );
  XOR2_X1 U335 ( .A(n395), .B(n394), .Z(n492) );
  NOR2_X1 U336 ( .A1(n492), .A2(n477), .ZN(n560) );
  XNOR2_X1 U337 ( .A(n451), .B(n450), .ZN(n500) );
  XNOR2_X1 U338 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U339 ( .A(n452), .B(G29GAT), .ZN(n453) );
  XNOR2_X1 U340 ( .A(n482), .B(n481), .ZN(G1349GAT) );
  XNOR2_X1 U341 ( .A(n454), .B(n453), .ZN(G1328GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT76), .B(KEYINPUT66), .Z(n290) );
  XNOR2_X1 U343 ( .A(G92GAT), .B(KEYINPUT77), .ZN(n289) );
  XNOR2_X1 U344 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .Z(n440) );
  XOR2_X1 U346 ( .A(n291), .B(n440), .Z(n293) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(G106GAT), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n298) );
  XOR2_X1 U349 ( .A(G29GAT), .B(G134GAT), .Z(n353) );
  XNOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n294), .B(KEYINPUT78), .ZN(n327) );
  XOR2_X1 U352 ( .A(n353), .B(n327), .Z(n296) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n306) );
  XOR2_X1 U356 ( .A(KEYINPUT7), .B(KEYINPUT70), .Z(n300) );
  XNOR2_X1 U357 ( .A(G50GAT), .B(G43GAT), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U359 ( .A(KEYINPUT8), .B(n301), .Z(n423) );
  XOR2_X1 U360 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n303) );
  XNOR2_X1 U361 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n423), .B(n304), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n553) );
  XNOR2_X1 U365 ( .A(n553), .B(KEYINPUT36), .ZN(n581) );
  XOR2_X1 U366 ( .A(G64GAT), .B(G57GAT), .Z(n308) );
  XNOR2_X1 U367 ( .A(G211GAT), .B(G78GAT), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U369 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n310) );
  XNOR2_X1 U370 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U372 ( .A(n312), .B(n311), .Z(n322) );
  XOR2_X1 U373 ( .A(G71GAT), .B(KEYINPUT13), .Z(n441) );
  XOR2_X1 U374 ( .A(G1GAT), .B(G127GAT), .Z(n352) );
  XOR2_X1 U375 ( .A(n441), .B(n352), .Z(n314) );
  XNOR2_X1 U376 ( .A(G183GAT), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U377 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U378 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n316) );
  NAND2_X1 U379 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U380 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n320) );
  XOR2_X1 U382 ( .A(G15GAT), .B(G22GAT), .Z(n422) );
  XOR2_X1 U383 ( .A(n422), .B(KEYINPUT15), .Z(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n578) );
  INV_X1 U386 ( .A(n578), .ZN(n550) );
  XNOR2_X1 U387 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n323), .B(G183GAT), .ZN(n324) );
  XOR2_X1 U389 ( .A(n324), .B(KEYINPUT17), .Z(n326) );
  XNOR2_X1 U390 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n391) );
  XOR2_X1 U392 ( .A(KEYINPUT98), .B(n327), .Z(n329) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U395 ( .A(KEYINPUT73), .B(G64GAT), .Z(n331) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G92GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U398 ( .A(G204GAT), .B(n332), .Z(n446) );
  XOR2_X1 U399 ( .A(n333), .B(n446), .Z(n338) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n417) );
  XOR2_X1 U401 ( .A(KEYINPUT91), .B(G218GAT), .Z(n335) );
  XNOR2_X1 U402 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U404 ( .A(G197GAT), .B(n336), .Z(n374) );
  XNOR2_X1 U405 ( .A(n417), .B(n374), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U407 ( .A(n391), .B(n339), .Z(n518) );
  XOR2_X1 U408 ( .A(KEYINPUT27), .B(n518), .Z(n401) );
  INV_X1 U409 ( .A(n401), .ZN(n363) );
  XOR2_X1 U410 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n341) );
  XNOR2_X1 U411 ( .A(KEYINPUT5), .B(KEYINPUT96), .ZN(n340) );
  XNOR2_X1 U412 ( .A(n341), .B(n340), .ZN(n342) );
  NAND2_X1 U413 ( .A1(G225GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n288), .B(n343), .ZN(n344) );
  XOR2_X1 U415 ( .A(n344), .B(KEYINPUT4), .Z(n351) );
  XOR2_X1 U416 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n346) );
  XNOR2_X1 U417 ( .A(G162GAT), .B(KEYINPUT93), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U419 ( .A(n347), .B(KEYINPUT3), .Z(n349) );
  XNOR2_X1 U420 ( .A(G141GAT), .B(G155GAT), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n378), .B(G85GAT), .ZN(n350) );
  XNOR2_X1 U423 ( .A(n351), .B(n350), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n356) );
  XNOR2_X1 U425 ( .A(G120GAT), .B(G148GAT), .ZN(n354) );
  XNOR2_X1 U426 ( .A(n354), .B(G57GAT), .ZN(n436) );
  XOR2_X1 U427 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n360) );
  XNOR2_X1 U428 ( .A(KEYINPUT0), .B(KEYINPUT83), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U430 ( .A(G113GAT), .B(n361), .ZN(n395) );
  XNOR2_X1 U431 ( .A(n362), .B(n395), .ZN(n405) );
  NAND2_X1 U432 ( .A1(n363), .A2(n516), .ZN(n364) );
  XOR2_X1 U433 ( .A(KEYINPUT99), .B(n364), .Z(n540) );
  XOR2_X1 U434 ( .A(KEYINPUT22), .B(G148GAT), .Z(n366) );
  XNOR2_X1 U435 ( .A(KEYINPUT90), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U437 ( .A(G106GAT), .B(G78GAT), .Z(n447) );
  XOR2_X1 U438 ( .A(n367), .B(n447), .Z(n369) );
  XNOR2_X1 U439 ( .A(G50GAT), .B(G22GAT), .ZN(n368) );
  XNOR2_X1 U440 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U441 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n371) );
  NAND2_X1 U442 ( .A1(G228GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U444 ( .A(n373), .B(n372), .Z(n376) );
  XNOR2_X1 U445 ( .A(n374), .B(KEYINPUT23), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U447 ( .A(n378), .B(n377), .Z(n475) );
  XNOR2_X1 U448 ( .A(n475), .B(KEYINPUT28), .ZN(n522) );
  XOR2_X1 U449 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n380) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(G127GAT), .ZN(n379) );
  XNOR2_X1 U451 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U452 ( .A(G120GAT), .B(G176GAT), .Z(n382) );
  XNOR2_X1 U453 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n381) );
  XNOR2_X1 U454 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U455 ( .A(n384), .B(n383), .Z(n393) );
  XOR2_X1 U456 ( .A(G190GAT), .B(G99GAT), .Z(n386) );
  XNOR2_X1 U457 ( .A(G43GAT), .B(G134GAT), .ZN(n385) );
  XNOR2_X1 U458 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U459 ( .A(G71GAT), .B(n387), .Z(n389) );
  NAND2_X1 U460 ( .A1(G227GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U461 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U462 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U464 ( .A1(n526), .A2(n492), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n396), .B(KEYINPUT100), .ZN(n408) );
  INV_X1 U466 ( .A(n518), .ZN(n471) );
  NOR2_X1 U467 ( .A1(n492), .A2(n471), .ZN(n397) );
  NOR2_X1 U468 ( .A1(n475), .A2(n397), .ZN(n398) );
  XOR2_X1 U469 ( .A(KEYINPUT25), .B(n398), .Z(n403) );
  XOR2_X1 U470 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n400) );
  NAND2_X1 U471 ( .A1(n475), .A2(n492), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n400), .B(n399), .ZN(n566) );
  NOR2_X1 U473 ( .A1(n566), .A2(n401), .ZN(n402) );
  NOR2_X1 U474 ( .A1(n403), .A2(n402), .ZN(n404) );
  XOR2_X1 U475 ( .A(KEYINPUT102), .B(n404), .Z(n406) );
  NAND2_X1 U476 ( .A1(n406), .A2(n405), .ZN(n407) );
  NAND2_X1 U477 ( .A1(n408), .A2(n407), .ZN(n485) );
  NAND2_X1 U478 ( .A1(n550), .A2(n485), .ZN(n409) );
  XOR2_X1 U479 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n515) );
  XOR2_X1 U481 ( .A(G1GAT), .B(G197GAT), .Z(n413) );
  XNOR2_X1 U482 ( .A(G113GAT), .B(G141GAT), .ZN(n412) );
  XOR2_X1 U483 ( .A(n413), .B(n412), .Z(n414) );
  XNOR2_X1 U484 ( .A(n414), .B(G36GAT), .ZN(n421) );
  XOR2_X1 U485 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n416) );
  NAND2_X1 U486 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XOR2_X1 U487 ( .A(n416), .B(n415), .Z(n419) );
  XNOR2_X1 U488 ( .A(n417), .B(G29GAT), .ZN(n418) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U491 ( .A(KEYINPUT68), .B(KEYINPUT71), .Z(n427) );
  XNOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n543) );
  INV_X1 U495 ( .A(n543), .ZN(n568) );
  INV_X1 U496 ( .A(KEYINPUT32), .ZN(n430) );
  NAND2_X1 U497 ( .A1(KEYINPUT75), .A2(n430), .ZN(n433) );
  INV_X1 U498 ( .A(KEYINPUT75), .ZN(n431) );
  NAND2_X1 U499 ( .A1(n431), .A2(KEYINPUT32), .ZN(n432) );
  NAND2_X1 U500 ( .A1(n433), .A2(n432), .ZN(n435) );
  XNOR2_X1 U501 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U504 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n438) );
  XNOR2_X1 U505 ( .A(n439), .B(n438), .ZN(n445) );
  XOR2_X1 U506 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n442) );
  XOR2_X1 U508 ( .A(n443), .B(n442), .Z(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n459) );
  NAND2_X1 U512 ( .A1(n568), .A2(n459), .ZN(n487) );
  NOR2_X1 U513 ( .A1(n515), .A2(n487), .ZN(n451) );
  XNOR2_X1 U514 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n450) );
  NAND2_X1 U515 ( .A1(n500), .A2(n516), .ZN(n454) );
  XOR2_X1 U516 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n452) );
  NOR2_X1 U517 ( .A1(n550), .A2(n581), .ZN(n455) );
  XNOR2_X1 U518 ( .A(KEYINPUT45), .B(n455), .ZN(n456) );
  NAND2_X1 U519 ( .A1(n456), .A2(n459), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n568), .A2(n457), .ZN(n458) );
  XOR2_X1 U521 ( .A(KEYINPUT113), .B(n458), .Z(n467) );
  XOR2_X1 U522 ( .A(n459), .B(KEYINPUT41), .Z(n545) );
  INV_X1 U523 ( .A(n545), .ZN(n478) );
  NAND2_X1 U524 ( .A1(n568), .A2(n478), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n460), .B(KEYINPUT46), .ZN(n462) );
  INV_X1 U526 ( .A(n553), .ZN(n559) );
  AND2_X1 U527 ( .A1(n550), .A2(n553), .ZN(n461) );
  AND2_X1 U528 ( .A1(n462), .A2(n461), .ZN(n465) );
  XNOR2_X1 U529 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n463) );
  NOR2_X1 U530 ( .A1(n467), .A2(n466), .ZN(n470) );
  INV_X1 U531 ( .A(n541), .ZN(n525) );
  NOR2_X1 U532 ( .A1(n525), .A2(n471), .ZN(n472) );
  XOR2_X1 U533 ( .A(n472), .B(KEYINPUT54), .Z(n473) );
  NOR2_X1 U534 ( .A1(n516), .A2(n473), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT65), .B(n474), .ZN(n565) );
  NOR2_X1 U536 ( .A1(n475), .A2(n565), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n476), .B(KEYINPUT55), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n560), .A2(n478), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n480) );
  XNOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n479) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(KEYINPUT82), .ZN(n484) );
  NOR2_X1 U543 ( .A1(n559), .A2(n550), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n503) );
  NAND2_X1 U546 ( .A1(n495), .A2(n516), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT103), .Z(n491) );
  NAND2_X1 U549 ( .A1(n495), .A2(n518), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  INV_X1 U552 ( .A(n492), .ZN(n527) );
  NAND2_X1 U553 ( .A1(n495), .A2(n527), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n522), .A2(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U557 ( .A1(n518), .A2(n500), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n500), .A2(n527), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  XOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U563 ( .A1(n500), .A2(n522), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1331GAT) );
  NAND2_X1 U565 ( .A1(n543), .A2(n478), .ZN(n514) );
  NOR2_X1 U566 ( .A1(n503), .A2(n514), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(KEYINPUT108), .ZN(n510) );
  NAND2_X1 U568 ( .A1(n510), .A2(n516), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n510), .A2(n518), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT109), .Z(n509) );
  NAND2_X1 U574 ( .A1(n527), .A2(n510), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U577 ( .A1(n510), .A2(n522), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n527), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n525), .A2(n528), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n536), .A2(n568), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n536), .A2(n478), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n534) );
  NAND2_X1 U599 ( .A1(n536), .A2(n578), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n559), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n566), .A2(n540), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n552) );
  NOR2_X1 U608 ( .A1(n543), .A2(n552), .ZN(n544) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n552), .A2(n545), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n550), .A2(n552), .ZN(n551) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U618 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n568), .A2(n560), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n578), .A2(n560), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT58), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(n562), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n572) );
  XOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT121), .B(n567), .ZN(n580) );
  INV_X1 U634 ( .A(n580), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n577), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n580), .A2(n459), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n574) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

