//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT70), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n463), .A2(new_n465), .A3(new_n470), .A4(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT69), .B(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n475), .B1(new_n474), .B2(new_n478), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n481), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n473), .ZN(new_n483));
  NOR3_X1   g058(.A1(new_n479), .A2(new_n480), .A3(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n472), .A2(new_n473), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n473), .B1(new_n469), .B2(new_n471), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n473), .A2(G138), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n481), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n467), .B1(new_n476), .B2(KEYINPUT3), .ZN(new_n498));
  AND4_X1   g073(.A1(new_n470), .A2(new_n463), .A3(new_n465), .A4(KEYINPUT3), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n500), .B2(KEYINPUT74), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n469), .B2(new_n471), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n497), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(KEYINPUT73), .B(G114), .Z(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(new_n473), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(G126), .B(G2105), .C1(new_n498), .C2(new_n499), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n488), .A2(KEYINPUT72), .A3(G126), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  AND3_X1   g091(.A1(KEYINPUT75), .A2(KEYINPUT6), .A3(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT6), .B1(KEYINPUT75), .B2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(new_n519), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n522), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(G62), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G166));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT77), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  INV_X1    g115(.A(new_n521), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n524), .A2(G89), .ZN(new_n543));
  NAND2_X1  g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n527), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G168));
  NOR2_X1   g121(.A1(new_n519), .A2(new_n527), .ZN(new_n547));
  AOI22_X1  g122(.A1(G90), .A2(new_n547), .B1(new_n521), .B2(G52), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT78), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n531), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n531), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n521), .A2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n547), .A2(G81), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT79), .ZN(G188));
  XNOR2_X1  g140(.A(new_n547), .B(KEYINPUT80), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n541), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n541), .B2(new_n570), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n527), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n571), .A2(new_n572), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n569), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n566), .A2(G87), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n528), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(G49), .B2(new_n521), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n566), .A2(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n527), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(G48), .A2(new_n521), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT82), .ZN(G305));
  NAND2_X1  g165(.A1(new_n547), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n521), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n531), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n566), .A2(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT83), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n527), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n612), .B2(G860), .ZN(G148));
  OAI21_X1  g188(.A(KEYINPUT85), .B1(new_n559), .B2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n612), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  MUX2_X1   g191(.A(KEYINPUT85), .B(new_n614), .S(new_n616), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n477), .A2(new_n481), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n488), .A2(G123), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n625));
  INV_X1    g200(.A(G135), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n625), .C1(new_n626), .C2(new_n485), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT87), .Z(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n639), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(G14), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  AOI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n662), .C2(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(G23), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(G22), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n679), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1971), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n679), .A2(G6), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G305), .B2(G16), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n689), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n486), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n488), .A2(G119), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G25), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  OR2_X1    g284(.A1(G16), .A2(G24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G290), .B2(new_n679), .ZN(new_n711));
  INV_X1    g286(.A(G1986), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(KEYINPUT89), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  NOR4_X1   g289(.A1(new_n708), .A2(new_n709), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n697), .A2(new_n698), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n486), .A2(G141), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n488), .A2(G129), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT26), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n477), .A2(G105), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n722), .A2(new_n723), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT95), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(KEYINPUT95), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n721), .B1(new_n732), .B2(new_n720), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n720), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n488), .A2(G128), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n473), .A2(G116), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  INV_X1    g316(.A(G140), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n739), .B1(new_n740), .B2(new_n741), .C1(new_n485), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT91), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT91), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n738), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2067), .ZN(new_n748));
  NOR2_X1   g323(.A1(G27), .A2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G164), .B2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2078), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n736), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n720), .A2(G33), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  INV_X1    g330(.A(G139), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n485), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT92), .Z(new_n758));
  AOI22_X1  g333(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n473), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n720), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2072), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n559), .B2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  INV_X1    g341(.A(G28), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT30), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(KEYINPUT30), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n766), .B(new_n772), .C1(new_n720), .C2(new_n627), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n720), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n679), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n679), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1961), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(G1961), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n773), .A2(new_n779), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n720), .A2(G35), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT98), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n492), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT29), .B(G2090), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n679), .A2(G21), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G168), .B2(new_n679), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT97), .Z(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n792), .B2(G1966), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n784), .B(new_n793), .C1(G1966), .C2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n679), .A2(G4), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n607), .B2(new_n679), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT90), .B(G1348), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n679), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT99), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n798), .B(new_n803), .C1(G2084), .C2(new_n778), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n763), .A2(new_n794), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n718), .A2(new_n719), .A3(new_n752), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n547), .A2(G93), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n521), .A2(G55), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n531), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n559), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n808), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT38), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n607), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n821), .A2(new_n822), .A3(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n812), .A2(G860), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT101), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  OR2_X1    g401(.A1(new_n823), .A2(new_n826), .ZN(G145));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n828));
  INV_X1    g403(.A(new_n761), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(KEYINPUT102), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n731), .B(new_n743), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G164), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n761), .A2(KEYINPUT103), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n488), .A2(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n473), .A2(G118), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G142), .B2(new_n486), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(new_n620), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n703), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n833), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n833), .B2(new_n835), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(G160), .B(new_n627), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G162), .ZN(new_n847));
  AOI21_X1  g422(.A(G37), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n845), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g425(.A(G305), .B(G290), .ZN(new_n851));
  XNOR2_X1  g426(.A(G288), .B(G303), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(KEYINPUT105), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(KEYINPUT105), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n607), .A2(G299), .A3(KEYINPUT104), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT104), .B1(new_n607), .B2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n607), .A2(G299), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n817), .B(new_n615), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n862), .B2(new_n866), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n858), .B(new_n868), .ZN(new_n869));
  MUX2_X1   g444(.A(new_n812), .B(new_n869), .S(G868), .Z(G295));
  MUX2_X1   g445(.A(new_n812), .B(new_n869), .S(G868), .Z(G331));
  INV_X1    g446(.A(KEYINPUT109), .ZN(new_n872));
  AOI21_X1  g447(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(KEYINPUT107), .B2(G301), .ZN(new_n874));
  OR3_X1    g449(.A1(G301), .A2(G286), .A3(KEYINPUT107), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n817), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT108), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n874), .A2(new_n816), .A3(new_n815), .A4(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(KEYINPUT108), .A3(new_n817), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n872), .B1(new_n865), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n884), .A2(KEYINPUT109), .A3(new_n864), .A4(new_n863), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n877), .B2(KEYINPUT110), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(KEYINPUT110), .B2(new_n877), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n862), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n889), .B2(new_n854), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n883), .A2(new_n885), .A3(new_n853), .A4(new_n888), .ZN(new_n891));
  XNOR2_X1  g466(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n882), .A2(new_n862), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n887), .B2(new_n865), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n895), .B2(new_n854), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(KEYINPUT44), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT111), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n892), .B1(new_n890), .B2(new_n891), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n891), .A3(new_n892), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n900), .B(new_n905), .C1(new_n901), .C2(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n899), .B1(new_n906), .B2(new_n908), .ZN(G397));
  INV_X1    g484(.A(G1384), .ZN(new_n910));
  INV_X1    g485(.A(new_n509), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n510), .A2(new_n511), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT72), .B1(new_n488), .B2(G126), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n497), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n494), .B1(new_n502), .B2(new_n503), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n500), .A2(KEYINPUT74), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n910), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G160), .A2(G40), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT125), .Z(new_n928));
  INV_X1    g503(.A(new_n923), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n743), .B(G2067), .Z(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n732), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n926), .B2(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n732), .A2(new_n924), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n731), .A2(G1996), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n704), .A2(new_n707), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n704), .A2(new_n707), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n923), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n929), .A2(G1986), .A3(G290), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n939), .B1(new_n937), .B2(new_n923), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n743), .A2(G2067), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n929), .B1(new_n950), .B2(KEYINPUT124), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(KEYINPUT124), .B2(new_n950), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n934), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n479), .A2(new_n480), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT121), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  INV_X1    g531(.A(new_n482), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(KEYINPUT120), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n473), .B1(new_n957), .B2(KEYINPUT120), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n954), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n954), .B2(new_n960), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n963));
  NOR4_X1   g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(G2078), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n515), .A2(KEYINPUT45), .A3(new_n910), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n921), .A2(new_n965), .ZN(new_n966));
  NOR4_X1   g541(.A1(new_n479), .A2(new_n480), .A3(new_n956), .A4(new_n483), .ZN(new_n967));
  INV_X1    g542(.A(G2078), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n921), .A2(new_n967), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n964), .A2(new_n966), .B1(new_n969), .B2(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n919), .A2(KEYINPUT112), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n515), .A2(new_n973), .A3(new_n910), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n967), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1961), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(KEYINPUT119), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT119), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  OAI211_X1 g555(.A(G301), .B(new_n970), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT122), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n978), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n977), .A2(KEYINPUT119), .A3(new_n978), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT122), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G301), .A4(new_n970), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n969), .A2(new_n963), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n505), .B2(new_n514), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n973), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT112), .B(G1384), .C1(new_n505), .C2(new_n514), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n920), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n965), .A2(new_n967), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT53), .A4(new_n968), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n983), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n982), .A2(new_n989), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n569), .A2(new_n1003), .A3(new_n576), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n569), .B2(new_n576), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n921), .A2(new_n967), .A3(new_n965), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT56), .B(G2072), .Z(new_n1009));
  OR2_X1    g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT116), .B(G1956), .Z(new_n1011));
  AOI21_X1  g586(.A(new_n972), .B1(new_n971), .B2(new_n974), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n967), .B1(new_n919), .B2(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1007), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT50), .B1(new_n992), .B2(new_n993), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1013), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1006), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n1004), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n606), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n977), .A2(new_n797), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n971), .A2(new_n967), .A3(new_n974), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(G2067), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1015), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT61), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1023), .B2(new_n1015), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1021), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1010), .A2(new_n1014), .A3(new_n1007), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(KEYINPUT61), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1008), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT58), .B(G1341), .Z(new_n1036));
  AOI22_X1  g611(.A1(new_n1035), .A2(new_n924), .B1(new_n1026), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n1037), .B2(new_n558), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1026), .A2(new_n1036), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1008), .A2(G1996), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1039), .B(new_n559), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1031), .A2(new_n1034), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1025), .A2(KEYINPUT60), .A3(new_n1027), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n607), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1025), .A2(new_n1027), .A3(KEYINPUT60), .A4(new_n606), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1046), .A2(new_n1047), .B1(new_n1048), .B2(new_n1028), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1029), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n971), .A2(new_n974), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n995), .B1(new_n1051), .B2(new_n920), .ZN(new_n1052));
  OAI22_X1  g627(.A1(G2084), .A2(new_n977), .B1(new_n1052), .B2(G1966), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G168), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(new_n1057), .C1(KEYINPUT117), .C2(KEYINPUT51), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n1057), .B2(KEYINPUT117), .ZN(new_n1059));
  OAI211_X1 g634(.A(G8), .B(new_n1059), .C1(new_n1053), .C2(G286), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n983), .A2(G301), .A3(new_n990), .A4(new_n997), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT54), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(G171), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G303), .A2(G8), .ZN(new_n1067));
  XOR2_X1   g642(.A(new_n1067), .B(KEYINPUT55), .Z(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1070));
  INV_X1    g645(.A(G2090), .ZN(new_n1071));
  INV_X1    g646(.A(G1971), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1070), .A2(new_n1071), .B1(new_n1072), .B2(new_n1008), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1073), .B2(new_n1055), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n589), .A2(G1981), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT114), .B(G86), .Z(new_n1076));
  OAI21_X1  g651(.A(new_n588), .B1(new_n529), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G1981), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1026), .A3(G8), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n678), .A2(G1976), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(G288), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1026), .A2(G8), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1026), .A2(G8), .A3(new_n1084), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(KEYINPUT52), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n922), .A2(G2090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n975), .A2(new_n976), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1008), .A2(new_n1072), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AND4_X1   g669(.A1(KEYINPUT113), .A2(new_n1094), .A3(G8), .A4(new_n1068), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1055), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT113), .B1(new_n1096), .B2(new_n1068), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1074), .B(new_n1090), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1066), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1002), .A2(new_n1050), .A3(new_n1062), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1062), .A2(KEYINPUT62), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1098), .A2(new_n999), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1058), .A2(new_n1103), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1097), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1096), .A2(KEYINPUT113), .A3(new_n1068), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1090), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1083), .A2(new_n1085), .A3(new_n678), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1075), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(G8), .A3(new_n1026), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1053), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1096), .A2(new_n1068), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1115), .A2(new_n1090), .A3(KEYINPUT115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1090), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1053), .A2(G8), .A3(G168), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1098), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1112), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1100), .A2(new_n1105), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G290), .B(G1986), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n923), .B1(new_n941), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n953), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT126), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(new_n953), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g708(.A1(G401), .A2(G229), .A3(new_n460), .A4(G227), .ZN(new_n1135));
  XOR2_X1   g709(.A(new_n1135), .B(KEYINPUT127), .Z(new_n1136));
  NAND3_X1  g710(.A1(new_n1136), .A2(new_n849), .A3(new_n904), .ZN(G225));
  INV_X1    g711(.A(G225), .ZN(G308));
endmodule


