//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n208), .B(new_n214), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n226), .B(new_n227), .Z(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G50), .B(G68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G58), .B(G77), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  NAND3_X1  g0039(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(new_n211), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT67), .ZN(new_n242));
  INV_X1    g0042(.A(G87), .ZN(new_n243));
  AND2_X1   g0043(.A1(new_n243), .A2(KEYINPUT15), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(KEYINPUT15), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT15), .B(G87), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n255), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n241), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT65), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT65), .A2(G1), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n262), .A2(G13), .A3(G20), .A4(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(KEYINPUT68), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT65), .B(G1), .Z(new_n268));
  AOI21_X1  g0068(.A(new_n241), .B1(new_n268), .B2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G77), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n264), .B2(G77), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n259), .A2(new_n267), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n277), .A2(G232), .B1(new_n280), .B2(G107), .ZN(new_n281));
  INV_X1    g0081(.A(G238), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n275), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  AND2_X1   g0088(.A1(G1), .A2(G13), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n262), .A2(new_n296), .A3(new_n263), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT66), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n262), .A2(new_n296), .A3(new_n299), .A4(new_n263), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n289), .A2(new_n290), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G244), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n287), .A2(new_n295), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n273), .A2(new_n274), .B1(new_n304), .B2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n241), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n246), .A2(new_n248), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n251), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n310), .B2(new_n257), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n270), .A2(new_n267), .A3(new_n272), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n311), .A2(new_n312), .A3(new_n274), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n304), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n304), .A2(G179), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n305), .A2(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n302), .A2(G226), .ZN(new_n320));
  INV_X1    g0120(.A(G223), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n284), .A2(new_n321), .B1(new_n266), .B2(new_n283), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G222), .B2(new_n277), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n295), .B(new_n320), .C1(new_n323), .C2(new_n301), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n316), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  INV_X1    g0126(.A(new_n256), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n254), .A2(new_n252), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G50), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n212), .B1(new_n201), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n241), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n269), .A2(G50), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n265), .A2(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n325), .B(new_n334), .C1(G179), .C2(new_n324), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n324), .A2(G200), .B1(new_n336), .B2(new_n334), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT9), .A4(new_n333), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n337), .B(new_n341), .C1(new_n306), .C2(new_n324), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(KEYINPUT10), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT10), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n324), .A2(new_n306), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n339), .B2(new_n340), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n346), .B2(new_n337), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n319), .B(new_n335), .C1(new_n343), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n225), .A2(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(G226), .B2(G1698), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n351), .B2(new_n280), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n286), .B1(new_n291), .B2(new_n294), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n298), .A2(G238), .A3(new_n300), .A4(new_n301), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT14), .B1(new_n358), .B2(new_n316), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n353), .A2(new_n355), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT13), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G68), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n251), .A2(G77), .B1(G20), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n256), .A2(G50), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n308), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g0171(.A(new_n371), .B(KEYINPUT11), .Z(new_n372));
  NAND2_X1  g0172(.A1(new_n265), .A2(new_n368), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n269), .A2(G68), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT71), .B1(new_n358), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n363), .A2(new_n380), .A3(G200), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n376), .B1(G190), .B2(new_n358), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n298), .A2(G232), .A3(new_n300), .A4(new_n301), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n295), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n295), .ZN(new_n390));
  INV_X1    g0190(.A(G1698), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n283), .A2(G223), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n283), .A2(G226), .A3(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G87), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(G190), .B1(new_n395), .B2(new_n286), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n286), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n295), .A3(new_n386), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n378), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n255), .A2(new_n264), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n269), .B2(new_n255), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n280), .B2(new_n212), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n278), .A2(new_n279), .A3(new_n406), .A4(G20), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G58), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n368), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n410), .B2(new_n201), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n256), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n308), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n404), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n401), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n275), .A2(new_n212), .A3(new_n276), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n406), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n368), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n416), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n418), .A3(new_n241), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n403), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n389), .A2(new_n430), .A3(new_n390), .A4(new_n398), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n399), .A2(new_n316), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT18), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n428), .A2(new_n403), .B1(new_n316), .B2(new_n399), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n431), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n401), .A2(new_n419), .A3(KEYINPUT17), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n422), .A2(new_n434), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n348), .A2(new_n385), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G116), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n240), .A2(new_n211), .B1(G20), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n443), .B(new_n212), .C1(G33), .C2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n442), .A2(KEYINPUT20), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT20), .B1(new_n442), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n262), .A2(G33), .A3(new_n263), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n264), .A2(new_n308), .A3(new_n449), .A4(G116), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n268), .A2(G13), .A3(G20), .A4(new_n441), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT77), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n445), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n442), .A2(KEYINPUT20), .A3(new_n445), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT77), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n451), .A4(new_n450), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(G264), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n462));
  OAI211_X1 g0262(.A(G257), .B(new_n391), .C1(new_n278), .C2(new_n279), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n465), .A2(new_n286), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n262), .A2(G45), .A3(new_n263), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G270), .B(new_n301), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n268), .A2(new_n291), .A3(G45), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n466), .A2(new_n474), .A3(new_n430), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n461), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT78), .ZN(new_n477));
  INV_X1    g0277(.A(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n465), .A2(new_n286), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n316), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n461), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G169), .B1(new_n466), .B2(new_n474), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n460), .B2(new_n453), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n485), .A2(new_n477), .A3(KEYINPUT21), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(new_n479), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n306), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n378), .B1(new_n478), .B2(new_n479), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n461), .A3(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n483), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n282), .A2(new_n391), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(G244), .B2(new_n391), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n493), .A2(new_n280), .B1(new_n250), .B2(new_n441), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n286), .ZN(new_n495));
  INV_X1    g0295(.A(G250), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n286), .B1(new_n467), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n262), .A2(G45), .A3(new_n288), .A4(new_n263), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n499), .A3(new_n306), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n286), .A2(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(G200), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n264), .A2(new_n308), .A3(new_n449), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G87), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n212), .B1(new_n349), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n243), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n212), .B(G68), .C1(new_n278), .C2(new_n279), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n506), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n506), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n308), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT75), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n264), .B1(new_n246), .B2(new_n248), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n506), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT74), .B1(new_n513), .B2(new_n506), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n511), .B(new_n510), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n241), .ZN(new_n526));
  INV_X1    g0326(.A(new_n521), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT75), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n502), .B(new_n505), .C1(new_n522), .C2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n501), .A2(new_n430), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G169), .B2(new_n501), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(KEYINPUT75), .A3(new_n527), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n309), .A2(new_n504), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT76), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT76), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n533), .A2(new_n534), .B1(new_n309), .B2(new_n504), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n529), .B(new_n539), .C1(new_n540), .C2(new_n532), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n268), .A2(G45), .A3(new_n472), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(G264), .A4(new_n301), .ZN(new_n545));
  OAI211_X1 g0345(.A(G264), .B(new_n301), .C1(new_n467), .C2(new_n470), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n549));
  OAI211_X1 g0349(.A(G250), .B(new_n391), .C1(new_n278), .C2(new_n279), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G294), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n467), .A2(new_n470), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n286), .B1(new_n553), .B2(new_n291), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n430), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n316), .B1(new_n554), .B2(new_n546), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n212), .B2(G107), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n559), .A2(new_n561), .B1(new_n251), .B2(G116), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n212), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n563));
  XNOR2_X1  g0363(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT24), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n563), .A2(new_n566), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(new_n562), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n308), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n264), .A2(G107), .ZN(new_n574));
  XOR2_X1   g0374(.A(KEYINPUT80), .B(KEYINPUT25), .Z(new_n575));
  OR2_X1    g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n577), .B1(G107), .B2(new_n504), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n556), .A2(new_n557), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n568), .A2(new_n572), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n241), .ZN(new_n582));
  AOI21_X1  g0382(.A(G200), .B1(new_n548), .B2(new_n554), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n554), .A2(new_n306), .A3(new_n546), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n578), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G250), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n586));
  OAI211_X1 g0386(.A(G244), .B(new_n391), .C1(new_n278), .C2(new_n279), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n443), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT4), .B1(new_n277), .B2(G244), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n286), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G257), .B(new_n301), .C1(new_n467), .C2(new_n470), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n592), .A2(new_n473), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n316), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n430), .A3(new_n593), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n327), .A2(new_n266), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT6), .ZN(new_n598));
  AND2_X1   g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n508), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n560), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n597), .B1(new_n602), .B2(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n424), .A2(new_n425), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(KEYINPUT73), .B1(new_n604), .B2(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT73), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n212), .B1(new_n600), .B2(new_n601), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n597), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n308), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n264), .A2(G97), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n444), .B2(new_n503), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n595), .B(new_n596), .C1(new_n609), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n602), .A2(G20), .ZN(new_n614));
  INV_X1    g0414(.A(new_n597), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(KEYINPUT73), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n604), .A2(G107), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n608), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n618), .B2(new_n241), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n594), .A2(G200), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n592), .A2(new_n473), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n587), .A2(new_n588), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(new_n443), .A4(new_n586), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n624), .B2(new_n286), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G190), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n619), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n580), .A2(new_n585), .A3(new_n613), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n440), .A2(new_n491), .A3(new_n542), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g0429(.A(new_n629), .B(KEYINPUT82), .Z(G372));
  AND3_X1   g0430(.A1(new_n435), .A2(new_n436), .A3(new_n431), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n436), .B1(new_n435), .B2(new_n431), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n361), .A2(G190), .A3(new_n362), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(new_n372), .A3(new_n374), .A4(new_n375), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n379), .B2(new_n381), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n317), .A2(new_n318), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n377), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n419), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT17), .B1(new_n401), .B2(new_n419), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n634), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n343), .A2(new_n347), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n335), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(G169), .B1(new_n591), .B2(new_n593), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n430), .B2(new_n625), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n618), .A2(new_n241), .ZN(new_n648));
  INV_X1    g0448(.A(new_n612), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT84), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n596), .B1(new_n625), .B2(G169), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT84), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n652), .A2(new_n619), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT83), .B1(new_n530), .B2(new_n537), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT83), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n529), .B(new_n657), .C1(new_n540), .C2(new_n532), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n613), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n542), .A2(KEYINPUT26), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT21), .B1(new_n485), .B2(new_n477), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n461), .A2(new_n480), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(KEYINPUT78), .A3(new_n482), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n667), .A3(new_n580), .A4(new_n476), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n613), .A2(new_n585), .A3(new_n627), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n656), .A3(new_n669), .A4(new_n658), .ZN(new_n670));
  INV_X1    g0470(.A(new_n537), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n645), .B1(new_n440), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT85), .Z(G369));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n665), .A2(new_n667), .A3(new_n476), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n212), .A2(G13), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n268), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n461), .A2(new_n684), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n677), .A2(new_n490), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n677), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n676), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n684), .B1(new_n579), .B2(new_n573), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n580), .A2(new_n585), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n580), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n694), .A2(KEYINPUT87), .A3(new_n684), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT87), .B1(new_n694), .B2(new_n684), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n684), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n677), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n699), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n206), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n509), .A2(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n209), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n684), .B1(new_n664), .B2(new_n672), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n659), .A2(KEYINPUT26), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n542), .A2(new_n660), .A3(new_n662), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n671), .A4(new_n670), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n699), .ZN(new_n715));
  MUX2_X1   g0515(.A(new_n711), .B(new_n715), .S(KEYINPUT29), .Z(new_n716));
  NAND4_X1  g0516(.A1(new_n542), .A2(new_n491), .A3(new_n628), .A4(new_n699), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n552), .A2(new_n286), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(new_n495), .A3(new_n499), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n475), .A2(new_n548), .A3(new_n719), .A4(new_n625), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n548), .A2(new_n501), .A3(new_n718), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .A3(new_n475), .A4(new_n625), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n501), .A2(G179), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n555), .A2(new_n725), .A3(new_n487), .A4(new_n594), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n727), .B2(new_n684), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n676), .B1(new_n717), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n716), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n710), .B1(new_n732), .B2(G1), .ZN(G364));
  AOI21_X1  g0533(.A(new_n261), .B1(new_n678), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n705), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n691), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n689), .A2(new_n676), .A3(new_n690), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n211), .B1(G20), .B2(new_n316), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n212), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n306), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n560), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n212), .A2(new_n430), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G190), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n378), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G20), .A3(new_n306), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G159), .ZN(new_n752));
  XOR2_X1   g0552(.A(KEYINPUT90), .B(KEYINPUT32), .Z(new_n753));
  OAI22_X1  g0553(.A1(new_n748), .A2(new_n329), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n744), .B(new_n754), .C1(G87), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n746), .A2(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n212), .B1(new_n749), .B2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G58), .B1(G97), .B2(new_n761), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n212), .A2(new_n430), .A3(new_n378), .A4(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n283), .B1(new_n764), .B2(new_n368), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n745), .A2(new_n306), .A3(new_n378), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G77), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n757), .A2(new_n758), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n747), .A2(G326), .B1(G294), .B2(new_n761), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT91), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n283), .B1(new_n767), .B2(G311), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  NOR2_X1   g0573(.A1(new_n764), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G329), .B2(new_n751), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n743), .B1(new_n755), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G322), .B2(new_n759), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n771), .A2(new_n772), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n741), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n736), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n740), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n235), .A2(new_n293), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n704), .A2(new_n283), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n293), .B2(new_n210), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n704), .A2(new_n280), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n441), .B2(new_n704), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n790), .A2(new_n793), .B1(KEYINPUT88), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(KEYINPUT88), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n789), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n781), .A2(new_n782), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n688), .B2(new_n786), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n739), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND3_X1  g0603(.A1(new_n317), .A2(new_n318), .A3(new_n699), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n314), .A2(new_n305), .B1(new_n273), .B2(new_n684), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n317), .A2(new_n318), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n711), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n717), .A2(new_n730), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G330), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n736), .B1(new_n809), .B2(new_n811), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n740), .A2(new_n783), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n736), .B1(G77), .B2(new_n816), .C1(new_n808), .C2(new_n784), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n743), .A2(new_n243), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n755), .A2(new_n560), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G294), .C2(new_n759), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n283), .B1(new_n767), .B2(G116), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n763), .A2(G283), .B1(new_n751), .B2(G311), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n747), .A2(G303), .B1(G97), .B2(new_n761), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n747), .A2(G137), .B1(G150), .B2(new_n763), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT92), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  INV_X1    g0627(.A(new_n759), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n826), .B1(new_n827), .B2(new_n828), .C1(new_n829), .C2(new_n766), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT93), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n283), .B1(new_n750), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT94), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n761), .A2(G58), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n743), .A2(new_n368), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G50), .B2(new_n756), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n833), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n832), .A2(KEYINPUT93), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n824), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT95), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n817), .B1(new_n844), .B2(new_n740), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n814), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  OR2_X1    g0647(.A1(new_n602), .A2(KEYINPUT35), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n602), .A2(KEYINPUT35), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n848), .A2(G116), .A3(new_n213), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT96), .B(KEYINPUT36), .Z(new_n851));
  XNOR2_X1  g0651(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OR3_X1    g0652(.A1(new_n209), .A2(new_n266), .A3(new_n410), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n329), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(G13), .B(new_n268), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n634), .A2(new_n682), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n376), .B(new_n684), .C1(new_n637), .C2(new_n367), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n376), .A2(new_n684), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n377), .A2(new_n384), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n684), .B(new_n807), .C1(new_n664), .C2(new_n672), .ZN(new_n862));
  INV_X1    g0662(.A(new_n804), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  INV_X1    g0665(.A(new_n682), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n429), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n633), .B2(new_n642), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT97), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n682), .B1(new_n428), .B2(new_n403), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n435), .B2(new_n431), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n420), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n420), .A2(new_n433), .A3(new_n867), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n872), .B2(KEYINPUT97), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n865), .B1(new_n868), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n439), .A2(new_n872), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n877), .A4(new_n874), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(KEYINPUT98), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT98), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(new_n865), .C1(new_n868), .C2(new_n878), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n857), .B1(new_n864), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n882), .B2(new_n884), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n367), .A2(new_n376), .A3(new_n699), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n875), .B(new_n869), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n865), .B1(new_n890), .B2(new_n868), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT39), .B1(new_n891), .B2(new_n881), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n645), .B1(new_n716), .B2(new_n440), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n881), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n807), .B1(new_n858), .B2(new_n860), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n810), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT40), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n810), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n884), .A3(new_n882), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n440), .A2(new_n810), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(G330), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n896), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n268), .B2(new_n678), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n896), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n856), .B1(new_n911), .B2(new_n912), .ZN(G367));
  OAI221_X1 g0713(.A(new_n788), .B1(new_n206), .B2(new_n249), .C1(new_n231), .C2(new_n792), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n782), .B1(new_n914), .B2(KEYINPUT104), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(KEYINPUT104), .B2(new_n914), .ZN(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT106), .B(G137), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n767), .A2(G50), .B1(new_n751), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n283), .C1(new_n829), .C2(new_n764), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n760), .A2(new_n368), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n743), .A2(new_n266), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n747), .A2(G143), .B1(new_n756), .B2(G58), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n326), .C2(new_n828), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n747), .A2(G311), .B1(G107), .B2(new_n761), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n444), .B2(new_n743), .C1(new_n777), .C2(new_n828), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT46), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n755), .A2(new_n927), .A3(new_n441), .ZN(new_n928));
  INV_X1    g0728(.A(G294), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n764), .A2(new_n929), .B1(new_n766), .B2(new_n776), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT46), .B1(new_n756), .B2(G116), .ZN(new_n931));
  XNOR2_X1  g0731(.A(KEYINPUT105), .B(G317), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n280), .B1(new_n932), .B2(new_n750), .ZN(new_n933));
  OR4_X1    g0733(.A1(new_n928), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n924), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n916), .B1(new_n936), .B2(new_n740), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n535), .A2(new_n505), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n684), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n656), .A2(new_n658), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n671), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n937), .B1(new_n941), .B2(new_n786), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n705), .B(new_n943), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n701), .A2(new_n702), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n613), .B(new_n627), .C1(new_n619), .C2(new_n699), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT99), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n662), .B2(new_n684), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT44), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n947), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n662), .A2(new_n684), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n701), .A3(new_n702), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT45), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n691), .A2(new_n697), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n697), .B(new_n700), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n691), .B(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n951), .A2(new_n957), .A3(new_n698), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n960), .A2(new_n732), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n944), .B1(new_n964), .B2(new_n732), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(new_n735), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT101), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n948), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n613), .B1(new_n952), .B2(new_n580), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n699), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT42), .B1(new_n948), .B2(new_n701), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT100), .Z(new_n976));
  AOI21_X1  g0776(.A(new_n969), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n967), .A2(new_n968), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n968), .A3(new_n967), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT102), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n959), .A2(new_n982), .A3(new_n954), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT102), .B1(new_n698), .B2(new_n948), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n981), .B(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n942), .B1(new_n966), .B2(new_n986), .ZN(G387));
  OR2_X1    g0787(.A1(new_n697), .A2(new_n786), .ZN(new_n988));
  INV_X1    g0788(.A(new_n794), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n989), .A2(new_n707), .B1(G107), .B2(new_n206), .ZN(new_n990));
  INV_X1    g0790(.A(new_n228), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n255), .A2(new_n329), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n707), .B(new_n293), .C1(new_n368), .C2(new_n266), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n791), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n991), .A2(G45), .B1(KEYINPUT107), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(KEYINPUT107), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n736), .B1(new_n998), .B2(new_n789), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n767), .A2(G303), .B1(new_n763), .B2(G311), .ZN(new_n1000));
  INV_X1    g0800(.A(G322), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n748), .B2(new_n1001), .C1(new_n828), .C2(new_n932), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n755), .A2(new_n929), .B1(new_n760), .B2(new_n776), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT109), .Z(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n743), .A2(new_n441), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n283), .B(new_n1012), .C1(G326), .C2(new_n751), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n828), .A2(new_n329), .B1(new_n743), .B2(new_n444), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n748), .A2(new_n829), .B1(new_n755), .B2(new_n266), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n309), .A2(new_n761), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT108), .B(G150), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n280), .B1(new_n751), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n767), .A2(G68), .B1(new_n763), .B2(new_n255), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n999), .B1(new_n1023), .B2(new_n740), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n962), .A2(new_n735), .B1(new_n988), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n962), .A2(new_n732), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n705), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n962), .A2(new_n732), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  NAND2_X1  g0829(.A1(new_n948), .A2(new_n787), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n788), .B1(new_n444), .B2(new_n206), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n238), .A2(new_n792), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n736), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT110), .Z(new_n1034));
  AOI22_X1  g0834(.A1(G311), .A2(new_n759), .B1(new_n747), .B2(G317), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT52), .Z(new_n1036));
  OAI22_X1  g0836(.A1(new_n764), .A2(new_n777), .B1(new_n760), .B2(new_n441), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT112), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n280), .B1(new_n750), .B2(new_n1001), .C1(new_n766), .C2(new_n929), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n744), .B(new_n1041), .C1(G283), .C2(new_n756), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G150), .A2(new_n747), .B1(new_n759), .B2(G159), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n766), .A2(new_n254), .B1(new_n750), .B2(new_n827), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n280), .B(new_n1047), .C1(G50), .C2(new_n763), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n760), .A2(new_n266), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1049), .B(new_n818), .C1(G68), .C2(new_n756), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1043), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT113), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n741), .B1(new_n1053), .B2(KEYINPUT113), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1034), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1030), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n960), .A2(new_n963), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n734), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n964), .A2(new_n705), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1026), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G390));
  OAI21_X1  g0863(.A(new_n736), .B1(new_n255), .B2(new_n816), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT116), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n283), .B1(new_n763), .B2(G107), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n444), .B2(new_n766), .C1(new_n929), .C2(new_n750), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n838), .B(new_n1067), .C1(G87), .C2(new_n756), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n748), .A2(new_n776), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1049), .B(new_n1069), .C1(G116), .C2(new_n759), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n756), .A2(new_n1019), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT53), .Z(new_n1072));
  AOI22_X1  g0872(.A1(new_n763), .A2(new_n917), .B1(new_n751), .B2(G125), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT54), .B(G143), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n283), .C1(new_n766), .C2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n828), .A2(new_n834), .B1(new_n760), .B2(new_n829), .ZN(new_n1076));
  INV_X1    g0876(.A(G128), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n748), .A2(new_n1077), .B1(new_n743), .B2(new_n329), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1068), .A2(new_n1070), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1065), .B1(new_n1080), .B2(new_n741), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n892), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1084), .B2(new_n783), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n731), .A2(new_n808), .A3(new_n861), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1086), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n864), .A2(new_n889), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n897), .A2(new_n889), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n714), .B(new_n699), .C1(new_n806), .C2(new_n805), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n804), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(new_n861), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1088), .B(new_n1092), .C1(new_n1093), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n861), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n673), .A2(new_n699), .A3(new_n808), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n804), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n889), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1101), .A2(new_n1102), .B1(new_n888), .B2(new_n892), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1096), .A2(new_n861), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1094), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1103), .A2(new_n1106), .A3(new_n1090), .A4(new_n1089), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1085), .B1(new_n1108), .B2(new_n735), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n440), .A2(new_n731), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT115), .Z(new_n1111));
  AOI21_X1  g0911(.A(new_n861), .B1(new_n731), .B2(new_n808), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1089), .A2(new_n1112), .B1(new_n862), .B2(new_n863), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1099), .B1(new_n811), .B2(new_n807), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1114), .A2(new_n804), .A3(new_n1086), .A4(new_n1095), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n895), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n705), .B1(new_n1108), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n1098), .B2(new_n1107), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1109), .B1(new_n1119), .B2(new_n1120), .ZN(G378));
  AOI21_X1  g0921(.A(new_n676), .B1(new_n901), .B2(new_n904), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n886), .B2(new_n893), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n885), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1101), .A2(new_n1124), .B1(new_n634), .B2(new_n682), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n903), .A2(new_n884), .A3(new_n882), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n900), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n902), .B1(new_n1127), .B2(new_n897), .ZN(new_n1128));
  OAI21_X1  g0928(.A(G330), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1082), .A2(new_n1102), .A3(new_n1083), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n343), .A2(new_n347), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n335), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n866), .A2(new_n334), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT118), .Z(new_n1135));
  XNOR2_X1  g0935(.A(new_n1133), .B(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1123), .A2(new_n1131), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n735), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n828), .A2(new_n560), .B1(new_n743), .B2(new_n409), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G116), .B2(new_n747), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n309), .A2(new_n767), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n280), .A2(new_n292), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n750), .A2(new_n776), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(G97), .C2(new_n763), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n920), .B1(G77), .B2(new_n756), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT58), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1146), .B(new_n329), .C1(G33), .C2(G41), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT117), .Z(new_n1155));
  AOI211_X1 g0955(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n829), .B2(new_n743), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n755), .A2(new_n1074), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n764), .A2(new_n834), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G137), .C2(new_n767), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n747), .A2(G125), .B1(G150), .B2(new_n761), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n1077), .C2(new_n828), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1157), .B1(new_n1162), .B2(KEYINPUT59), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(KEYINPUT59), .B2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n740), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n782), .B1(new_n329), .B2(new_n815), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n1138), .C2(new_n784), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1142), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1123), .A2(new_n1131), .A3(new_n1138), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1138), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n886), .A2(new_n1122), .A3(new_n893), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1129), .B1(new_n1130), .B2(new_n1125), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n895), .A2(new_n1111), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1171), .B(new_n1175), .C1(new_n1120), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  OAI211_X1 g0978(.A(KEYINPUT119), .B(new_n705), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1087), .B(new_n1091), .C1(new_n1103), .C2(new_n1106), .ZN(new_n1182));
  AND4_X1   g0982(.A1(new_n1090), .A2(new_n1103), .A3(new_n1089), .A4(new_n1106), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1118), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1176), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1141), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT119), .B1(new_n1187), .B2(new_n705), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1170), .B1(new_n1181), .B2(new_n1188), .ZN(G375));
  AOI21_X1  g0989(.A(new_n782), .B1(new_n368), .B2(new_n815), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n283), .B1(new_n751), .B2(G303), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n767), .A2(G107), .B1(new_n763), .B2(G116), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1018), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n828), .A2(new_n776), .B1(new_n748), .B2(new_n929), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n755), .A2(new_n444), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n921), .A4(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT121), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n748), .A2(new_n834), .B1(new_n743), .B2(new_n409), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n283), .B1(new_n764), .B2(new_n1074), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n766), .A2(new_n326), .B1(new_n750), .B2(new_n1077), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n759), .A2(new_n917), .B1(G50), .B2(new_n761), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n829), .C2(new_n755), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1197), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(KEYINPUT121), .B2(new_n1196), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1190), .B1(new_n741), .B2(new_n1205), .C1(new_n861), .C2(new_n784), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n734), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(KEYINPUT120), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(KEYINPUT120), .B2(new_n1207), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1116), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1176), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n944), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1117), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1213), .ZN(G381));
  INV_X1    g1014(.A(G387), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n802), .B(new_n1025), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1215), .A2(new_n846), .A3(new_n1062), .A4(new_n1217), .ZN(new_n1218));
  OR4_X1    g1018(.A1(G378), .A2(G375), .A3(new_n1218), .A4(G381), .ZN(G407));
  NAND2_X1  g1019(.A1(new_n683), .A2(G213), .ZN(new_n1220));
  OR3_X1    g1020(.A1(G375), .A2(G378), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(new_n1220), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G378), .B(new_n1170), .C1(new_n1181), .C2(new_n1188), .ZN(new_n1226));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1177), .A2(new_n944), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1169), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1232), .A2(new_n1211), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n705), .B1(new_n1232), .B2(new_n1211), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1209), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n846), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G384), .B(new_n1209), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1230), .A2(new_n1231), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1236), .A2(KEYINPUT123), .A3(new_n1238), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1225), .A2(G2897), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT123), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1242), .B1(new_n1230), .B2(new_n1250), .ZN(new_n1251));
  XOR2_X1   g1051(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1230), .B2(new_n1240), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1241), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(new_n1217), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n983), .A2(new_n984), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n981), .B(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n735), .B2(new_n965), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1259), .A2(new_n942), .A3(new_n1062), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1062), .B1(new_n1259), .B2(new_n942), .ZN(new_n1261));
  OAI211_X1 g1061(.A(KEYINPUT125), .B(new_n1256), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(G390), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1256), .A2(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1259), .A2(new_n942), .A3(new_n1062), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1255), .B2(new_n1217), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1230), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1250), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(KEYINPUT124), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1220), .A3(new_n1240), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1230), .A2(KEYINPUT63), .A3(new_n1240), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1273), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1262), .A2(new_n1242), .A3(new_n1268), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1262), .A2(new_n1268), .A3(KEYINPUT126), .A4(new_n1242), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1230), .A2(new_n1250), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1284), .B1(KEYINPUT124), .B2(new_n1285), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1254), .A2(new_n1270), .B1(new_n1279), .B2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1227), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1226), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(new_n1240), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1240), .ZN(new_n1291));
  OR3_X1    g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1269), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1269), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(G402));
endmodule


