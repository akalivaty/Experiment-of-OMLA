//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT86), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n220), .C1(KEYINPUT15), .C2(new_n208), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n211), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(KEYINPUT84), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n214), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(KEYINPUT83), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n228), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n223), .A2(new_n226), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n206), .B1(new_n230), .B2(new_n220), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT17), .B1(new_n222), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n214), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n233), .A2(KEYINPUT14), .B1(new_n224), .B2(new_n214), .ZN(new_n234));
  NAND2_X1  g033(.A1(G29gat), .A2(G36gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT85), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n207), .A4(new_n210), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n243));
  INV_X1    g042(.A(new_n226), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n225), .B1(new_n224), .B2(new_n214), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n227), .A2(new_n229), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n239), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n242), .B(new_n243), .C1(new_n248), .C2(new_n206), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G99gat), .B(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT96), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G85gat), .A3(G92gat), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT7), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT7), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(KEYINPUT96), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G85gat), .ZN(new_n260));
  INV_X1    g059(.A(G92gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT8), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n252), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT7), .ZN(new_n267));
  AOI22_X1  g066(.A1(KEYINPUT8), .A2(new_n263), .B1(new_n260), .B2(new_n261), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n251), .A3(new_n259), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT97), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n222), .A2(new_n231), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n266), .A2(new_n269), .ZN(new_n276));
  AND2_X1   g075(.A1(G232gat), .A2(G233gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n275), .A2(new_n276), .B1(KEYINPUT41), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G190gat), .B(G218gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(KEYINPUT98), .A3(new_n283), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n279), .A2(KEYINPUT98), .A3(new_n280), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT99), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n277), .A2(KEYINPUT41), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(G134gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n284), .A2(new_n285), .A3(new_n288), .A4(new_n292), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G8gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT88), .ZN(new_n298));
  INV_X1    g097(.A(G1gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT87), .A3(KEYINPUT16), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT16), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(G1gat), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G15gat), .ZN(new_n305));
  INV_X1    g104(.A(G15gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G22gat), .ZN(new_n307));
  AND4_X1   g106(.A1(new_n300), .A2(new_n303), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n297), .A2(KEYINPUT88), .ZN(new_n309));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n298), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n300), .A3(new_n303), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(new_n307), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G1gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n298), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .A4(new_n309), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G71gat), .B(G78gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n322));
  AND2_X1   g121(.A1(G57gat), .A2(G64gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G57gat), .A2(G64gat), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  XNOR2_X1  g127(.A(G57gat), .B(G64gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n320), .B(new_n328), .C1(new_n329), .C2(new_n322), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n319), .B1(KEYINPUT21), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n327), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G155gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g137(.A1(G231gat), .A2(G233gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT95), .ZN(new_n340));
  XOR2_X1   g139(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G183gat), .B(G211gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n337), .A2(new_n338), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n344), .B1(new_n337), .B2(new_n338), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n296), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G230gat), .A2(G233gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT101), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n269), .A2(KEYINPUT100), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n276), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n270), .A2(new_n331), .A3(new_n352), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT10), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n276), .A2(KEYINPUT10), .A3(new_n331), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n351), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT102), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT102), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n351), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n350), .A3(new_n355), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G120gat), .B(G148gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G176gat), .B(G204gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n359), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT103), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT103), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n359), .A2(new_n371), .A3(new_n361), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n358), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n367), .B1(new_n374), .B2(new_n363), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n348), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT37), .ZN(new_n379));
  OR2_X1    g178(.A1(G197gat), .A2(G204gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(G197gat), .A2(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  NAND2_X1  g181(.A1(G211gat), .A2(G218gat), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT72), .ZN(new_n385));
  INV_X1    g184(.A(new_n383), .ZN(new_n386));
  NOR2_X1   g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n385), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G226gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n395), .A2(KEYINPUT23), .ZN(new_n396));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(KEYINPUT23), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT66), .B(G183gat), .ZN(new_n400));
  INV_X1    g199(.A(G190gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT67), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n404), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407));
  INV_X1    g206(.A(G183gat), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n407), .A2(new_n408), .A3(new_n401), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n410), .A2(KEYINPUT65), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(KEYINPUT65), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n399), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT26), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n418), .A2(new_n395), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n395), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n408), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n400), .B2(new_n422), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n401), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT28), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT27), .B(G183gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT28), .A3(new_n401), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n421), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n409), .B1(new_n408), .B2(new_n401), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n410), .A2(KEYINPUT64), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n410), .A2(KEYINPUT64), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n399), .A2(KEYINPUT25), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n394), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n414), .B2(new_n415), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n430), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n442), .A2(new_n392), .A3(new_n393), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n391), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n394), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n442), .A2(KEYINPUT29), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n390), .B(new_n445), .C1(new_n446), .C2(new_n394), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT73), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(KEYINPUT73), .A3(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n379), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT79), .B(KEYINPUT37), .Z(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT38), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n454), .A2(new_n461), .A3(new_n458), .A4(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464));
  XNOR2_X1  g263(.A(G141gat), .B(G148gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n466), .A2(KEYINPUT2), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G155gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n291), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT74), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(KEYINPUT74), .A3(new_n466), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n472), .B(new_n471), .C1(new_n465), .C2(new_n467), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G113gat), .B(G120gat), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(KEYINPUT1), .ZN(new_n480));
  XNOR2_X1  g279(.A(G127gat), .B(G134gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n478), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n477), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n482), .A2(new_n477), .A3(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n478), .A2(KEYINPUT3), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n482), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n491), .A2(new_n485), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n496), .A2(new_n489), .A3(new_n485), .A4(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(new_n497), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n486), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G1gat), .B(G29gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT0), .ZN(new_n504));
  XNOR2_X1  g303(.A(G57gat), .B(G85gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n464), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  AOI211_X1 g307(.A(new_n506), .B(new_n486), .C1(new_n498), .C2(new_n501), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n502), .A2(KEYINPUT6), .A3(new_n507), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n458), .B1(new_n444), .B2(new_n447), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n460), .A2(new_n463), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n493), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n478), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n439), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n390), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(G228gat), .A3(G233gat), .A4(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n384), .A2(new_n388), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n439), .B1(new_n384), .B2(new_n388), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n493), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n478), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n518), .A2(new_n523), .B1(G228gat), .B2(G233gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G78gat), .B(G106gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n202), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n532), .A2(new_n533), .A3(new_n304), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n304), .B2(new_n532), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n528), .A2(new_n535), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n444), .A2(KEYINPUT73), .A3(new_n447), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT73), .B1(new_n444), .B2(new_n447), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n458), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n491), .A2(new_n496), .ZN(new_n547));
  INV_X1    g346(.A(new_n485), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n483), .A2(new_n485), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n549), .A2(KEYINPUT39), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT39), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n552), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n506), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n546), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n509), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(KEYINPUT39), .A3(new_n550), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n557), .A2(KEYINPUT40), .A3(new_n506), .A4(new_n553), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n539), .B1(new_n545), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n508), .A2(new_n509), .ZN(new_n561));
  INV_X1    g360(.A(new_n511), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n512), .B(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n542), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n514), .A2(new_n560), .B1(new_n566), .B2(new_n539), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n416), .A2(KEYINPUT68), .A3(new_n431), .A4(new_n437), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n441), .B2(new_n430), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n495), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n438), .A2(new_n569), .A3(new_n482), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G227gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n393), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT34), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n575), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n571), .A2(KEYINPUT70), .A3(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT34), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n582), .B2(KEYINPUT34), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT32), .B1(new_n573), .B2(new_n580), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n573), .B2(new_n580), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G99gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT69), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n306), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G43gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  OAI221_X1 g394(.A(KEYINPUT32), .B1(new_n588), .B2(new_n593), .C1(new_n573), .C2(new_n580), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n582), .A2(KEYINPUT34), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT71), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT34), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n597), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n577), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n598), .A2(new_n604), .A3(KEYINPUT36), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT36), .B1(new_n598), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n567), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n586), .A2(new_n597), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n603), .B1(new_n602), .B2(new_n577), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n566), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n610), .A2(KEYINPUT35), .A3(new_n611), .A4(new_n538), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n538), .A3(new_n604), .A4(new_n598), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT35), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g416(.A(G169gat), .B(G197gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT81), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n618), .B(KEYINPUT81), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n617), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n625), .A3(new_n617), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  INV_X1    g430(.A(new_n628), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n626), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n222), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n230), .A2(new_n220), .ZN(new_n636));
  INV_X1    g435(.A(new_n206), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n243), .B1(new_n638), .B2(new_n242), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n318), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n317), .B(new_n312), .C1(new_n222), .C2(new_n231), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n640), .A2(KEYINPUT18), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n318), .A2(new_n638), .A3(new_n242), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n642), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n641), .B(KEYINPUT13), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT89), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(KEYINPUT89), .A3(new_n646), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n643), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n634), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT91), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n319), .B1(new_n232), .B2(new_n249), .ZN(new_n658));
  INV_X1    g457(.A(new_n641), .ZN(new_n659));
  INV_X1    g458(.A(new_n642), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n661), .A2(KEYINPUT90), .A3(KEYINPUT18), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT90), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n652), .B2(new_n653), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AND4_X1   g464(.A1(new_n634), .A2(new_n643), .A3(new_n649), .A4(new_n650), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n657), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT90), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n663), .A3(new_n653), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n643), .A2(new_n649), .A3(new_n634), .A4(new_n650), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n670), .A2(KEYINPUT91), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n656), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n616), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT92), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n616), .A2(KEYINPUT92), .A3(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n378), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n563), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND3_X1   g481(.A1(new_n678), .A2(new_n545), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n297), .B1(new_n678), .B2(new_n545), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  NAND3_X1  g485(.A1(new_n678), .A2(new_n306), .A3(new_n610), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT36), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n608), .B2(new_n609), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n598), .A2(new_n604), .A3(KEYINPUT36), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n678), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n687), .B1(new_n694), .B2(new_n306), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n539), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  NAND2_X1  g497(.A1(new_n377), .A2(new_n347), .ZN(new_n699));
  INV_X1    g498(.A(new_n296), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT104), .Z(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n676), .B2(new_n677), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n213), .A3(new_n679), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n616), .A2(new_n296), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n616), .A2(KEYINPUT44), .A3(new_n296), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT91), .B1(new_n670), .B2(new_n671), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n666), .A2(new_n657), .A3(new_n668), .A4(new_n669), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n655), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n563), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n705), .A2(new_n706), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n707), .A2(new_n718), .A3(new_n719), .ZN(G1328gat));
  INV_X1    g519(.A(new_n545), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(G36gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n717), .B2(new_n721), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(G1329gat));
  NAND2_X1  g531(.A1(new_n704), .A2(new_n610), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n204), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n712), .A2(G43gat), .A3(new_n692), .A4(new_n716), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT47), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1330gat));
  NAND2_X1  g539(.A1(new_n704), .A2(new_n539), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n202), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n712), .A2(G50gat), .A3(new_n539), .A4(new_n716), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1331gat));
  NAND3_X1  g547(.A1(new_n348), .A2(new_n715), .A3(new_n376), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n691), .A2(new_n567), .B1(new_n614), .B2(new_n613), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n612), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n679), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n545), .B(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756));
  INV_X1    g555(.A(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT107), .Z(new_n759));
  NAND2_X1  g558(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n757), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1333gat));
  NAND2_X1  g561(.A1(new_n751), .A2(new_n610), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  AOI21_X1  g563(.A(G71gat), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n751), .A2(G71gat), .A3(new_n692), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT50), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n751), .A2(new_n539), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  INV_X1    g573(.A(new_n347), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n673), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n616), .A2(new_n296), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n616), .A2(KEYINPUT51), .A3(new_n296), .A4(new_n776), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n376), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n679), .A2(new_n260), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n673), .A2(new_n377), .A3(new_n775), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n710), .A2(new_n711), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n679), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n787), .A2(new_n788), .B1(new_n260), .B2(new_n791), .ZN(G1336gat));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n779), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n700), .B1(new_n750), .B2(new_n612), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n785), .A3(KEYINPUT51), .A4(new_n776), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n795), .A2(new_n780), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n755), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(G92gat), .A3(new_n377), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n793), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT111), .B(new_n801), .C1(new_n783), .C2(new_n786), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n710), .A2(new_n711), .A3(new_n755), .A4(new_n789), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n805), .B2(G92gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n798), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n802), .B1(new_n808), .B2(new_n794), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n261), .B1(new_n790), .B2(new_n545), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(G1337gat));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n692), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G99gat), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n813), .A2(new_n814), .ZN(new_n817));
  INV_X1    g616(.A(new_n610), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(G99gat), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n816), .A2(new_n817), .B1(new_n787), .B2(new_n819), .ZN(G1338gat));
  NAND4_X1  g619(.A1(new_n710), .A2(new_n539), .A3(new_n711), .A4(new_n789), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n821), .B2(G106gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n377), .A2(new_n538), .A3(G106gat), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n799), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n794), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n824), .B(KEYINPUT114), .Z(new_n827));
  AOI22_X1  g626(.A1(new_n826), .A2(new_n827), .B1(G106gat), .B2(new_n821), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n356), .A2(new_n357), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n350), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n359), .A3(new_n361), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n366), .B1(new_n374), .B2(new_n831), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT55), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n373), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n834), .B2(new_n835), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n715), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n713), .A2(new_n714), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n645), .A2(new_n646), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT115), .Z(new_n842));
  AOI21_X1  g641(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n628), .B(new_n627), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n376), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n700), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n838), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n296), .A2(new_n373), .A3(new_n847), .A4(new_n836), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n840), .A2(new_n844), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n775), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n378), .A2(new_n673), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT116), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  INV_X1    g653(.A(new_n852), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n848), .A2(new_n849), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n373), .A2(new_n836), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n673), .A2(new_n857), .A3(new_n847), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n376), .A2(new_n840), .A3(new_n844), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n700), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n854), .B(new_n855), .C1(new_n861), .C2(new_n775), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n539), .A3(new_n818), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n755), .A2(new_n563), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n673), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n376), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n775), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n721), .A2(new_n296), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G134gat), .A3(new_n563), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT117), .Z(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n866), .A2(new_n296), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G134gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(G1343gat));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n853), .A2(new_n539), .A3(new_n862), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G141gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n691), .A2(new_n865), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n673), .A4(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n538), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n834), .A2(new_n835), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(new_n892), .B2(KEYINPUT119), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(KEYINPUT119), .B2(new_n892), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n673), .A3(new_n857), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n296), .B1(new_n895), .B2(new_n859), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n347), .B1(new_n896), .B2(new_n856), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n852), .B1(new_n897), .B2(KEYINPUT120), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(KEYINPUT120), .B2(new_n897), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n890), .A2(KEYINPUT118), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n901), .A3(new_n889), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n886), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(new_n673), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n882), .B(new_n888), .C1(new_n904), .C2(new_n885), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n885), .B1(new_n903), .B2(new_n673), .ZN(new_n906));
  INV_X1    g705(.A(new_n888), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT58), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(G1344gat));
  XOR2_X1   g708(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n910));
  INV_X1    g709(.A(new_n891), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n538), .B1(new_n897), .B2(new_n855), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n863), .A2(new_n911), .B1(new_n912), .B2(KEYINPUT57), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n376), .A3(new_n887), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n890), .A2(KEYINPUT118), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n891), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n902), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n376), .A3(new_n887), .ZN(new_n919));
  INV_X1    g718(.A(G148gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT59), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n884), .A2(new_n920), .A3(new_n376), .A4(new_n887), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT122), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  INV_X1    g725(.A(new_n921), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n903), .B2(new_n376), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n926), .B(new_n923), .C1(new_n928), .C2(new_n915), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(G1345gat));
  AND2_X1   g729(.A1(new_n903), .A2(new_n775), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n884), .A2(new_n887), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n775), .A2(new_n469), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n931), .A2(new_n469), .B1(new_n932), .B2(new_n933), .ZN(G1346gat));
  AND2_X1   g733(.A1(new_n903), .A2(new_n296), .ZN(new_n935));
  OR4_X1    g734(.A1(G162gat), .A2(new_n692), .A3(new_n563), .A4(new_n873), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n935), .A2(new_n291), .B1(new_n883), .B2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n863), .A2(new_n679), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n818), .A2(new_n539), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(G169gat), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n673), .A4(new_n755), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n938), .A2(new_n545), .A3(new_n939), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n715), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n945), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT123), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n942), .B(new_n948), .C1(new_n945), .C2(new_n941), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1348gat));
  NAND2_X1  g749(.A1(new_n940), .A2(new_n755), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n951), .A2(G176gat), .A3(new_n377), .ZN(new_n952));
  OAI21_X1  g751(.A(G176gat), .B1(new_n944), .B2(new_n377), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n944), .A2(new_n347), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n775), .A2(new_n428), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n955), .A2(new_n400), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  OAI221_X1 g758(.A(new_n959), .B1(new_n951), .B2(new_n956), .C1(new_n955), .C2(new_n400), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1350gat));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n943), .A2(new_n296), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n401), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT124), .B(G190gat), .C1(new_n944), .C2(new_n700), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(KEYINPUT61), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n962), .B(new_n967), .C1(new_n963), .C2(new_n401), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n940), .A2(new_n401), .A3(new_n296), .A4(new_n755), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(G1351gat));
  NOR3_X1   g769(.A1(new_n692), .A2(new_n679), .A3(new_n721), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n913), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(G197gat), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n972), .A2(new_n973), .A3(new_n715), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n692), .A2(new_n538), .A3(new_n800), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n938), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n938), .A2(KEYINPUT125), .A3(new_n975), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n673), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n974), .B1(new_n981), .B2(new_n973), .ZN(G1352gat));
  OAI21_X1  g781(.A(G204gat), .B1(new_n972), .B2(new_n377), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n976), .A2(G204gat), .A3(new_n377), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT126), .A3(new_n984), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT126), .B1(new_n985), .B2(new_n984), .ZN(new_n987));
  OAI221_X1 g786(.A(new_n983), .B1(new_n984), .B2(new_n985), .C1(new_n986), .C2(new_n987), .ZN(G1353gat));
  OAI21_X1  g787(.A(G211gat), .B1(new_n972), .B2(new_n347), .ZN(new_n989));
  XOR2_X1   g788(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  INV_X1    g789(.A(G211gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n980), .A2(new_n991), .A3(new_n775), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1354gat));
  NOR2_X1   g792(.A1(new_n700), .A2(G218gat), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n913), .A2(new_n296), .A3(new_n971), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n996), .A2(G218gat), .ZN(new_n997));
  OR3_X1    g796(.A1(new_n995), .A2(KEYINPUT127), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(KEYINPUT127), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1355gat));
endmodule


