

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753;

  XNOR2_X1 U372 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n380) );
  INV_X1 U373 ( .A(G953), .ZN(n745) );
  NOR2_X1 U374 ( .A1(n720), .A2(n597), .ZN(n593) );
  XNOR2_X1 U375 ( .A(n548), .B(KEYINPUT35), .ZN(n566) );
  BUF_X1 U376 ( .A(G128), .Z(n349) );
  AND2_X2 U377 ( .A1(n363), .A2(n744), .ZN(n624) );
  NAND2_X2 U378 ( .A1(n661), .A2(n623), .ZN(n363) );
  XNOR2_X1 U379 ( .A(n512), .B(n365), .ZN(n552) );
  XNOR2_X1 U380 ( .A(G119), .B(G113), .ZN(n376) );
  XNOR2_X1 U381 ( .A(G101), .B(KEYINPUT67), .ZN(n375) );
  BUF_X1 U382 ( .A(n487), .Z(n350) );
  XNOR2_X1 U383 ( .A(n351), .B(n352), .ZN(n482) );
  NOR2_X1 U384 ( .A1(n653), .A2(n444), .ZN(n351) );
  NAND2_X1 U385 ( .A1(n445), .A2(G210), .ZN(n352) );
  XNOR2_X2 U386 ( .A(n353), .B(KEYINPUT0), .ZN(n543) );
  NOR2_X2 U387 ( .A1(n598), .A2(n507), .ZN(n353) );
  XNOR2_X2 U388 ( .A(n354), .B(G469), .ZN(n487) );
  NOR2_X2 U389 ( .A1(n672), .A2(G902), .ZN(n354) );
  XNOR2_X2 U390 ( .A(n433), .B(n381), .ZN(n741) );
  XNOR2_X2 U391 ( .A(n380), .B(n450), .ZN(n433) );
  XNOR2_X2 U392 ( .A(n397), .B(n396), .ZN(n672) );
  XNOR2_X2 U393 ( .A(n741), .B(G146), .ZN(n397) );
  NOR2_X1 U394 ( .A1(n594), .A2(n753), .ZN(n596) );
  NAND2_X1 U395 ( .A1(n356), .A2(n565), .ZN(n359) );
  BUF_X1 U396 ( .A(n517), .Z(n585) );
  AND2_X1 U397 ( .A1(n622), .A2(n621), .ZN(n744) );
  INV_X1 U398 ( .A(KEYINPUT22), .ZN(n365) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n460) );
  XNOR2_X1 U400 ( .A(n596), .B(n366), .ZN(n616) );
  XNOR2_X1 U401 ( .A(G146), .B(G125), .ZN(n435) );
  XNOR2_X1 U402 ( .A(n483), .B(KEYINPUT85), .ZN(n502) );
  NAND2_X1 U403 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U404 ( .A(n413), .B(n412), .ZN(n517) );
  XNOR2_X1 U405 ( .A(n502), .B(KEYINPUT19), .ZN(n598) );
  XNOR2_X1 U406 ( .A(G104), .B(G107), .ZN(n392) );
  XNOR2_X1 U407 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U408 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U409 ( .A(n538), .B(n364), .ZN(n556) );
  INV_X1 U410 ( .A(KEYINPUT103), .ZN(n364) );
  XOR2_X1 U411 ( .A(n401), .B(n400), .Z(n355) );
  AND2_X1 U412 ( .A1(n564), .A2(n563), .ZN(n356) );
  AND2_X1 U413 ( .A1(n551), .A2(n515), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n579), .B(KEYINPUT45), .ZN(n358) );
  NAND2_X1 U415 ( .A1(n360), .A2(n359), .ZN(n578) );
  NAND2_X1 U416 ( .A1(n362), .A2(n361), .ZN(n360) );
  AND2_X1 U417 ( .A1(n561), .A2(n565), .ZN(n361) );
  NOR2_X1 U418 ( .A1(n564), .A2(KEYINPUT65), .ZN(n362) );
  NAND2_X1 U419 ( .A1(n363), .A2(n628), .ZN(n629) );
  XNOR2_X1 U420 ( .A(n556), .B(G110), .ZN(G12) );
  NAND2_X1 U421 ( .A1(n552), .A2(n357), .ZN(n572) );
  INV_X1 U422 ( .A(n482), .ZN(n480) );
  XNOR2_X1 U423 ( .A(n443), .B(n668), .ZN(n653) );
  XOR2_X1 U424 ( .A(n595), .B(KEYINPUT46), .Z(n366) );
  AND2_X1 U425 ( .A1(n685), .A2(n537), .ZN(n367) );
  AND2_X1 U426 ( .A1(n551), .A2(n550), .ZN(n368) );
  INV_X1 U427 ( .A(G137), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n379) );
  INV_X1 U430 ( .A(KEYINPUT34), .ZN(n544) );
  BUF_X1 U431 ( .A(n516), .Z(n685) );
  AND2_X1 U432 ( .A1(n430), .A2(n429), .ZN(n498) );
  BUF_X1 U433 ( .A(n566), .Z(n558) );
  XOR2_X1 U434 ( .A(KEYINPUT5), .B(KEYINPUT72), .Z(n370) );
  NAND2_X1 U435 ( .A1(n460), .A2(G210), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n374) );
  XNOR2_X1 U437 ( .A(G116), .B(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n378) );
  XNOR2_X1 U439 ( .A(KEYINPUT88), .B(KEYINPUT3), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n441) );
  XNOR2_X1 U441 ( .A(n379), .B(n441), .ZN(n382) );
  XNOR2_X2 U442 ( .A(G143), .B(G128), .ZN(n450) );
  XNOR2_X1 U443 ( .A(G134), .B(G131), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n397), .ZN(n639) );
  INV_X1 U445 ( .A(G902), .ZN(n457) );
  NAND2_X1 U446 ( .A1(n639), .A2(n457), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n383), .B(G472), .ZN(n522) );
  INV_X1 U448 ( .A(G237), .ZN(n384) );
  NAND2_X1 U449 ( .A1(n457), .A2(n384), .ZN(n445) );
  AND2_X1 U450 ( .A1(n445), .A2(G214), .ZN(n490) );
  NAND2_X1 U451 ( .A1(n522), .A2(n481), .ZN(n386) );
  INV_X1 U452 ( .A(KEYINPUT30), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n430) );
  NAND2_X1 U454 ( .A1(n745), .A2(G227), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n387), .B(KEYINPUT90), .ZN(n390) );
  INV_X1 U456 ( .A(G140), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n388), .B(G137), .ZN(n406) );
  INV_X1 U458 ( .A(n406), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n395) );
  INV_X1 U460 ( .A(G101), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n391), .B(G110), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  INV_X1 U464 ( .A(n350), .ZN(n590) );
  XOR2_X1 U465 ( .A(KEYINPUT24), .B(G110), .Z(n399) );
  XNOR2_X1 U466 ( .A(n349), .B(G119), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n402) );
  XOR2_X1 U468 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n401) );
  XNOR2_X1 U469 ( .A(KEYINPUT91), .B(KEYINPUT78), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n402), .B(n355), .ZN(n405) );
  NAND2_X1 U471 ( .A1(G234), .A2(n745), .ZN(n403) );
  XOR2_X1 U472 ( .A(KEYINPUT8), .B(n403), .Z(n454) );
  NAND2_X1 U473 ( .A1(G221), .A2(n454), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U475 ( .A(n435), .B(KEYINPUT10), .ZN(n464) );
  XNOR2_X1 U476 ( .A(n464), .B(n406), .ZN(n742) );
  XNOR2_X1 U477 ( .A(n407), .B(n742), .ZN(n636) );
  NAND2_X1 U478 ( .A1(n636), .A2(n457), .ZN(n413) );
  XOR2_X1 U479 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n409) );
  XNOR2_X1 U480 ( .A(G902), .B(KEYINPUT15), .ZN(n627) );
  NAND2_X1 U481 ( .A1(G234), .A2(n627), .ZN(n408) );
  XNOR2_X1 U482 ( .A(n409), .B(n408), .ZN(n422) );
  NAND2_X1 U483 ( .A1(G217), .A2(n422), .ZN(n411) );
  INV_X1 U484 ( .A(KEYINPUT25), .ZN(n410) );
  XNOR2_X1 U485 ( .A(n411), .B(n410), .ZN(n412) );
  NAND2_X1 U486 ( .A1(G237), .A2(G234), .ZN(n414) );
  XNOR2_X1 U487 ( .A(n414), .B(KEYINPUT14), .ZN(n683) );
  NAND2_X1 U488 ( .A1(G902), .A2(n683), .ZN(n415) );
  NOR2_X1 U489 ( .A1(G900), .A2(n415), .ZN(n416) );
  NAND2_X1 U490 ( .A1(G953), .A2(n416), .ZN(n417) );
  XOR2_X1 U491 ( .A(KEYINPUT104), .B(n417), .Z(n420) );
  INV_X1 U492 ( .A(n683), .ZN(n418) );
  NAND2_X1 U493 ( .A1(n745), .A2(G952), .ZN(n504) );
  NOR2_X1 U494 ( .A1(n418), .A2(n504), .ZN(n419) );
  NOR2_X1 U495 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U496 ( .A(n421), .B(KEYINPUT75), .ZN(n425) );
  NAND2_X1 U497 ( .A1(G221), .A2(n422), .ZN(n424) );
  INV_X1 U498 ( .A(KEYINPUT21), .ZN(n423) );
  XNOR2_X1 U499 ( .A(n424), .B(n423), .ZN(n688) );
  NAND2_X1 U500 ( .A1(n425), .A2(n688), .ZN(n586) );
  INV_X1 U501 ( .A(n586), .ZN(n426) );
  AND2_X1 U502 ( .A1(n585), .A2(n426), .ZN(n427) );
  NAND2_X1 U503 ( .A1(n590), .A2(n427), .ZN(n428) );
  XNOR2_X1 U504 ( .A(n428), .B(KEYINPUT73), .ZN(n429) );
  NAND2_X1 U505 ( .A1(n745), .A2(G224), .ZN(n431) );
  XNOR2_X1 U506 ( .A(n431), .B(KEYINPUT74), .ZN(n432) );
  XNOR2_X1 U507 ( .A(n433), .B(n432), .ZN(n437) );
  XNOR2_X1 U508 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  XNOR2_X1 U509 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U510 ( .A(n437), .B(n436), .ZN(n443) );
  XNOR2_X2 U511 ( .A(G122), .B(G104), .ZN(n468) );
  XNOR2_X2 U512 ( .A(G116), .B(G107), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n468), .B(n451), .ZN(n440) );
  XNOR2_X1 U514 ( .A(KEYINPUT68), .B(KEYINPUT16), .ZN(n438) );
  INV_X1 U515 ( .A(G110), .ZN(n539) );
  XNOR2_X1 U516 ( .A(n438), .B(n539), .ZN(n439) );
  XNOR2_X1 U517 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U518 ( .A(n442), .B(n441), .ZN(n668) );
  INV_X1 U519 ( .A(n627), .ZN(n444) );
  XOR2_X1 U520 ( .A(KEYINPUT7), .B(KEYINPUT98), .Z(n447) );
  XNOR2_X1 U521 ( .A(G134), .B(G122), .ZN(n446) );
  XNOR2_X1 U522 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U523 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n448) );
  XNOR2_X1 U524 ( .A(n449), .B(n448), .ZN(n453) );
  XNOR2_X1 U525 ( .A(n450), .B(n451), .ZN(n452) );
  XNOR2_X1 U526 ( .A(n453), .B(n452), .ZN(n456) );
  NAND2_X1 U527 ( .A1(n454), .A2(G217), .ZN(n455) );
  XNOR2_X1 U528 ( .A(n456), .B(n455), .ZN(n632) );
  NAND2_X1 U529 ( .A1(n632), .A2(n457), .ZN(n459) );
  XOR2_X1 U530 ( .A(KEYINPUT100), .B(G478), .Z(n458) );
  XNOR2_X1 U531 ( .A(n459), .B(n458), .ZN(n509) );
  INV_X1 U532 ( .A(n509), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT13), .B(G475), .ZN(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n462) );
  NAND2_X1 U535 ( .A1(G214), .A2(n460), .ZN(n461) );
  XNOR2_X1 U536 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U537 ( .A(n463), .B(KEYINPUT97), .Z(n465) );
  XNOR2_X1 U538 ( .A(n465), .B(n464), .ZN(n471) );
  XOR2_X1 U539 ( .A(G140), .B(G143), .Z(n467) );
  XNOR2_X1 U540 ( .A(G113), .B(G131), .ZN(n466) );
  XNOR2_X1 U541 ( .A(n467), .B(n466), .ZN(n469) );
  XOR2_X1 U542 ( .A(n469), .B(n468), .Z(n470) );
  XNOR2_X1 U543 ( .A(n471), .B(n470), .ZN(n647) );
  OR2_X1 U544 ( .A1(G902), .A2(n647), .ZN(n472) );
  XNOR2_X1 U545 ( .A(n473), .B(n472), .ZN(n508) );
  INV_X1 U546 ( .A(n508), .ZN(n501) );
  AND2_X1 U547 ( .A1(n474), .A2(n501), .ZN(n546) );
  INV_X1 U548 ( .A(n546), .ZN(n475) );
  NOR2_X1 U549 ( .A1(n480), .A2(n475), .ZN(n476) );
  NAND2_X1 U550 ( .A1(n498), .A2(n476), .ZN(n604) );
  XOR2_X1 U551 ( .A(G143), .B(KEYINPUT111), .Z(n477) );
  XNOR2_X1 U552 ( .A(n604), .B(n477), .ZN(G45) );
  NAND2_X1 U553 ( .A1(n509), .A2(n501), .ZN(n570) );
  NOR2_X1 U554 ( .A1(n586), .A2(n570), .ZN(n479) );
  XNOR2_X1 U555 ( .A(n522), .B(KEYINPUT6), .ZN(n551) );
  NOR2_X1 U556 ( .A1(n585), .A2(n551), .ZN(n478) );
  NAND2_X1 U557 ( .A1(n479), .A2(n478), .ZN(n491) );
  INV_X1 U558 ( .A(n490), .ZN(n481) );
  INV_X1 U559 ( .A(n502), .ZN(n484) );
  NOR2_X1 U560 ( .A1(n491), .A2(n484), .ZN(n486) );
  XNOR2_X1 U561 ( .A(KEYINPUT84), .B(KEYINPUT36), .ZN(n485) );
  XNOR2_X1 U562 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U563 ( .A(n487), .B(KEYINPUT1), .ZN(n516) );
  INV_X1 U564 ( .A(n685), .ZN(n549) );
  NAND2_X1 U565 ( .A1(n488), .A2(n549), .ZN(n602) );
  XOR2_X1 U566 ( .A(G125), .B(KEYINPUT37), .Z(n489) );
  XNOR2_X1 U567 ( .A(n602), .B(n489), .ZN(G27) );
  NOR2_X1 U568 ( .A1(n491), .A2(n490), .ZN(n492) );
  NAND2_X1 U569 ( .A1(n492), .A2(n685), .ZN(n495) );
  XOR2_X1 U570 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n493) );
  XNOR2_X1 U571 ( .A(n493), .B(KEYINPUT105), .ZN(n494) );
  XNOR2_X1 U572 ( .A(n495), .B(n494), .ZN(n496) );
  NAND2_X1 U573 ( .A1(n496), .A2(n480), .ZN(n620) );
  XNOR2_X1 U574 ( .A(n620), .B(G140), .ZN(G42) );
  XNOR2_X1 U575 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n497) );
  XNOR2_X1 U576 ( .A(n480), .B(n497), .ZN(n704) );
  NAND2_X1 U577 ( .A1(n498), .A2(n704), .ZN(n500) );
  XNOR2_X1 U578 ( .A(KEYINPUT81), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U579 ( .A(n500), .B(n499), .ZN(n533) );
  OR2_X1 U580 ( .A1(n509), .A2(n501), .ZN(n569) );
  OR2_X1 U581 ( .A1(n533), .A2(n569), .ZN(n619) );
  XNOR2_X1 U582 ( .A(n619), .B(G134), .ZN(G36) );
  NOR2_X1 U583 ( .A1(G898), .A2(n745), .ZN(n503) );
  XOR2_X1 U584 ( .A(KEYINPUT89), .B(n503), .Z(n667) );
  NAND2_X1 U585 ( .A1(n667), .A2(G902), .ZN(n505) );
  NAND2_X1 U586 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U587 ( .A1(n506), .A2(n683), .ZN(n507) );
  AND2_X1 U588 ( .A1(n509), .A2(n508), .ZN(n583) );
  NAND2_X1 U589 ( .A1(n583), .A2(n688), .ZN(n510) );
  XNOR2_X1 U590 ( .A(n510), .B(KEYINPUT101), .ZN(n511) );
  NAND2_X1 U591 ( .A1(n543), .A2(n511), .ZN(n512) );
  INV_X1 U592 ( .A(KEYINPUT102), .ZN(n513) );
  XNOR2_X1 U593 ( .A(n585), .B(n513), .ZN(n690) );
  INV_X1 U594 ( .A(n690), .ZN(n514) );
  AND2_X1 U595 ( .A1(n685), .A2(n514), .ZN(n515) );
  XNOR2_X1 U596 ( .A(n572), .B(G101), .ZN(G3) );
  INV_X1 U597 ( .A(n516), .ZN(n519) );
  NAND2_X1 U598 ( .A1(n517), .A2(n688), .ZN(n684) );
  INV_X1 U599 ( .A(n684), .ZN(n518) );
  NAND2_X1 U600 ( .A1(n519), .A2(n518), .ZN(n521) );
  INV_X1 U601 ( .A(KEYINPUT71), .ZN(n520) );
  XNOR2_X1 U602 ( .A(n521), .B(n520), .ZN(n540) );
  INV_X1 U603 ( .A(n540), .ZN(n523) );
  BUF_X1 U604 ( .A(n522), .Z(n695) );
  AND2_X1 U605 ( .A1(n523), .A2(n695), .ZN(n698) );
  NAND2_X1 U606 ( .A1(n543), .A2(n698), .ZN(n525) );
  XNOR2_X1 U607 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n524) );
  XNOR2_X1 U608 ( .A(n525), .B(n524), .ZN(n568) );
  INV_X1 U609 ( .A(n570), .ZN(n737) );
  NAND2_X1 U610 ( .A1(n568), .A2(n737), .ZN(n526) );
  XNOR2_X1 U611 ( .A(n526), .B(G113), .ZN(G15) );
  INV_X1 U612 ( .A(n569), .ZN(n733) );
  NAND2_X1 U613 ( .A1(n568), .A2(n733), .ZN(n528) );
  XOR2_X1 U614 ( .A(G116), .B(KEYINPUT113), .Z(n527) );
  XNOR2_X1 U615 ( .A(n528), .B(n527), .ZN(G18) );
  OR2_X1 U616 ( .A1(n350), .A2(n684), .ZN(n529) );
  NOR2_X1 U617 ( .A1(n695), .A2(n529), .ZN(n530) );
  NAND2_X1 U618 ( .A1(n543), .A2(n530), .ZN(n531) );
  XNOR2_X1 U619 ( .A(n531), .B(KEYINPUT95), .ZN(n729) );
  NAND2_X1 U620 ( .A1(n729), .A2(n737), .ZN(n532) );
  XNOR2_X1 U621 ( .A(n532), .B(G104), .ZN(G6) );
  INV_X1 U622 ( .A(n533), .ZN(n534) );
  NAND2_X1 U623 ( .A1(n534), .A2(n737), .ZN(n536) );
  INV_X1 U624 ( .A(KEYINPUT40), .ZN(n535) );
  XNOR2_X1 U625 ( .A(n536), .B(n535), .ZN(n594) );
  XOR2_X1 U626 ( .A(G131), .B(n594), .Z(G33) );
  NOR2_X1 U627 ( .A1(n695), .A2(n585), .ZN(n537) );
  NAND2_X1 U628 ( .A1(n552), .A2(n367), .ZN(n538) );
  OR2_X2 U629 ( .A1(n540), .A2(n551), .ZN(n542) );
  XNOR2_X1 U630 ( .A(KEYINPUT86), .B(KEYINPUT33), .ZN(n541) );
  XNOR2_X2 U631 ( .A(n542), .B(n541), .ZN(n712) );
  NAND2_X1 U632 ( .A1(n712), .A2(n543), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n545), .B(n544), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U635 ( .A(n558), .B(G122), .Z(G24) );
  AND2_X1 U636 ( .A1(n549), .A2(n690), .ZN(n550) );
  NAND2_X1 U637 ( .A1(n552), .A2(n368), .ZN(n554) );
  INV_X1 U638 ( .A(KEYINPUT32), .ZN(n553) );
  XOR2_X1 U639 ( .A(G119), .B(n555), .Z(G21) );
  INV_X1 U640 ( .A(n555), .ZN(n557) );
  NAND2_X1 U641 ( .A1(n557), .A2(n556), .ZN(n564) );
  INV_X1 U642 ( .A(n558), .ZN(n560) );
  INV_X1 U643 ( .A(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n561) );
  INV_X1 U645 ( .A(KEYINPUT65), .ZN(n562) );
  NAND2_X1 U646 ( .A1(n562), .A2(KEYINPUT44), .ZN(n563) );
  NAND2_X1 U647 ( .A1(n559), .A2(KEYINPUT65), .ZN(n565) );
  NAND2_X1 U648 ( .A1(n566), .A2(KEYINPUT44), .ZN(n567) );
  XNOR2_X1 U649 ( .A(n567), .B(KEYINPUT83), .ZN(n575) );
  OR2_X1 U650 ( .A1(n729), .A2(n568), .ZN(n571) );
  AND2_X1 U651 ( .A1(n570), .A2(n569), .ZN(n708) );
  XNOR2_X1 U652 ( .A(n708), .B(KEYINPUT77), .ZN(n610) );
  NAND2_X1 U653 ( .A1(n571), .A2(n610), .ZN(n573) );
  NAND2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X2 U655 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U656 ( .A(n576), .B(KEYINPUT82), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n578), .A2(n577), .ZN(n580) );
  INV_X1 U658 ( .A(KEYINPUT80), .ZN(n579) );
  XNOR2_X2 U659 ( .A(n580), .B(n358), .ZN(n679) );
  NOR2_X2 U660 ( .A1(n679), .A2(n627), .ZN(n582) );
  INV_X1 U661 ( .A(KEYINPUT79), .ZN(n581) );
  XNOR2_X1 U662 ( .A(n582), .B(n581), .ZN(n625) );
  INV_X1 U663 ( .A(n583), .ZN(n706) );
  NAND2_X1 U664 ( .A1(n704), .A2(n481), .ZN(n707) );
  NOR2_X1 U665 ( .A1(n706), .A2(n707), .ZN(n584) );
  XNOR2_X1 U666 ( .A(KEYINPUT41), .B(n584), .ZN(n720) );
  NOR2_X1 U667 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n695), .A2(n587), .ZN(n588) );
  XNOR2_X1 U669 ( .A(KEYINPUT107), .B(n588), .ZN(n589) );
  XNOR2_X1 U670 ( .A(KEYINPUT28), .B(n589), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n592) );
  XNOR2_X1 U673 ( .A(n593), .B(n592), .ZN(n753) );
  INV_X1 U674 ( .A(KEYINPUT64), .ZN(n595) );
  INV_X1 U675 ( .A(n597), .ZN(n600) );
  INV_X1 U676 ( .A(n598), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n608), .A2(KEYINPUT47), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n708), .A2(KEYINPUT47), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT76), .ZN(n606) );
  OR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n614) );
  INV_X1 U684 ( .A(n608), .ZN(n738) );
  INV_X1 U685 ( .A(KEYINPUT47), .ZN(n609) );
  AND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n738), .A2(n611), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT69), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n618) );
  INV_X1 U691 ( .A(KEYINPUT48), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n622) );
  AND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  INV_X1 U694 ( .A(n679), .ZN(n661) );
  INV_X1 U695 ( .A(n744), .ZN(n680) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n626) );
  NOR2_X1 U697 ( .A1(n680), .A2(n626), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n630) );
  NOR2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X2 U700 ( .A1(n630), .A2(n629), .ZN(n671) );
  NAND2_X1 U701 ( .A1(n671), .A2(G478), .ZN(n631) );
  XOR2_X1 U702 ( .A(n632), .B(n631), .Z(n634) );
  INV_X1 U703 ( .A(G952), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n633), .A2(G953), .ZN(n657) );
  INV_X1 U705 ( .A(n657), .ZN(n677) );
  NOR2_X1 U706 ( .A1(n634), .A2(n677), .ZN(G63) );
  NAND2_X1 U707 ( .A1(n671), .A2(G217), .ZN(n635) );
  XOR2_X1 U708 ( .A(n636), .B(n635), .Z(n637) );
  NOR2_X1 U709 ( .A1(n637), .A2(n677), .ZN(G66) );
  NAND2_X1 U710 ( .A1(n671), .A2(G472), .ZN(n641) );
  XOR2_X1 U711 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n638) );
  XNOR2_X1 U712 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n642), .A2(n657), .ZN(n644) );
  XOR2_X1 U714 ( .A(KEYINPUT109), .B(KEYINPUT63), .Z(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n671), .A2(G475), .ZN(n649) );
  XNOR2_X1 U717 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n645) );
  XOR2_X1 U718 ( .A(n645), .B(KEYINPUT59), .Z(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n650), .A2(n657), .ZN(n652) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G60) );
  NAND2_X1 U724 ( .A1(n671), .A2(G210), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n653), .B(n654), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n660) );
  INV_X1 U729 ( .A(KEYINPUT56), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G51) );
  NAND2_X1 U731 ( .A1(n661), .A2(n745), .ZN(n666) );
  NAND2_X1 U732 ( .A1(G224), .A2(G953), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(KEYINPUT124), .ZN(n663) );
  XNOR2_X1 U734 ( .A(KEYINPUT61), .B(n663), .ZN(n664) );
  NAND2_X1 U735 ( .A1(G898), .A2(n664), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n670), .B(n669), .ZN(G69) );
  NAND2_X1 U739 ( .A1(n671), .A2(G469), .ZN(n676) );
  XNOR2_X1 U740 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT58), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n672), .B(n674), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(G54) );
  BUF_X1 U745 ( .A(n679), .Z(n681) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U747 ( .A(n682), .B(KEYINPUT2), .ZN(n725) );
  NAND2_X1 U748 ( .A1(G952), .A2(n683), .ZN(n718) );
  NAND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n686), .B(KEYINPUT50), .ZN(n687) );
  XNOR2_X1 U751 ( .A(KEYINPUT115), .B(n687), .ZN(n694) );
  INV_X1 U752 ( .A(n688), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n691), .B(KEYINPUT114), .ZN(n692) );
  XNOR2_X1 U755 ( .A(KEYINPUT49), .B(n692), .ZN(n693) );
  NOR2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n697) );
  INV_X1 U757 ( .A(n695), .ZN(n696) );
  AND2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n699) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U760 ( .A(KEYINPUT117), .B(n700), .Z(n702) );
  XOR2_X1 U761 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n701) );
  XNOR2_X1 U762 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n720), .A2(n703), .ZN(n715) );
  NOR2_X1 U764 ( .A1(n704), .A2(n481), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT118), .ZN(n713) );
  INV_X1 U769 ( .A(n712), .ZN(n719) );
  NOR2_X1 U770 ( .A1(n713), .A2(n719), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n716), .B(KEYINPUT52), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U774 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U776 ( .A(KEYINPUT119), .B(n723), .Z(n724) );
  NAND2_X1 U777 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n726), .B(KEYINPUT120), .ZN(n727) );
  NOR2_X1 U779 ( .A1(n727), .A2(G953), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U781 ( .A1(n729), .A2(n733), .ZN(n731) );
  XOR2_X1 U782 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n730) );
  XNOR2_X1 U783 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(G107), .B(n732), .ZN(G9) );
  XOR2_X1 U785 ( .A(KEYINPUT29), .B(KEYINPUT110), .Z(n735) );
  NAND2_X1 U786 ( .A1(n738), .A2(n733), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n349), .B(n736), .ZN(G30) );
  NAND2_X1 U789 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(KEYINPUT112), .ZN(n740) );
  XNOR2_X1 U791 ( .A(G146), .B(n740), .ZN(G48) );
  XNOR2_X1 U792 ( .A(n741), .B(n742), .ZN(n748) );
  XNOR2_X1 U793 ( .A(n748), .B(KEYINPUT125), .ZN(n743) );
  XNOR2_X1 U794 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n747), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U797 ( .A(n748), .B(G227), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U799 ( .A1(G953), .A2(n750), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U801 ( .A(G137), .B(n753), .Z(G39) );
endmodule

