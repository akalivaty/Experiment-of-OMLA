//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n447, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n594,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n652, new_n653, new_n656, new_n658, new_n659, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  AND2_X1   g052(.A1(new_n464), .A2(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n467), .B2(new_n474), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(G124), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n464), .A2(new_n466), .A3(new_n474), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT67), .A4(new_n474), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(G136), .A3(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n482), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n478), .A2(KEYINPUT4), .A3(G138), .A4(new_n474), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n474), .B2(G114), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n504), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n496), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(new_n511), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT71), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n520), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  AOI211_X1 g106(.A(new_n531), .B(new_n512), .C1(new_n514), .C2(new_n516), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n514), .A2(new_n516), .ZN(new_n533));
  INV_X1    g108(.A(new_n512), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT73), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(G63), .B(G651), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT6), .B1(KEYINPUT71), .B2(G651), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT74), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n524), .A2(new_n540), .A3(new_n525), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n541), .A3(G543), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(KEYINPUT75), .A2(G89), .ZN(new_n546));
  NOR2_X1   g121(.A1(KEYINPUT75), .A2(G89), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n533), .A2(new_n526), .A3(new_n534), .A4(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n550), .B1(new_n549), .B2(new_n552), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n536), .B(new_n545), .C1(new_n554), .C2(new_n555), .ZN(G286));
  INV_X1    g131(.A(G286), .ZN(G168));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n539), .A2(new_n541), .A3(G52), .A4(G543), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n533), .A2(new_n526), .A3(G90), .A4(new_n534), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n558), .A3(new_n560), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G64), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n515), .B1(new_n511), .B2(G543), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n513), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n534), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(new_n531), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n565), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G77), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n564), .A2(new_n574), .ZN(G301));
  INV_X1    g150(.A(G301), .ZN(G171));
  OAI21_X1  g151(.A(G56), .B1(new_n532), .B2(new_n535), .ZN(new_n577));
  NAND2_X1  g152(.A1(G68), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n519), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n517), .A2(new_n526), .ZN(new_n580));
  INV_X1    g155(.A(G81), .ZN(new_n581));
  INV_X1    g156(.A(G43), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n580), .A2(new_n581), .B1(new_n542), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT78), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G56), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n569), .B2(new_n570), .ZN(new_n586));
  INV_X1    g161(.A(new_n578), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  INV_X1    g164(.A(new_n583), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G860), .ZN(G153));
  AND3_X1   g168(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G36), .ZN(G176));
  NAND2_X1  g170(.A1(G1), .A2(G3), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT8), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT79), .ZN(G188));
  AND3_X1   g174(.A1(new_n539), .A2(new_n541), .A3(G543), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT9), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(G53), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G78), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G65), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n568), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  INV_X1    g182(.A(new_n580), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G91), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n539), .A2(new_n541), .A3(G53), .A4(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(KEYINPUT80), .B2(new_n601), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n603), .A2(new_n607), .A3(new_n609), .A4(new_n611), .ZN(G299));
  AOI22_X1  g187(.A1(new_n608), .A2(G87), .B1(new_n600), .B2(G49), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n569), .A2(new_n570), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G74), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n519), .ZN(G288));
  AND3_X1   g191(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n617));
  NAND2_X1  g192(.A1(G73), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G61), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n568), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n620), .B2(G651), .ZN(new_n621));
  INV_X1    g196(.A(G86), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n580), .ZN(G305));
  INV_X1    g198(.A(G60), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n569), .B2(new_n570), .ZN(new_n625));
  NAND2_X1  g200(.A1(G72), .A2(G543), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT81), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(G60), .B1(new_n532), .B2(new_n535), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(new_n630), .A3(new_n626), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n628), .A2(G651), .A3(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G85), .ZN(new_n633));
  INV_X1    g208(.A(G47), .ZN(new_n634));
  OAI22_X1  g209(.A1(new_n580), .A2(new_n633), .B1(new_n542), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n636), .ZN(G290));
  NAND2_X1  g212(.A1(G301), .A2(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(G79), .A2(G543), .ZN(new_n639));
  INV_X1    g214(.A(G66), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n568), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n641), .A2(G651), .B1(new_n600), .B2(G54), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n643));
  INV_X1    g218(.A(G92), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n580), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .A4(new_n526), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n638), .B1(G868), .B2(new_n649), .ZN(G284));
  OAI21_X1  g225(.A(new_n638), .B1(G868), .B2(new_n649), .ZN(G321));
  NAND2_X1  g226(.A1(G286), .A2(G868), .ZN(new_n652));
  INV_X1    g227(.A(G299), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(G868), .ZN(G297));
  OAI21_X1  g229(.A(new_n652), .B1(new_n653), .B2(G868), .ZN(G280));
  INV_X1    g230(.A(G559), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n649), .B1(new_n656), .B2(G860), .ZN(G148));
  NAND2_X1  g232(.A1(new_n649), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G868), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n592), .B2(G868), .ZN(G323));
  XNOR2_X1  g235(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g236(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT12), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT13), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2100), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n480), .A2(G123), .A3(new_n481), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n485), .A2(G135), .A3(new_n486), .ZN(new_n667));
  OR2_X1    g242(.A1(G99), .A2(G2105), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n668), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n671), .ZN(G156));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT83), .B(G2438), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2427), .B(G2430), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT14), .ZN(new_n678));
  XOR2_X1   g253(.A(G2451), .B(G2454), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1341), .B(G1348), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2443), .B(G2446), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G14), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G401));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  XOR2_X1   g264(.A(G2084), .B(G2090), .Z(new_n690));
  XNOR2_X1  g265(.A(G2067), .B(G2678), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n692), .B2(KEYINPUT18), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2096), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2100), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(KEYINPUT17), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  AOI21_X1  g272(.A(KEYINPUT18), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G227));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G1981), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT85), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT19), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1961), .B(G1966), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT86), .ZN(new_n708));
  XOR2_X1   g283(.A(G1956), .B(G2474), .Z(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n711), .A2(new_n712), .B1(new_n706), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n706), .A2(KEYINPUT20), .A3(new_n710), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n706), .A2(new_n710), .A3(new_n713), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G1986), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1991), .B(G1996), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(new_n718), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n702), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n726), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n728), .A2(new_n701), .A3(new_n724), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(G229));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G27), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G164), .B2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G2078), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n731), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2090), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n480), .A2(new_n481), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G128), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n485), .A2(new_n486), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G140), .ZN(new_n742));
  NOR2_X1   g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT90), .Z(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT91), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n731), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(G2067), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(G2067), .B1(new_n748), .B2(new_n751), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n734), .B(new_n738), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G32), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT26), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n480), .A2(G129), .A3(new_n481), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n485), .A2(G141), .A3(new_n486), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n765), .B(new_n766), .Z(new_n767));
  OR2_X1    g342(.A1(new_n733), .A2(G2078), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n649), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G4), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1348), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .C1(new_n737), .C2(G2090), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n755), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n774));
  NOR2_X1   g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT24), .A2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(G29), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(G160), .A2(G29), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n774), .B2(new_n778), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT99), .Z(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n592), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n787));
  INV_X1    g362(.A(G16), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n653), .B2(new_n788), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1956), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT31), .B(G11), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT98), .B1(G5), .B2(G16), .ZN(new_n795));
  OR3_X1    g370(.A1(KEYINPUT98), .A2(G5), .A3(G16), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n795), .B(new_n796), .C1(G301), .C2(new_n788), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1961), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n485), .A2(G139), .A3(new_n486), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT25), .Z(new_n801));
  NAND2_X1  g376(.A1(G115), .A2(G2104), .ZN(new_n802));
  INV_X1    g377(.A(G127), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n467), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n804), .A2(KEYINPUT93), .A3(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT93), .B1(new_n804), .B2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n799), .B(new_n801), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G33), .B(new_n807), .S(G29), .Z(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G2072), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n670), .A2(new_n731), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT97), .Z(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT30), .B(G28), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n731), .B2(new_n812), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n794), .A2(new_n798), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n773), .A2(new_n783), .A3(new_n793), .A4(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n770), .A2(new_n771), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  MUX2_X1   g393(.A(G6), .B(G305), .S(G16), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G16), .A2(G23), .ZN(new_n824));
  INV_X1    g399(.A(G288), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT33), .B(G1976), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n788), .A2(G22), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G166), .B2(new_n788), .ZN(new_n830));
  INV_X1    g405(.A(G1971), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n818), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n820), .B(new_n821), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n835), .A2(KEYINPUT34), .A3(new_n832), .A4(new_n828), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NAND2_X1  g413(.A1(G290), .A2(G16), .ZN(new_n839));
  INV_X1    g414(.A(G24), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT88), .B1(new_n840), .B2(G16), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n840), .A2(KEYINPUT88), .A3(G16), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n843), .A2(G1986), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(G1986), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n731), .A2(G25), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n739), .A2(G119), .ZN(new_n847));
  OR2_X1    g422(.A1(G95), .A2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT87), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n741), .A2(G131), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n846), .B1(new_n853), .B2(new_n731), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT35), .B(G1991), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n844), .A2(new_n845), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n837), .A2(new_n838), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n838), .B1(new_n837), .B2(new_n857), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n816), .B(new_n817), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n780), .A2(new_n781), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n788), .A2(G21), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(G168), .B2(new_n788), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT96), .B(G1966), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(G311));
  INV_X1    g442(.A(new_n859), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n837), .A2(new_n838), .A3(new_n857), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n815), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n861), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n865), .A4(new_n817), .ZN(G150));
  NAND2_X1  g447(.A1(new_n608), .A2(G93), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT102), .B(G55), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n600), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n614), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n519), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(G860), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT37), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n649), .A2(G559), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT39), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n873), .A2(new_n875), .ZN(new_n885));
  OAI21_X1  g460(.A(G67), .B1(new_n532), .B2(new_n535), .ZN(new_n886));
  INV_X1    g461(.A(G80), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n887), .B2(new_n513), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(G651), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n584), .B2(new_n591), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n579), .A2(new_n583), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n877), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n884), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n880), .B1(new_n894), .B2(new_n878), .ZN(G145));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n492), .A2(KEYINPUT104), .A3(new_n495), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT104), .B1(new_n492), .B2(new_n495), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n505), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT105), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(new_n505), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n746), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n739), .A2(G130), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n741), .A2(G142), .ZN(new_n906));
  OR2_X1    g481(.A1(G106), .A2(G2105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(G2104), .C1(G118), .C2(new_n474), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n900), .A2(new_n746), .A3(new_n902), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n900), .A2(new_n746), .A3(new_n902), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(new_n903), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n896), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n914), .A3(new_n896), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G160), .A2(new_n670), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n476), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n490), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(G162), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n763), .A2(new_n807), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n763), .B1(new_n924), .B2(new_n807), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n922), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n807), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n764), .B1(new_n929), .B2(KEYINPUT106), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n919), .A2(G162), .A3(new_n920), .ZN(new_n931));
  AOI21_X1  g506(.A(G162), .B1(new_n919), .B2(new_n920), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n930), .B(new_n925), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n933), .A3(new_n852), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n663), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n852), .B1(new_n928), .B2(new_n933), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n853), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n663), .B1(new_n940), .B2(new_n934), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n918), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n663), .A3(new_n934), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n916), .A4(new_n917), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT108), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g524(.A(new_n893), .B(new_n658), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n648), .A2(G299), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n610), .B(new_n602), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n606), .A2(G651), .B1(new_n608), .B2(G91), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n642), .A4(new_n647), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n951), .A2(KEYINPUT41), .A3(new_n954), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT41), .B1(new_n951), .B2(new_n954), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(new_n950), .ZN(new_n960));
  XNOR2_X1  g535(.A(G303), .B(G305), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n632), .A2(new_n636), .A3(G288), .ZN(new_n962));
  AOI21_X1  g537(.A(G288), .B1(new_n632), .B2(new_n636), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n962), .A2(new_n963), .A3(KEYINPUT109), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(new_n825), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n632), .A2(new_n636), .A3(G288), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n965), .A3(new_n967), .ZN(new_n971));
  INV_X1    g546(.A(new_n961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT42), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(KEYINPUT42), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n970), .A2(KEYINPUT42), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT109), .B1(new_n962), .B2(new_n963), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n977), .B2(new_n971), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n962), .A2(new_n963), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n961), .B1(new_n979), .B2(new_n965), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n975), .B(new_n976), .C1(new_n978), .C2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n960), .A2(new_n974), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n960), .B1(new_n974), .B2(new_n981), .ZN(new_n983));
  OAI21_X1  g558(.A(G868), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(G868), .B2(new_n889), .ZN(G295));
  OAI21_X1  g560(.A(new_n984), .B1(G868), .B2(new_n889), .ZN(G331));
  NAND2_X1  g561(.A1(new_n549), .A2(new_n552), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT76), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n544), .B1(new_n988), .B2(new_n553), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n559), .A2(new_n558), .A3(new_n560), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n561), .ZN(new_n991));
  OAI21_X1  g566(.A(G64), .B1(new_n532), .B2(new_n535), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n519), .B1(new_n992), .B2(new_n572), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n989), .B(new_n536), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(G286), .A2(new_n564), .A3(new_n574), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n583), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n877), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n889), .B1(new_n579), .B2(new_n583), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n994), .A2(new_n995), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n890), .B2(new_n892), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n959), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(new_n1003), .A3(new_n955), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n969), .A3(new_n973), .A4(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1001), .A2(new_n955), .A3(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n959), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1010));
  OAI22_X1  g585(.A1(new_n1009), .A2(new_n1010), .B1(new_n978), .B2(new_n980), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1011), .A3(new_n946), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1008), .A2(new_n1011), .A3(new_n1014), .A4(new_n946), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(KEYINPUT44), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1017), .A3(new_n1015), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1020), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g596(.A(new_n746), .B(G2067), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n763), .B(G1996), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n852), .A2(new_n855), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n852), .A2(new_n855), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G290), .A2(G1986), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G290), .A2(G1986), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n900), .A2(new_n902), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n900), .B2(new_n902), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n470), .A2(new_n475), .A3(G40), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1033), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1039), .B2(KEYINPUT45), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G164), .A2(G1384), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT113), .B1(new_n1048), .B2(KEYINPUT45), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(new_n1038), .C1(G164), .C2(G1384), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(KEYINPUT118), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n899), .A2(new_n1035), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT50), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n508), .B(new_n506), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1054), .B(new_n1035), .C1(new_n1058), .C2(new_n496), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1055), .A2(new_n1057), .A3(new_n1061), .A4(new_n1043), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(G2090), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1053), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT114), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n1067));
  NAND4_X1  g642(.A1(G303), .A2(new_n1067), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(G166), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1066), .A2(KEYINPUT115), .A3(new_n1068), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1064), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n899), .A2(new_n1035), .A3(new_n1043), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(G8), .C1(new_n1080), .C2(G288), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(G1976), .B2(new_n825), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G305), .A2(G1981), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  INV_X1    g660(.A(G1981), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT117), .B(G86), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n608), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n621), .B2(new_n1088), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n1084), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1079), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1073), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1085), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1081), .A2(new_n1095), .A3(KEYINPUT52), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1081), .B2(KEYINPUT52), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1083), .B(new_n1094), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n899), .A2(new_n1054), .A3(new_n1035), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n1043), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(G2090), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1076), .B(G8), .C1(new_n1053), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1966), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT45), .B(new_n1035), .C1(new_n1058), .C2(new_n496), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1043), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT45), .B1(new_n899), .B2(new_n1035), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1100), .A2(new_n1101), .A3(new_n781), .A4(new_n1043), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(G168), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G8), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT51), .ZN(new_n1113));
  AOI21_X1  g688(.A(G168), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  OAI211_X1 g690(.A(G8), .B(new_n1111), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AND4_X1   g692(.A1(new_n1078), .A2(new_n1099), .A3(new_n1104), .A4(new_n1117), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1119));
  INV_X1    g694(.A(G2078), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1042), .A2(KEYINPUT53), .A3(new_n1120), .A4(new_n1047), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1039), .A2(KEYINPUT45), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1122), .A2(new_n1052), .A3(new_n1120), .A4(new_n1043), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g699(.A(G1961), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1123), .A2(new_n1124), .B1(new_n1125), .B2(new_n1102), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1121), .A2(new_n1126), .A3(G301), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1107), .A2(new_n1108), .A3(G2078), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1128), .A2(KEYINPUT123), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(KEYINPUT123), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT53), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(G301), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1119), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(new_n1131), .A3(G301), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT54), .B(new_n1134), .C1(new_n1135), .C2(G301), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1118), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1047), .A2(new_n1052), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1956), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1062), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G299), .B(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1139), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT61), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(KEYINPUT120), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n648), .A2(KEYINPUT121), .ZN(new_n1153));
  INV_X1    g728(.A(G2067), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1102), .A2(new_n771), .B1(new_n1091), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1155), .B2(KEYINPUT60), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(KEYINPUT60), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n648), .B(KEYINPUT121), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1996), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1047), .A2(new_n1161), .A3(new_n1052), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT58), .B(G1341), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1091), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n592), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1164), .A2(new_n1167), .A3(new_n592), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1150), .A2(new_n1152), .A3(new_n1160), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1144), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1155), .A2(new_n648), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1147), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT119), .Z(new_n1174));
  AOI21_X1  g749(.A(new_n1137), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1112), .A2(G286), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1078), .A2(new_n1099), .A3(new_n1104), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(G8), .B1(new_n1053), .B2(new_n1103), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1180), .B2(new_n1077), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1181), .A2(new_n1104), .A3(new_n1099), .A4(new_n1176), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT124), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1078), .A2(new_n1099), .A3(new_n1104), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1113), .A2(new_n1116), .A3(new_n1184), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1132), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1185), .A2(KEYINPUT124), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1104), .A2(new_n1098), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1094), .A2(new_n1080), .A3(new_n825), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1193), .B1(G1981), .B2(G305), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1092), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1183), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1046), .B1(new_n1175), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1045), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1026), .B1(new_n1198), .B2(new_n1024), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n746), .A2(G2067), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1199), .A2(KEYINPUT125), .A3(new_n1200), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1203), .A2(new_n1045), .A3(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1198), .A2(new_n1032), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1206), .A2(KEYINPUT48), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(KEYINPUT48), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1207), .B(new_n1208), .C1(new_n1198), .C2(new_n1029), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1045), .A2(new_n1161), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1211));
  OR2_X1    g786(.A1(new_n1211), .A2(KEYINPUT46), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1210), .B(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT47), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1022), .A2(new_n763), .ZN(new_n1215));
  AOI22_X1  g790(.A1(new_n1045), .A2(new_n1215), .B1(new_n1211), .B2(KEYINPUT46), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1214), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1205), .B(new_n1209), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1197), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g796(.A1(new_n727), .A2(new_n729), .A3(new_n699), .ZN(new_n1223));
  NAND4_X1  g797(.A1(new_n947), .A2(new_n1223), .A3(G319), .A4(new_n687), .ZN(new_n1224));
  OAI21_X1  g798(.A(KEYINPUT127), .B1(new_n1020), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g799(.A(new_n1224), .ZN(new_n1226));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  NAND4_X1  g801(.A1(new_n1226), .A2(new_n1227), .A3(new_n1019), .A4(new_n1018), .ZN(new_n1228));
  AND2_X1   g802(.A1(new_n1225), .A2(new_n1228), .ZN(G308));
  NAND2_X1  g803(.A1(new_n1225), .A2(new_n1228), .ZN(G225));
endmodule


