

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n544), .A2(n543), .ZN(G164) );
  AND2_X1 U551 ( .A1(n715), .A2(G2072), .ZN(n703) );
  NOR2_X1 U552 ( .A1(n977), .A2(n693), .ZN(n695) );
  INV_X1 U553 ( .A(KEYINPUT28), .ZN(n710) );
  INV_X1 U554 ( .A(KEYINPUT97), .ZN(n730) );
  NOR2_X1 U555 ( .A1(G1384), .A2(G164), .ZN(n689) );
  INV_X1 U556 ( .A(G2104), .ZN(n522) );
  NOR2_X2 U557 ( .A1(G2105), .A2(n522), .ZN(n893) );
  NOR2_X1 U558 ( .A1(n638), .A2(G651), .ZN(n648) );
  NOR2_X1 U559 ( .A1(n527), .A2(n526), .ZN(G160) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X1 U561 ( .A(KEYINPUT17), .B(n517), .Z(n518) );
  XNOR2_X1 U562 ( .A(KEYINPUT66), .B(n518), .ZN(n608) );
  NAND2_X1 U563 ( .A1(G137), .A2(n608), .ZN(n521) );
  NAND2_X1 U564 ( .A1(G101), .A2(n893), .ZN(n519) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n519), .Z(n520) );
  NAND2_X1 U566 ( .A1(n521), .A2(n520), .ZN(n527) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U568 ( .A1(G113), .A2(n887), .ZN(n525) );
  NAND2_X1 U569 ( .A1(n522), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U570 ( .A(n523), .B(KEYINPUT65), .ZN(n889) );
  NAND2_X1 U571 ( .A1(G125), .A2(n889), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n526) );
  INV_X1 U573 ( .A(G96), .ZN(G221) );
  XOR2_X1 U574 ( .A(G2427), .B(G2435), .Z(n529) );
  XNOR2_X1 U575 ( .A(G2454), .B(G2443), .ZN(n528) );
  XNOR2_X1 U576 ( .A(n529), .B(n528), .ZN(n536) );
  XOR2_X1 U577 ( .A(G2451), .B(KEYINPUT103), .Z(n531) );
  XNOR2_X1 U578 ( .A(G2430), .B(G2438), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U580 ( .A(n532), .B(G2446), .Z(n534) );
  XNOR2_X1 U581 ( .A(G1348), .B(G1341), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U583 ( .A(n536), .B(n535), .ZN(n537) );
  AND2_X1 U584 ( .A1(n537), .A2(G14), .ZN(G401) );
  AND2_X1 U585 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U586 ( .A1(G114), .A2(n887), .ZN(n538) );
  XNOR2_X1 U587 ( .A(n538), .B(KEYINPUT88), .ZN(n540) );
  NAND2_X1 U588 ( .A1(G138), .A2(n608), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U590 ( .A1(G102), .A2(n893), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G126), .A2(n889), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  INV_X1 U594 ( .A(G651), .ZN(n551) );
  NOR2_X1 U595 ( .A1(n638), .A2(n551), .ZN(n655) );
  NAND2_X1 U596 ( .A1(n655), .A2(G76), .ZN(n545) );
  XNOR2_X1 U597 ( .A(KEYINPUT74), .B(n545), .ZN(n548) );
  NOR2_X1 U598 ( .A1(G543), .A2(G651), .ZN(n651) );
  NAND2_X1 U599 ( .A1(n651), .A2(G89), .ZN(n546) );
  XNOR2_X1 U600 ( .A(KEYINPUT4), .B(n546), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U602 ( .A(n549), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U603 ( .A1(n648), .A2(G51), .ZN(n550) );
  XOR2_X1 U604 ( .A(KEYINPUT75), .B(n550), .Z(n554) );
  NOR2_X1 U605 ( .A1(G543), .A2(n551), .ZN(n552) );
  XOR2_X1 U606 ( .A(KEYINPUT1), .B(n552), .Z(n647) );
  NAND2_X1 U607 ( .A1(n647), .A2(G63), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U611 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U614 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U615 ( .A(G223), .B(KEYINPUT72), .Z(n834) );
  NAND2_X1 U616 ( .A1(n834), .A2(G567), .ZN(n560) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U618 ( .A1(n651), .A2(G81), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G68), .A2(n655), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT13), .B(n564), .Z(n568) );
  NAND2_X1 U623 ( .A1(G56), .A2(n647), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT73), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT14), .ZN(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n648), .A2(G43), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n977) );
  INV_X1 U629 ( .A(G860), .ZN(n599) );
  OR2_X1 U630 ( .A1(n977), .A2(n599), .ZN(G153) );
  NAND2_X1 U631 ( .A1(G64), .A2(n647), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G52), .A2(n648), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n651), .A2(G90), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n573), .B(KEYINPUT68), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G77), .A2(n655), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U640 ( .A(KEYINPUT69), .B(n579), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U642 ( .A1(G92), .A2(n651), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G79), .A2(n655), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G66), .A2(n647), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G54), .A2(n648), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U649 ( .A(KEYINPUT15), .B(n586), .Z(n976) );
  OR2_X1 U650 ( .A1(n976), .A2(G868), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G78), .A2(n655), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G65), .A2(n647), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U655 ( .A1(n651), .A2(G91), .ZN(n591) );
  XOR2_X1 U656 ( .A(KEYINPUT70), .B(n591), .Z(n592) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U658 ( .A1(n648), .A2(G53), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(G299) );
  INV_X1 U660 ( .A(G868), .ZN(n667) );
  NOR2_X1 U661 ( .A1(G286), .A2(n667), .ZN(n597) );
  NOR2_X1 U662 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U664 ( .A(KEYINPUT76), .B(n598), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n600), .A2(n976), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U668 ( .A1(n976), .A2(G868), .ZN(n602) );
  XOR2_X1 U669 ( .A(KEYINPUT77), .B(n602), .Z(n603) );
  NOR2_X1 U670 ( .A1(G559), .A2(n603), .ZN(n604) );
  XNOR2_X1 U671 ( .A(n604), .B(KEYINPUT78), .ZN(n606) );
  NOR2_X1 U672 ( .A1(n977), .A2(G868), .ZN(n605) );
  NOR2_X1 U673 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U674 ( .A1(n889), .A2(G123), .ZN(n607) );
  XNOR2_X1 U675 ( .A(n607), .B(KEYINPUT18), .ZN(n610) );
  BUF_X1 U676 ( .A(n608), .Z(n896) );
  NAND2_X1 U677 ( .A1(G135), .A2(n896), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G99), .A2(n893), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G111), .A2(n887), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(n613), .Z(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n926) );
  XNOR2_X1 U684 ( .A(n926), .B(G2096), .ZN(n616) );
  INV_X1 U685 ( .A(G2100), .ZN(n847) );
  NAND2_X1 U686 ( .A1(n616), .A2(n847), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G67), .A2(n647), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G55), .A2(n648), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G93), .A2(n651), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G80), .A2(n655), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(n621), .Z(n622) );
  NOR2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n666) );
  XNOR2_X1 U695 ( .A(KEYINPUT80), .B(n977), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n976), .A2(G559), .ZN(n664) );
  XNOR2_X1 U697 ( .A(n624), .B(n664), .ZN(n625) );
  NOR2_X1 U698 ( .A1(G860), .A2(n625), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n666), .B(n626), .ZN(G145) );
  NAND2_X1 U700 ( .A1(G73), .A2(n655), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT2), .ZN(n634) );
  NAND2_X1 U702 ( .A1(G61), .A2(n647), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G48), .A2(n648), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n651), .A2(G86), .ZN(n630) );
  XOR2_X1 U706 ( .A(KEYINPUT82), .B(n630), .Z(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U709 ( .A1(G49), .A2(n648), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n647), .A2(n637), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G88), .A2(n651), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G75), .A2(n655), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G62), .A2(n647), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G50), .A2(n648), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G60), .A2(n647), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G47), .A2(n648), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U725 ( .A1(G85), .A2(n651), .ZN(n652) );
  XNOR2_X1 U726 ( .A(KEYINPUT67), .B(n652), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n655), .A2(G72), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n657), .A2(n656), .ZN(G290) );
  XNOR2_X1 U730 ( .A(n666), .B(n977), .ZN(n663) );
  XNOR2_X1 U731 ( .A(G288), .B(KEYINPUT19), .ZN(n659) );
  XOR2_X1 U732 ( .A(G299), .B(G166), .Z(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U734 ( .A(n660), .B(G290), .Z(n661) );
  XNOR2_X1 U735 ( .A(G305), .B(n661), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n840) );
  XNOR2_X1 U737 ( .A(n664), .B(n840), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U741 ( .A(KEYINPUT83), .B(n670), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U749 ( .A1(G108), .A2(G120), .ZN(n675) );
  NOR2_X1 U750 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(G69), .A2(n676), .ZN(n838) );
  NAND2_X1 U752 ( .A1(G567), .A2(n838), .ZN(n677) );
  XOR2_X1 U753 ( .A(KEYINPUT86), .B(n677), .Z(n684) );
  NAND2_X1 U754 ( .A1(G132), .A2(G82), .ZN(n678) );
  XNOR2_X1 U755 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  XNOR2_X1 U756 ( .A(n679), .B(KEYINPUT84), .ZN(n680) );
  NOR2_X1 U757 ( .A1(G218), .A2(n680), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(KEYINPUT85), .ZN(n682) );
  OR2_X1 U759 ( .A1(G221), .A2(n682), .ZN(n839) );
  AND2_X1 U760 ( .A1(n839), .A2(G2106), .ZN(n683) );
  NOR2_X1 U761 ( .A1(n684), .A2(n683), .ZN(G319) );
  INV_X1 U762 ( .A(G319), .ZN(n917) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n917), .A2(n685), .ZN(n686) );
  XOR2_X1 U765 ( .A(KEYINPUT87), .B(n686), .Z(n837) );
  NAND2_X1 U766 ( .A1(n837), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U768 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n833) );
  INV_X1 U769 ( .A(KEYINPUT64), .ZN(n688) );
  XNOR2_X1 U770 ( .A(n689), .B(n688), .ZN(n782) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n781) );
  NOR2_X2 U772 ( .A1(n782), .A2(n781), .ZN(n715) );
  AND2_X1 U773 ( .A1(n715), .A2(G1996), .ZN(n690) );
  XOR2_X1 U774 ( .A(n690), .B(KEYINPUT26), .Z(n692) );
  INV_X1 U775 ( .A(n715), .ZN(n734) );
  NAND2_X1 U776 ( .A1(n734), .A2(G1341), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U778 ( .A1(n695), .A2(n976), .ZN(n694) );
  XNOR2_X1 U779 ( .A(n694), .B(KEYINPUT95), .ZN(n701) );
  NAND2_X1 U780 ( .A1(n695), .A2(n976), .ZN(n699) );
  NOR2_X1 U781 ( .A1(n715), .A2(G1348), .ZN(n697) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n734), .ZN(n696) );
  NOR2_X1 U783 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U785 ( .A1(n701), .A2(n700), .ZN(n708) );
  INV_X1 U786 ( .A(G299), .ZN(n986) );
  XNOR2_X1 U787 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n702) );
  XNOR2_X1 U788 ( .A(n703), .B(n702), .ZN(n705) );
  XOR2_X1 U789 ( .A(G1956), .B(KEYINPUT93), .Z(n947) );
  NAND2_X1 U790 ( .A1(n734), .A2(n947), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U792 ( .A(KEYINPUT94), .B(n706), .Z(n709) );
  NAND2_X1 U793 ( .A1(n986), .A2(n709), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U795 ( .A1(n986), .A2(n709), .ZN(n711) );
  XNOR2_X1 U796 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U797 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U798 ( .A(n714), .B(KEYINPUT29), .ZN(n719) );
  NAND2_X1 U799 ( .A1(G1961), .A2(n734), .ZN(n717) );
  XOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .Z(n1008) );
  NAND2_X1 U801 ( .A1(n715), .A2(n1008), .ZN(n716) );
  NAND2_X1 U802 ( .A1(n717), .A2(n716), .ZN(n720) );
  NOR2_X1 U803 ( .A1(G301), .A2(n720), .ZN(n718) );
  NOR2_X1 U804 ( .A1(n719), .A2(n718), .ZN(n729) );
  NAND2_X1 U805 ( .A1(G301), .A2(n720), .ZN(n721) );
  XOR2_X1 U806 ( .A(KEYINPUT96), .B(n721), .Z(n726) );
  NAND2_X1 U807 ( .A1(G8), .A2(n734), .ZN(n771) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n771), .ZN(n745) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n734), .ZN(n743) );
  NOR2_X1 U810 ( .A1(n745), .A2(n743), .ZN(n722) );
  NAND2_X1 U811 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U813 ( .A1(G168), .A2(n724), .ZN(n725) );
  NOR2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U815 ( .A(n727), .B(KEYINPUT31), .ZN(n728) );
  NOR2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U817 ( .A(n731), .B(n730), .ZN(n744) );
  INV_X1 U818 ( .A(n744), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n732), .A2(G286), .ZN(n741) );
  INV_X1 U820 ( .A(G8), .ZN(n739) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n771), .ZN(n733) );
  XNOR2_X1 U822 ( .A(n733), .B(KEYINPUT98), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n734), .A2(G2090), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n737), .A2(G303), .ZN(n738) );
  OR2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U828 ( .A(n742), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X1 U829 ( .A1(G8), .A2(n743), .ZN(n747) );
  NOR2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n763) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n985) );
  AND2_X1 U833 ( .A1(n763), .A2(n985), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n762), .A2(n748), .ZN(n752) );
  INV_X1 U835 ( .A(n985), .ZN(n750) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n758) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n758), .A2(n749), .ZN(n990) );
  OR2_X1 U839 ( .A1(n750), .A2(n990), .ZN(n751) );
  AND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n753), .A2(n771), .ZN(n754) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  NOR2_X1 U843 ( .A1(KEYINPUT99), .A2(n755), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(KEYINPUT33), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n775) );
  INV_X1 U846 ( .A(n771), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n758), .A2(KEYINPUT99), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n761), .A2(KEYINPUT33), .ZN(n768) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n766) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G8), .A2(n764), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n767), .A2(n771), .ZN(n776) );
  AND2_X1 U855 ( .A1(n768), .A2(n776), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U857 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n779) );
  INV_X1 U859 ( .A(n779), .ZN(n772) );
  AND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n817) );
  INV_X1 U862 ( .A(n776), .ZN(n778) );
  XOR2_X1 U863 ( .A(G1981), .B(KEYINPUT100), .Z(n777) );
  XNOR2_X1 U864 ( .A(G305), .B(n777), .ZN(n972) );
  OR2_X1 U865 ( .A1(n778), .A2(n972), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n815) );
  XNOR2_X1 U867 ( .A(G1986), .B(G290), .ZN(n992) );
  INV_X1 U868 ( .A(n781), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n810) );
  INV_X1 U870 ( .A(n810), .ZN(n828) );
  AND2_X1 U871 ( .A1(n992), .A2(n828), .ZN(n813) );
  NAND2_X1 U872 ( .A1(G104), .A2(n893), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G140), .A2(n896), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT34), .B(n786), .ZN(n792) );
  NAND2_X1 U876 ( .A1(n887), .A2(G116), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT89), .B(n787), .Z(n789) );
  NAND2_X1 U878 ( .A1(n889), .A2(G128), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U880 ( .A(n790), .B(KEYINPUT35), .Z(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U882 ( .A(KEYINPUT36), .B(n793), .Z(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT90), .B(n794), .Z(n913) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U885 ( .A1(n913), .A2(n826), .ZN(n942) );
  NAND2_X1 U886 ( .A1(n828), .A2(n942), .ZN(n824) );
  NAND2_X1 U887 ( .A1(G95), .A2(n893), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G131), .A2(n896), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G107), .A2(n887), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G119), .A2(n889), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n909) );
  XNOR2_X1 U894 ( .A(KEYINPUT91), .B(G1991), .ZN(n1005) );
  NOR2_X1 U895 ( .A1(n909), .A2(n1005), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n889), .A2(G129), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G141), .A2(n896), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n893), .A2(G105), .ZN(n803) );
  XOR2_X1 U900 ( .A(KEYINPUT38), .B(n803), .Z(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n887), .A2(G117), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n885) );
  AND2_X1 U904 ( .A1(G1996), .A2(n885), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n928) );
  NOR2_X1 U906 ( .A1(n928), .A2(n810), .ZN(n821) );
  INV_X1 U907 ( .A(n821), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n824), .A2(n811), .ZN(n812) );
  OR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n831) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n885), .ZN(n923) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n1005), .A2(n909), .ZN(n818) );
  XNOR2_X1 U915 ( .A(n818), .B(KEYINPUT101), .ZN(n930) );
  NOR2_X1 U916 ( .A1(n819), .A2(n930), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n923), .A2(n822), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n913), .A2(n826), .ZN(n931) );
  NAND2_X1 U922 ( .A1(n827), .A2(n931), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G82), .ZN(G220) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n842) );
  XNOR2_X1 U940 ( .A(n976), .B(n840), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U942 ( .A(G286), .B(G301), .Z(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  NOR2_X1 U944 ( .A1(G37), .A2(n845), .ZN(n846) );
  XOR2_X1 U945 ( .A(KEYINPUT117), .B(n846), .Z(G397) );
  XNOR2_X1 U946 ( .A(n847), .B(G2096), .ZN(n849) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1966), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n858), .B(KEYINPUT104), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1971), .B(G1976), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(G1981), .B(G1956), .Z(n862) );
  XNOR2_X1 U962 ( .A(G1986), .B(G1961), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U965 ( .A(KEYINPUT105), .B(G2474), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U967 ( .A1(n896), .A2(G136), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n867), .B(KEYINPUT106), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G100), .A2(n893), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT108), .B(n868), .Z(n871) );
  NAND2_X1 U971 ( .A1(n889), .A2(G124), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT44), .B(n869), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G112), .A2(n887), .ZN(n874) );
  XNOR2_X1 U976 ( .A(KEYINPUT107), .B(n874), .ZN(n875) );
  NOR2_X1 U977 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G106), .A2(n893), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G142), .A2(n896), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT45), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G118), .A2(n887), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G130), .A2(n889), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U985 ( .A(KEYINPUT109), .B(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n902) );
  NAND2_X1 U988 ( .A1(n887), .A2(G115), .ZN(n888) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n888), .Z(n891) );
  NAND2_X1 U990 ( .A1(n889), .A2(G127), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n892), .B(KEYINPUT47), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n899) );
  NAND2_X1 U995 ( .A1(n896), .A2(G139), .ZN(n897) );
  XOR2_X1 U996 ( .A(KEYINPUT110), .B(n897), .Z(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(n900), .Z(n933) );
  XOR2_X1 U999 ( .A(G164), .B(n933), .Z(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(G160), .B(G162), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n903), .B(n926), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n905), .B(n904), .Z(n911) );
  XOR2_X1 U1004 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n916), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(n917), .A2(G401), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT118), .B(n918), .Z(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(n919), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n924), .Z(n940) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n935) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n933), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n936), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1035 ( .A(KEYINPUT52), .B(n943), .Z(n944) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(KEYINPUT119), .B(n945), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n946), .A2(G29), .ZN(n1001) );
  XOR2_X1 U1039 ( .A(G1981), .B(G6), .Z(n949) );
  XOR2_X1 U1040 ( .A(n947), .B(G20), .Z(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G19), .B(G1341), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1044 ( .A(KEYINPUT126), .B(n952), .Z(n956) );
  XNOR2_X1 U1045 ( .A(KEYINPUT59), .B(KEYINPUT127), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(n953), .B(G4), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G1348), .B(n954), .ZN(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n957), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(G1961), .B(G5), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT61), .B(n969), .Z(n970) );
  NOR2_X1 U1062 ( .A1(G16), .A2(n970), .ZN(n999) );
  XNOR2_X1 U1063 ( .A(KEYINPUT56), .B(G16), .ZN(n996) );
  XOR2_X1 U1064 ( .A(G1966), .B(G168), .Z(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT123), .B(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n975), .B(n974), .ZN(n981) );
  XOR2_X1 U1069 ( .A(G1348), .B(n976), .Z(n979) );
  XNOR2_X1 U1070 ( .A(n977), .B(G1341), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1073 ( .A(G1961), .B(G171), .Z(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n994) );
  NAND2_X1 U1075 ( .A1(G1971), .A2(G303), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G1956), .B(n986), .Z(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(KEYINPUT125), .B(n997), .ZN(n998) );
  NOR2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1085 ( .A1(n1001), .A2(n1000), .ZN(n1027) );
  XOR2_X1 U1086 ( .A(G2090), .B(G35), .Z(n1018) );
  XNOR2_X1 U1087 ( .A(G2067), .B(G26), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(G2072), .B(G33), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(n1004), .B(KEYINPUT120), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(n1005), .B(G25), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XNOR2_X1 U1093 ( .A(G1996), .B(G32), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(n1008), .B(G27), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(n1011), .B(KEYINPUT121), .ZN(n1012) );
  NOR2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(G28), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1015), .B(KEYINPUT53), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(n1016), .B(KEYINPUT122), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(G34), .B(G2084), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(KEYINPUT54), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(KEYINPUT55), .B(n1022), .ZN(n1024) );
  INV_X1 U1106 ( .A(G29), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(G11), .ZN(n1026) );
  NOR2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(n1028), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

