//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915;
  NOR2_X1   g000(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n204));
  OR3_X1    g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(new_n207), .A3(new_n209), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n204), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n204), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT17), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n219), .B(new_n220), .C1(G1gat), .C2(new_n217), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n215), .A2(KEYINPUT17), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n216), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n215), .A2(new_n223), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n203), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(new_n228), .A3(new_n226), .A4(new_n203), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n215), .B(new_n223), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n228), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235));
  INV_X1    g034(.A(G197gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT11), .B(G169gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT12), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OR3_X1    g040(.A1(new_n229), .A2(new_n234), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n229), .B2(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G15gat), .B(G43gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(new_n247), .Z(new_n248));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n251), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n252), .A2(KEYINPUT68), .B1(new_n253), .B2(KEYINPUT67), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT68), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n256));
  OAI22_X1  g055(.A1(new_n255), .A2(new_n256), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(KEYINPUT23), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(KEYINPUT23), .ZN(new_n262));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n261), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT25), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n269));
  INV_X1    g068(.A(G183gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n272));
  AOI21_X1  g071(.A(G190gat), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n268), .B1(new_n273), .B2(KEYINPUT69), .ZN(new_n274));
  INV_X1    g073(.A(new_n268), .ZN(new_n275));
  INV_X1    g074(.A(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n272), .ZN(new_n277));
  NOR2_X1   g076(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n259), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(KEYINPUT71), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n259), .A2(new_n283), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n284), .A2(new_n263), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n274), .A2(new_n281), .A3(new_n250), .A4(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT64), .B(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT23), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT65), .ZN(new_n292));
  INV_X1    g091(.A(new_n252), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(new_n253), .C1(G183gat), .C2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n263), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n260), .A2(new_n295), .A3(KEYINPUT25), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n289), .A2(new_n297), .A3(KEYINPUT23), .A4(new_n290), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n292), .A2(new_n294), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n267), .A2(new_n288), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n302));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n304), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n249), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n248), .B1(new_n307), .B2(KEYINPUT33), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n249), .A3(new_n306), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(new_n248), .C1(new_n307), .C2(KEYINPUT33), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n314));
  OR3_X1    g113(.A1(new_n307), .A2(new_n314), .A3(KEYINPUT34), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT34), .B1(new_n307), .B2(new_n314), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n311), .A2(new_n315), .A3(new_n312), .A4(new_n316), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT31), .B(G50gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT79), .ZN(new_n325));
  INV_X1    g124(.A(G22gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G141gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(G148gat), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n335), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n332), .A2(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n329), .B2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G155gat), .B(G162gat), .Z(new_n341));
  AOI22_X1  g140(.A1(new_n333), .A2(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT76), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G148gat), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n332), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n338), .B1(new_n348), .B2(new_n329), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n340), .A2(new_n341), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT76), .A4(new_n343), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n327), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  INV_X1    g153(.A(G204gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n236), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G197gat), .A2(G204gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n365), .A2(new_n366), .A3(new_n359), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n365), .B2(new_n359), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n359), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT72), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n356), .A2(new_n357), .B1(new_n360), .B2(new_n359), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(new_n366), .A3(new_n359), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n354), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n349), .A2(new_n350), .A3(new_n343), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n379), .B2(new_n351), .ZN(new_n380));
  INV_X1    g179(.A(new_n375), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n349), .A2(new_n350), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n369), .A2(new_n374), .A3(new_n327), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT80), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n387), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n349), .A2(new_n393), .A3(new_n350), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n393), .B1(new_n349), .B2(new_n350), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n351), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n381), .B1(new_n398), .B2(new_n327), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n326), .B1(new_n390), .B2(new_n401), .ZN(new_n402));
  AOI211_X1 g201(.A(G22gat), .B(new_n400), .C1(new_n386), .C2(new_n389), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n325), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n385), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n353), .A2(new_n375), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(KEYINPUT81), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n388), .B1(new_n407), .B2(new_n376), .ZN(new_n408));
  OAI21_X1  g207(.A(G22gat), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n326), .A3(new_n401), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n324), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n321), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT82), .B1(new_n413), .B2(new_n325), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n320), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G226gat), .ZN(new_n418));
  INV_X1    g217(.A(G233gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n300), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n267), .A2(new_n299), .A3(new_n288), .A4(KEYINPUT73), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n420), .A2(KEYINPUT29), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n300), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n375), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n300), .A2(new_n421), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n424), .ZN(new_n430));
  INV_X1    g229(.A(new_n426), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n429), .B(new_n381), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT30), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n437), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n304), .A2(new_n383), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n342), .A2(new_n393), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n444), .B2(new_n304), .ZN(new_n445));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT77), .B(KEYINPUT5), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(KEYINPUT3), .ZN(new_n448));
  INV_X1    g247(.A(new_n303), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n302), .B(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n379), .B2(new_n351), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n342), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n455), .A3(new_n342), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n446), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT77), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n304), .B1(new_n394), .B2(new_n395), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n446), .B1(new_n460), .B2(new_n453), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT78), .ZN(new_n465));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466));
  INV_X1    g265(.A(G85gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT0), .B(G57gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n447), .A2(new_n458), .A3(new_n463), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n458), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n465), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n464), .A2(KEYINPUT78), .B1(new_n474), .B2(new_n462), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n471), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g280(.A(new_n477), .B(new_n471), .C1(new_n479), .C2(new_n473), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n440), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT86), .B(new_n320), .C1(new_n412), .C2(new_n414), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n417), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  INV_X1    g286(.A(new_n439), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(new_n438), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n478), .A2(new_n480), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n482), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n415), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n428), .A2(KEYINPUT37), .A3(new_n432), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT37), .B1(new_n428), .B2(new_n432), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(new_n437), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT38), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT85), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(new_n437), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n496), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT38), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n375), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n425), .A2(new_n375), .A3(new_n427), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n488), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n506), .A2(new_n481), .A3(new_n483), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n404), .A2(new_n411), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g314(.A(new_n414), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n446), .B1(new_n452), .B2(new_n457), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n470), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n445), .A2(new_n446), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n448), .A2(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(KEYINPUT39), .C1(new_n522), .C2(new_n446), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n517), .B1(new_n524), .B2(KEYINPUT84), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526));
  AOI211_X1 g325(.A(new_n526), .B(KEYINPUT40), .C1(new_n520), .C2(new_n523), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n480), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n515), .A2(new_n516), .B1(new_n528), .B2(new_n440), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n318), .A2(KEYINPUT36), .A3(new_n319), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT36), .B1(new_n318), .B2(new_n319), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n489), .B1(new_n491), .B2(new_n482), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n412), .A2(new_n414), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n245), .B1(new_n495), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G134gat), .B(G162gat), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT91), .B(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(G92gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n467), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G99gat), .B(G106gat), .Z(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n542), .B1(new_n215), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n555), .A2(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(KEYINPUT92), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n224), .A2(new_n554), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n216), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT93), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n556), .A2(new_n557), .B1(new_n216), .B2(new_n559), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n563), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n541), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G64gat), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n569), .A2(G57gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(G57gat), .ZN(new_n571));
  AND2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  OAI22_X1  g371(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT9), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT90), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n580), .B(new_n584), .Z(new_n585));
  OAI21_X1  g384(.A(new_n223), .B1(new_n577), .B2(new_n576), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n561), .A2(KEYINPUT94), .A3(new_n564), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n566), .B2(new_n563), .ZN(new_n595));
  INV_X1    g394(.A(new_n541), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n566), .B2(new_n563), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n593), .A2(new_n595), .A3(new_n597), .A4(KEYINPUT95), .ZN(new_n601));
  AOI211_X1 g400(.A(new_n568), .B(new_n592), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n576), .B1(new_n552), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n554), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n552), .B(new_n553), .C1(new_n576), .C2(new_n604), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT10), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n554), .A2(new_n609), .A3(new_n576), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n603), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n606), .A2(G230gat), .A3(G233gat), .A4(new_n607), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n612), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n615), .B(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n538), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n481), .A2(new_n483), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT100), .B(G1gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1324gat));
  INV_X1    g430(.A(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n440), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(G8gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT16), .B(G8gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  MUX2_X1   g436(.A(new_n635), .B(KEYINPUT42), .S(new_n637), .Z(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n533), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n627), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n632), .A2(new_n320), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n639), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n632), .A2(new_n535), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT101), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT43), .B(G22gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  AOI21_X1  g446(.A(new_n568), .B1(new_n600), .B2(new_n601), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n592), .A3(new_n623), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n538), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n628), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT45), .Z(new_n654));
  INV_X1    g453(.A(new_n592), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n245), .A2(new_n655), .A3(new_n622), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n495), .A2(KEYINPUT103), .A3(new_n537), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n493), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n530), .A2(new_n536), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n495), .A2(new_n537), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n666), .B2(new_n649), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n656), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668), .B2(new_n628), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n669), .ZN(G1328gat));
  NOR3_X1   g469(.A1(new_n652), .A2(G36gat), .A3(new_n489), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT46), .ZN(new_n672));
  OAI21_X1  g471(.A(G36gat), .B1(new_n668), .B2(new_n489), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(G1329gat));
  INV_X1    g473(.A(G43gat), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n533), .B(new_n656), .C1(new_n664), .C2(new_n667), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n538), .A2(new_n675), .A3(new_n320), .A4(new_n651), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(KEYINPUT47), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(G43gat), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(KEYINPUT47), .B2(new_n683), .ZN(G1330gat));
  INV_X1    g483(.A(new_n535), .ZN(new_n685));
  OAI21_X1  g484(.A(G50gat), .B1(new_n668), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(G50gat), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT105), .Z(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  OAI22_X1  g489(.A1(new_n652), .A2(new_n689), .B1(new_n690), .B2(KEYINPUT48), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(KEYINPUT48), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT107), .Z(new_n695));
  XOR2_X1   g494(.A(new_n693), .B(new_n695), .Z(G1331gat));
  NOR2_X1   g495(.A1(new_n623), .A2(new_n244), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n602), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n659), .B2(new_n663), .ZN(new_n699));
  INV_X1    g498(.A(new_n628), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g501(.A(new_n489), .B(KEYINPUT108), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT49), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n569), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n569), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1333gat));
  AOI21_X1  g508(.A(G71gat), .B1(new_n699), .B2(new_n320), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n533), .A2(G71gat), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n699), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1334gat));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n535), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g515(.A1(new_n623), .A2(new_n244), .A3(new_n655), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n664), .B2(new_n667), .ZN(new_n718));
  OAI21_X1  g517(.A(G85gat), .B1(new_n718), .B2(new_n628), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n649), .B1(new_n661), .B2(new_n662), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT111), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n722), .B(new_n649), .C1(new_n661), .C2(new_n662), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n655), .B(new_n244), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n728), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n721), .A2(new_n730), .A3(new_n723), .A4(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n628), .A2(new_n623), .A3(G85gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT113), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n719), .B1(new_n732), .B2(new_n734), .ZN(G1336gat));
  OAI211_X1 g534(.A(new_n703), .B(new_n717), .C1(new_n664), .C2(new_n667), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT52), .B1(new_n736), .B2(G92gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n703), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(G92gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n729), .A2(new_n622), .A3(new_n731), .A4(new_n739), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n440), .B(new_n717), .C1(new_n664), .C2(new_n667), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G92gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT114), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT52), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n737), .A2(new_n740), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n746), .A2(new_n751), .ZN(G1337gat));
  INV_X1    g551(.A(new_n320), .ZN(new_n753));
  OR4_X1    g552(.A1(G99gat), .A2(new_n732), .A3(new_n753), .A4(new_n623), .ZN(new_n754));
  OAI21_X1  g553(.A(G99gat), .B1(new_n718), .B2(new_n640), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1338gat));
  OAI211_X1 g555(.A(new_n535), .B(new_n717), .C1(new_n664), .C2(new_n667), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n757), .A2(G106gat), .B1(KEYINPUT115), .B2(KEYINPUT53), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n685), .A2(G106gat), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n729), .A2(new_n622), .A3(new_n731), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1339gat));
  NAND4_X1  g562(.A1(new_n648), .A2(new_n245), .A3(new_n655), .A4(new_n623), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n602), .A2(KEYINPUT116), .A3(new_n245), .A4(new_n623), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n617), .B(KEYINPUT97), .Z(new_n770));
  OR3_X1    g569(.A1(new_n608), .A2(new_n603), .A3(new_n610), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(KEYINPUT54), .A3(new_n611), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n603), .C1(new_n608), .C2(new_n610), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n774), .A2(KEYINPUT117), .A3(new_n615), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT117), .B1(new_n774), .B2(new_n615), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT55), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n779), .B(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n770), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n244), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n227), .A2(new_n228), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n231), .A2(new_n232), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n239), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n622), .A2(new_n242), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n649), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n777), .A2(KEYINPUT55), .ZN(new_n788));
  INV_X1    g587(.A(new_n780), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n618), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n242), .A2(new_n785), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n648), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n592), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n769), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n415), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n794), .A2(new_n700), .A3(new_n795), .A4(new_n738), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n796), .B2(new_n245), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT118), .Z(new_n798));
  AND2_X1   g597(.A1(new_n769), .A2(new_n793), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n417), .A2(new_n485), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n628), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n738), .ZN(new_n802));
  INV_X1    g601(.A(G113gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n244), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n804), .ZN(G1340gat));
  INV_X1    g604(.A(G120gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n806), .A3(new_n622), .ZN(new_n807));
  OAI21_X1  g606(.A(G120gat), .B1(new_n796), .B2(new_n623), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1341gat));
  INV_X1    g608(.A(G127gat), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n796), .A2(new_n810), .A3(new_n592), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n802), .A2(new_n655), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n810), .ZN(G1342gat));
  NAND2_X1  g612(.A1(new_n649), .A2(new_n489), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(G134gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT56), .Z(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n796), .B2(new_n648), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT119), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(KEYINPUT119), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(G1343gat));
  NAND2_X1  g620(.A1(new_n700), .A2(new_n640), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n703), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n794), .A2(new_n535), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n332), .A3(new_n244), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n794), .A2(new_n535), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n827), .B2(KEYINPUT57), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n244), .B1(new_n781), .B2(KEYINPUT120), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n831), .B(new_n770), .C1(new_n778), .C2(new_n780), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n786), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n792), .B1(new_n833), .B2(new_n648), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n769), .B1(new_n834), .B2(new_n655), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(new_n535), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n828), .A2(new_n836), .A3(new_n245), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n826), .B1(new_n837), .B2(new_n332), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g638(.A(new_n331), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n840), .A3(new_n622), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n829), .B1(new_n794), .B2(new_n535), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n626), .A2(new_n245), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n592), .B1(new_n834), .B2(KEYINPUT122), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n846), .B(new_n792), .C1(new_n833), .C2(new_n648), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n685), .A2(KEYINPUT57), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n623), .B(new_n843), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n823), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n842), .B1(new_n851), .B2(G148gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n828), .A2(new_n836), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT59), .B(new_n840), .C1(new_n853), .C2(new_n622), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n841), .B1(new_n852), .B2(new_n854), .ZN(G1345gat));
  AOI21_X1  g654(.A(G155gat), .B1(new_n825), .B2(new_n655), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n592), .A2(new_n335), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1346gat));
  OR4_X1    g657(.A1(G162gat), .A2(new_n827), .A3(new_n814), .A4(new_n822), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n828), .A2(new_n836), .A3(new_n648), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n336), .ZN(G1347gat));
  NOR4_X1   g660(.A1(new_n799), .A2(new_n700), .A3(new_n800), .A4(new_n738), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n244), .A3(new_n289), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n700), .B1(new_n769), .B2(new_n793), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n440), .A3(new_n795), .ZN(new_n865));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865), .B2(new_n245), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(G1348gat));
  NOR3_X1   g666(.A1(new_n865), .A2(new_n290), .A3(new_n623), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n862), .A2(new_n622), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n290), .ZN(G1349gat));
  OAI211_X1 g669(.A(new_n862), .B(new_n655), .C1(new_n278), .C2(new_n277), .ZN(new_n871));
  OAI21_X1  g670(.A(G183gat), .B1(new_n865), .B2(new_n592), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(KEYINPUT123), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n865), .B2(new_n648), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT61), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n862), .A2(new_n276), .A3(new_n649), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1351gat));
  NAND2_X1  g677(.A1(new_n848), .A2(new_n849), .ZN(new_n879));
  INV_X1    g678(.A(new_n843), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n700), .A2(new_n489), .A3(new_n533), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G197gat), .B1(new_n882), .B2(new_n245), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n685), .A2(new_n533), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n703), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n236), .A3(new_n244), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(G1352gat));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n355), .B1(new_n850), .B2(new_n881), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n623), .A2(G204gat), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n864), .A2(new_n703), .A3(new_n884), .A4(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT62), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n892), .B2(KEYINPUT62), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n895), .A2(new_n896), .B1(KEYINPUT62), .B2(new_n892), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n889), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n892), .A2(KEYINPUT62), .ZN(new_n899));
  INV_X1    g698(.A(new_n896), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n894), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n622), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n901), .B(KEYINPUT125), .C1(new_n902), .C2(new_n355), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n898), .A2(new_n903), .ZN(G1353gat));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n363), .A3(new_n655), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n879), .A2(new_n880), .A3(new_n655), .A4(new_n881), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT63), .B1(new_n906), .B2(G211gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1354gat));
  OAI21_X1  g708(.A(new_n364), .B1(new_n885), .B2(new_n648), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT126), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n882), .A2(KEYINPUT127), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n649), .A2(G218gat), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n882), .A2(KEYINPUT127), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(G1355gat));
endmodule


