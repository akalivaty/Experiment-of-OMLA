

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n609), .A2(n608), .ZN(n623) );
  XNOR2_X1 U553 ( .A(n630), .B(n629), .ZN(n633) );
  XNOR2_X1 U554 ( .A(n648), .B(KEYINPUT30), .ZN(n650) );
  NAND2_X1 U555 ( .A1(n665), .A2(n664), .ZN(n667) );
  OR2_X1 U556 ( .A1(n657), .A2(n720), .ZN(n519) );
  OR2_X1 U557 ( .A1(n681), .A2(KEYINPUT33), .ZN(n520) );
  XOR2_X1 U558 ( .A(KEYINPUT31), .B(n654), .Z(n521) );
  INV_X1 U559 ( .A(KEYINPUT94), .ZN(n629) );
  AND2_X1 U560 ( .A1(n692), .A2(n691), .ZN(n640) );
  INV_X1 U561 ( .A(G168), .ZN(n649) );
  AND2_X1 U562 ( .A1(n650), .A2(n649), .ZN(n653) );
  INV_X1 U563 ( .A(KEYINPUT32), .ZN(n666) );
  NOR2_X1 U564 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U565 ( .A1(n721), .A2(n519), .ZN(n722) );
  NOR2_X2 U566 ( .A1(G2105), .A2(n526), .ZN(n881) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(n523), .ZN(n884) );
  NOR2_X1 U568 ( .A1(G651), .A2(n573), .ZN(n797) );
  INV_X1 U569 ( .A(KEYINPUT40), .ZN(n753) );
  INV_X1 U570 ( .A(G2104), .ZN(n526) );
  AND2_X1 U571 ( .A1(n526), .A2(G2105), .ZN(n876) );
  NAND2_X1 U572 ( .A1(n876), .A2(G125), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U574 ( .A(n522), .B(KEYINPUT64), .Z(n523) );
  NAND2_X1 U575 ( .A1(G137), .A2(n884), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n531) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  NAND2_X1 U578 ( .A1(n877), .A2(G113), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G101), .A2(n881), .ZN(n527) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n527), .Z(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G160) );
  NOR2_X1 U583 ( .A1(G543), .A2(G651), .ZN(n802) );
  NAND2_X1 U584 ( .A1(n802), .A2(G89), .ZN(n532) );
  XNOR2_X1 U585 ( .A(n532), .B(KEYINPUT4), .ZN(n534) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n573) );
  INV_X1 U587 ( .A(G651), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n573), .A2(n536), .ZN(n801) );
  NAND2_X1 U589 ( .A1(G76), .A2(n801), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n535), .B(KEYINPUT5), .ZN(n543) );
  NAND2_X1 U592 ( .A1(G51), .A2(n797), .ZN(n540) );
  NOR2_X1 U593 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U594 ( .A(KEYINPUT66), .B(n537), .Z(n538) );
  XNOR2_X1 U595 ( .A(KEYINPUT1), .B(n538), .ZN(n798) );
  NAND2_X1 U596 ( .A1(G63), .A2(n798), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n544), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U601 ( .A1(n881), .A2(G102), .ZN(n546) );
  NAND2_X1 U602 ( .A1(G138), .A2(n884), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G126), .A2(n876), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G114), .A2(n877), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n550), .A2(n549), .ZN(G164) );
  NAND2_X1 U608 ( .A1(G78), .A2(n801), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G53), .A2(n797), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n802), .A2(G91), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT68), .B(n553), .Z(n554) );
  NOR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G65), .A2(n798), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U616 ( .A1(G52), .A2(n797), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G64), .A2(n798), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G77), .A2(n801), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G90), .A2(n802), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U622 ( .A(KEYINPUT9), .B(n562), .ZN(n563) );
  XNOR2_X1 U623 ( .A(KEYINPUT67), .B(n563), .ZN(n564) );
  NOR2_X1 U624 ( .A1(n565), .A2(n564), .ZN(G171) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U626 ( .A1(G50), .A2(n797), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G62), .A2(n798), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G75), .A2(n801), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G88), .A2(n802), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n572), .B(KEYINPUT76), .ZN(G166) );
  INV_X1 U634 ( .A(G166), .ZN(G303) );
  NAND2_X1 U635 ( .A1(G87), .A2(n573), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U638 ( .A1(n798), .A2(n576), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n797), .A2(G49), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U641 ( .A1(n801), .A2(G73), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT2), .B(n579), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G86), .A2(n802), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G61), .A2(n798), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT74), .B(n582), .Z(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U648 ( .A(n585), .B(KEYINPUT75), .ZN(n587) );
  NAND2_X1 U649 ( .A1(G48), .A2(n797), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G85), .A2(n802), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G60), .A2(n798), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G72), .A2(n801), .ZN(n590) );
  XNOR2_X1 U655 ( .A(KEYINPUT65), .B(n590), .ZN(n591) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n797), .A2(G47), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(G290) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n692) );
  NAND2_X1 U660 ( .A1(G40), .A2(G160), .ZN(n595) );
  XNOR2_X1 U661 ( .A(KEYINPUT81), .B(n595), .ZN(n691) );
  NAND2_X1 U662 ( .A1(n692), .A2(n691), .ZN(n658) );
  NAND2_X1 U663 ( .A1(n658), .A2(G1341), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n596), .B(KEYINPUT96), .ZN(n606) );
  NAND2_X1 U665 ( .A1(n802), .A2(G81), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n597), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U667 ( .A1(G68), .A2(n801), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n600), .B(KEYINPUT13), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G43), .A2(n797), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n798), .A2(G56), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT14), .B(n603), .Z(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n944) );
  NAND2_X1 U675 ( .A1(n606), .A2(n944), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G1996), .A2(n640), .ZN(n607) );
  XOR2_X1 U677 ( .A(n607), .B(KEYINPUT26), .Z(n608) );
  NAND2_X1 U678 ( .A1(G79), .A2(n801), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G92), .A2(n802), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G54), .A2(n797), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G66), .A2(n798), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U685 ( .A(KEYINPUT15), .B(n616), .Z(n900) );
  NAND2_X1 U686 ( .A1(n623), .A2(n900), .ZN(n621) );
  AND2_X1 U687 ( .A1(n640), .A2(G2067), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n617), .B(KEYINPUT97), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n658), .A2(G1348), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n622), .B(KEYINPUT98), .ZN(n625) );
  OR2_X1 U693 ( .A1(n900), .A2(n623), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n632) );
  INV_X1 U695 ( .A(G299), .ZN(n943) );
  NAND2_X1 U696 ( .A1(n640), .A2(G2072), .ZN(n626) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(n626), .Z(n628) );
  NAND2_X1 U698 ( .A1(G1956), .A2(n658), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n943), .A2(n633), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n637) );
  NOR2_X1 U702 ( .A1(n943), .A2(n633), .ZN(n635) );
  XNOR2_X1 U703 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U705 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U706 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n645) );
  XOR2_X1 U708 ( .A(G2078), .B(KEYINPUT25), .Z(n970) );
  NOR2_X1 U709 ( .A1(n970), .A2(n658), .ZN(n642) );
  XNOR2_X1 U710 ( .A(KEYINPUT92), .B(G1961), .ZN(n1000) );
  NOR2_X1 U711 ( .A1(n640), .A2(n1000), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U713 ( .A(KEYINPUT93), .B(n643), .ZN(n651) );
  NAND2_X1 U714 ( .A1(n651), .A2(G171), .ZN(n644) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n655) );
  NAND2_X1 U716 ( .A1(G8), .A2(n658), .ZN(n657) );
  NOR2_X1 U717 ( .A1(n657), .A2(G1966), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT91), .ZN(n669) );
  INV_X1 U719 ( .A(G8), .ZN(n663) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n658), .ZN(n668) );
  NOR2_X1 U721 ( .A1(n663), .A2(n668), .ZN(n647) );
  AND2_X1 U722 ( .A1(n669), .A2(n647), .ZN(n648) );
  NOR2_X1 U723 ( .A1(G171), .A2(n651), .ZN(n652) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n521), .ZN(n670) );
  AND2_X1 U726 ( .A1(G286), .A2(G8), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n670), .A2(n656), .ZN(n665) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n657), .ZN(n660) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n658), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U731 ( .A1(G303), .A2(n661), .ZN(n662) );
  OR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n667), .B(n666), .ZN(n674) );
  NAND2_X1 U734 ( .A1(G8), .A2(n668), .ZN(n672) );
  AND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U738 ( .A(n675), .B(KEYINPUT100), .ZN(n725) );
  NOR2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n719) );
  NOR2_X1 U740 ( .A1(G303), .A2(G1971), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n719), .A2(n676), .ZN(n950) );
  NAND2_X1 U742 ( .A1(n725), .A2(n950), .ZN(n677) );
  XNOR2_X1 U743 ( .A(n677), .B(KEYINPUT101), .ZN(n680) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n949) );
  INV_X1 U745 ( .A(n657), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n949), .A2(n678), .ZN(n679) );
  XOR2_X1 U747 ( .A(G1981), .B(G305), .Z(n939) );
  NAND2_X1 U748 ( .A1(G128), .A2(n876), .ZN(n683) );
  NAND2_X1 U749 ( .A1(G116), .A2(n877), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n684), .B(KEYINPUT35), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n881), .A2(G104), .ZN(n686) );
  NAND2_X1 U753 ( .A1(G140), .A2(n884), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U755 ( .A(KEYINPUT34), .B(n687), .Z(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT36), .ZN(n896) );
  XOR2_X1 U758 ( .A(KEYINPUT37), .B(G2067), .Z(n734) );
  NAND2_X1 U759 ( .A1(n896), .A2(n734), .ZN(n922) );
  INV_X1 U760 ( .A(n691), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(KEYINPUT82), .ZN(n748) );
  INV_X1 U763 ( .A(n748), .ZN(n717) );
  NOR2_X1 U764 ( .A1(n922), .A2(n717), .ZN(n695) );
  XNOR2_X1 U765 ( .A(n695), .B(KEYINPUT83), .ZN(n741) );
  NAND2_X1 U766 ( .A1(G119), .A2(n876), .ZN(n697) );
  NAND2_X1 U767 ( .A1(G107), .A2(n877), .ZN(n696) );
  NAND2_X1 U768 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U769 ( .A(KEYINPUT84), .B(n698), .Z(n702) );
  NAND2_X1 U770 ( .A1(n884), .A2(G131), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n881), .A2(G95), .ZN(n699) );
  AND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n892) );
  AND2_X1 U774 ( .A1(n892), .A2(G1991), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n877), .A2(G117), .ZN(n703) );
  XOR2_X1 U776 ( .A(KEYINPUT85), .B(n703), .Z(n705) );
  NAND2_X1 U777 ( .A1(n876), .A2(G129), .ZN(n704) );
  NAND2_X1 U778 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U779 ( .A(KEYINPUT86), .B(n706), .ZN(n711) );
  XOR2_X1 U780 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n708) );
  NAND2_X1 U781 ( .A1(G105), .A2(n881), .ZN(n707) );
  XNOR2_X1 U782 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U783 ( .A(KEYINPUT87), .B(n709), .Z(n710) );
  NOR2_X1 U784 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U785 ( .A1(G141), .A2(n884), .ZN(n712) );
  NAND2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U787 ( .A(KEYINPUT89), .B(n714), .Z(n889) );
  AND2_X1 U788 ( .A1(n889), .A2(G1996), .ZN(n715) );
  NOR2_X1 U789 ( .A1(n716), .A2(n715), .ZN(n916) );
  NOR2_X1 U790 ( .A1(n717), .A2(n916), .ZN(n738) );
  INV_X1 U791 ( .A(n738), .ZN(n718) );
  AND2_X1 U792 ( .A1(n741), .A2(n718), .ZN(n733) );
  AND2_X1 U793 ( .A1(n939), .A2(n733), .ZN(n721) );
  NAND2_X1 U794 ( .A1(n719), .A2(KEYINPUT33), .ZN(n720) );
  NAND2_X1 U795 ( .A1(n520), .A2(n722), .ZN(n747) );
  NOR2_X1 U796 ( .A1(G303), .A2(G2090), .ZN(n723) );
  NAND2_X1 U797 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U799 ( .A1(n726), .A2(n657), .ZN(n731) );
  NOR2_X1 U800 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U801 ( .A(n727), .B(KEYINPUT90), .Z(n728) );
  XNOR2_X1 U802 ( .A(KEYINPUT24), .B(n728), .ZN(n729) );
  OR2_X1 U803 ( .A1(n657), .A2(n729), .ZN(n730) );
  NAND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n745) );
  NOR2_X1 U806 ( .A1(n896), .A2(n734), .ZN(n735) );
  XOR2_X1 U807 ( .A(KEYINPUT102), .B(n735), .Z(n931) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n889), .ZN(n925) );
  NOR2_X1 U809 ( .A1(G1991), .A2(n892), .ZN(n921) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n921), .A2(n736), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n925), .A2(n739), .ZN(n740) );
  XNOR2_X1 U814 ( .A(n740), .B(KEYINPUT39), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n931), .A2(n743), .ZN(n744) );
  AND2_X1 U817 ( .A1(n744), .A2(n748), .ZN(n750) );
  NOR2_X1 U818 ( .A1(n745), .A2(n750), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n747), .A2(n746), .ZN(n752) );
  XNOR2_X1 U820 ( .A(G1986), .B(G290), .ZN(n948) );
  NAND2_X1 U821 ( .A1(n948), .A2(n748), .ZN(n749) );
  OR2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n754) );
  XNOR2_X1 U824 ( .A(n754), .B(n753), .ZN(G329) );
  XOR2_X1 U825 ( .A(G2438), .B(KEYINPUT104), .Z(n756) );
  XNOR2_X1 U826 ( .A(G2454), .B(G2435), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n756), .B(n755), .ZN(n757) );
  XOR2_X1 U828 ( .A(n757), .B(G2430), .Z(n759) );
  XNOR2_X1 U829 ( .A(G1341), .B(G1348), .ZN(n758) );
  XNOR2_X1 U830 ( .A(n759), .B(n758), .ZN(n763) );
  XOR2_X1 U831 ( .A(G2446), .B(KEYINPUT105), .Z(n761) );
  XNOR2_X1 U832 ( .A(G2451), .B(G2427), .ZN(n760) );
  XNOR2_X1 U833 ( .A(n761), .B(n760), .ZN(n762) );
  XOR2_X1 U834 ( .A(n763), .B(n762), .Z(n765) );
  XNOR2_X1 U835 ( .A(KEYINPUT103), .B(G2443), .ZN(n764) );
  XNOR2_X1 U836 ( .A(n765), .B(n764), .ZN(n766) );
  AND2_X1 U837 ( .A1(n766), .A2(G14), .ZN(G401) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  INV_X1 U840 ( .A(G132), .ZN(G219) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  XOR2_X1 U842 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n768) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U844 ( .A(n768), .B(n767), .ZN(G223) );
  INV_X1 U845 ( .A(G223), .ZN(n828) );
  NAND2_X1 U846 ( .A1(n828), .A2(G567), .ZN(n769) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  NAND2_X1 U848 ( .A1(n944), .A2(G860), .ZN(G153) );
  INV_X1 U849 ( .A(G171), .ZN(G301) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U851 ( .A(n900), .ZN(n956) );
  INV_X1 U852 ( .A(G868), .ZN(n810) );
  NAND2_X1 U853 ( .A1(n956), .A2(n810), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n771), .A2(n770), .ZN(G284) );
  NOR2_X1 U855 ( .A1(G286), .A2(n810), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G868), .A2(G299), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G297) );
  INV_X1 U858 ( .A(G860), .ZN(n837) );
  NAND2_X1 U859 ( .A1(n837), .A2(G559), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n774), .A2(n900), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U862 ( .A1(n900), .A2(G868), .ZN(n776) );
  NOR2_X1 U863 ( .A1(G559), .A2(n776), .ZN(n778) );
  AND2_X1 U864 ( .A1(n810), .A2(n944), .ZN(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(G282) );
  XOR2_X1 U866 ( .A(KEYINPUT70), .B(KEYINPUT18), .Z(n780) );
  NAND2_X1 U867 ( .A1(G123), .A2(n876), .ZN(n779) );
  XNOR2_X1 U868 ( .A(n780), .B(n779), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n877), .A2(G111), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G135), .A2(n884), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n881), .A2(G99), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n918) );
  XOR2_X1 U875 ( .A(n918), .B(G2096), .Z(n788) );
  XNOR2_X1 U876 ( .A(G2100), .B(KEYINPUT71), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G559), .A2(n900), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n789), .B(KEYINPUT72), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n944), .B(n790), .ZN(n836) );
  XNOR2_X1 U881 ( .A(KEYINPUT19), .B(KEYINPUT77), .ZN(n792) );
  XNOR2_X1 U882 ( .A(G288), .B(KEYINPUT78), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n792), .B(n791), .ZN(n793) );
  XNOR2_X1 U884 ( .A(n943), .B(n793), .ZN(n795) );
  XNOR2_X1 U885 ( .A(G290), .B(G303), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n795), .B(n794), .ZN(n796) );
  XNOR2_X1 U887 ( .A(n796), .B(G305), .ZN(n808) );
  NAND2_X1 U888 ( .A1(G55), .A2(n797), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G67), .A2(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G80), .A2(n801), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(KEYINPUT73), .ZN(n838) );
  XNOR2_X1 U896 ( .A(n808), .B(n838), .ZN(n903) );
  XNOR2_X1 U897 ( .A(n836), .B(n903), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n809), .A2(G868), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n838), .A2(n810), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n817) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n817), .Z(n818) );
  NOR2_X1 U909 ( .A1(G218), .A2(n818), .ZN(n819) );
  NAND2_X1 U910 ( .A1(G96), .A2(n819), .ZN(n835) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n835), .ZN(n824) );
  NAND2_X1 U912 ( .A1(G120), .A2(G69), .ZN(n820) );
  NOR2_X1 U913 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U914 ( .A1(G108), .A2(n821), .ZN(n834) );
  NAND2_X1 U915 ( .A1(G567), .A2(n834), .ZN(n822) );
  XOR2_X1 U916 ( .A(KEYINPUT79), .B(n822), .Z(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U918 ( .A(KEYINPUT80), .B(n825), .Z(G319) );
  INV_X1 U919 ( .A(G319), .ZN(n827) );
  NAND2_X1 U920 ( .A1(G661), .A2(G483), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n833) );
  NAND2_X1 U922 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n828), .ZN(G217) );
  INV_X1 U924 ( .A(G661), .ZN(n830) );
  NAND2_X1 U925 ( .A1(G2), .A2(G15), .ZN(n829) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U927 ( .A(KEYINPUT106), .B(n831), .Z(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U930 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  NAND2_X1 U936 ( .A1(n837), .A2(n836), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(G145) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1966), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n842), .B(G2474), .Z(n844) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(G1981), .Z(n846) );
  XNOR2_X1 U945 ( .A(G1956), .B(G1961), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U948 ( .A(G2100), .B(G2096), .Z(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2072), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2084), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(G227) );
  NAND2_X1 U957 ( .A1(G112), .A2(n877), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(KEYINPUT108), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G124), .A2(n876), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n881), .A2(G100), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G136), .A2(n884), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n875) );
  NAND2_X1 U967 ( .A1(n881), .A2(G106), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G142), .A2(n884), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT45), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G130), .A2(n876), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G118), .A2(n877), .ZN(n870) );
  XNOR2_X1 U974 ( .A(KEYINPUT109), .B(n870), .ZN(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n873), .B(KEYINPUT110), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G127), .A2(n876), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G115), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n880), .B(KEYINPUT47), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G103), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G139), .A2(n884), .ZN(n885) );
  XNOR2_X1 U985 ( .A(KEYINPUT111), .B(n885), .ZN(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n912) );
  XOR2_X1 U987 ( .A(n888), .B(n912), .Z(n891) );
  XOR2_X1 U988 ( .A(G164), .B(n889), .Z(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n895) );
  XNOR2_X1 U990 ( .A(G162), .B(n892), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(n918), .ZN(n894) );
  XOR2_X1 U992 ( .A(n895), .B(n894), .Z(n898) );
  XNOR2_X1 U993 ( .A(G160), .B(n896), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U996 ( .A(G286), .B(G171), .Z(n902) );
  XNOR2_X1 U997 ( .A(n900), .B(n944), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n906) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n906), .Z(n907) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n907), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n908), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(KEYINPUT112), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1010 ( .A(G2072), .B(n912), .Z(n914) );
  XOR2_X1 U1011 ( .A(G164), .B(G2078), .Z(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT50), .B(n915), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n933) );
  XNOR2_X1 U1015 ( .A(G160), .B(G2084), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n929) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G162), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(KEYINPUT113), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT51), .B(n927), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1026 ( .A(KEYINPUT52), .B(n934), .Z(n935) );
  NOR2_X1 U1027 ( .A1(KEYINPUT55), .A2(n935), .ZN(n936) );
  XOR2_X1 U1028 ( .A(KEYINPUT114), .B(n936), .Z(n937) );
  NAND2_X1 U1029 ( .A1(G29), .A2(n937), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(KEYINPUT115), .B(n938), .ZN(n1021) );
  XNOR2_X1 U1031 ( .A(KEYINPUT56), .B(G16), .ZN(n965) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G168), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT57), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT118), .B(n942), .ZN(n963) );
  XNOR2_X1 U1036 ( .A(n943), .B(G1956), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(n944), .B(G1341), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n955) );
  AND2_X1 U1040 ( .A1(G303), .A2(G1971), .ZN(n952) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(n953), .B(KEYINPUT120), .ZN(n954) );
  NAND2_X1 U1044 ( .A1(n955), .A2(n954), .ZN(n961) );
  XNOR2_X1 U1045 ( .A(n956), .B(G1348), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(G301), .B(G1961), .ZN(n957) );
  NOR2_X1 U1047 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(n959), .B(KEYINPUT119), .ZN(n960) );
  NOR2_X1 U1049 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1050 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1052 ( .A1(n966), .A2(G11), .ZN(n988) );
  XOR2_X1 U1053 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n985) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G35), .ZN(n979) );
  XOR2_X1 U1055 ( .A(G25), .B(G1991), .Z(n967) );
  NAND2_X1 U1056 ( .A1(n967), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1057 ( .A(G1996), .B(G32), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n974) );
  XNOR2_X1 U1060 ( .A(G2067), .B(G26), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G27), .B(n970), .ZN(n971) );
  NOR2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n977), .ZN(n978) );
  NOR2_X1 U1066 ( .A1(n979), .A2(n978), .ZN(n983) );
  XOR2_X1 U1067 ( .A(G34), .B(KEYINPUT116), .Z(n981) );
  XNOR2_X1 U1068 ( .A(G2084), .B(KEYINPUT54), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n981), .B(n980), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(n985), .B(n984), .ZN(n986) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n986), .ZN(n987) );
  NOR2_X1 U1073 ( .A1(n988), .A2(n987), .ZN(n1018) );
  XOR2_X1 U1074 ( .A(KEYINPUT123), .B(G4), .Z(n990) );
  XNOR2_X1 U1075 ( .A(G1348), .B(KEYINPUT59), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(n990), .B(n989), .ZN(n994) );
  XNOR2_X1 U1077 ( .A(G1341), .B(G19), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G6), .B(G1981), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n997) );
  XNOR2_X1 U1081 ( .A(KEYINPUT122), .B(G1956), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(G20), .B(n995), .ZN(n996) );
  NOR2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT60), .B(n998), .ZN(n1009) );
  XOR2_X1 U1085 ( .A(KEYINPUT121), .B(G5), .Z(n999) );
  XNOR2_X1 U1086 ( .A(n1000), .B(n999), .ZN(n1007) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XOR2_X1 U1090 ( .A(G1986), .B(G24), .Z(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(G1966), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G21), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(KEYINPUT61), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT125), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(G16), .A2(n1015), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1016), .Z(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1019), .Z(n1020) );
  NOR2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

