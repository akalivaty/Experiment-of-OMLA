//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n623, new_n624, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  XNOR2_X1  g016(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g027(.A1(G221), .A2(G218), .A3(G219), .ZN(new_n453));
  NAND3_X1  g028(.A1(new_n437), .A2(new_n453), .A3(new_n438), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(G137), .ZN(new_n470));
  OAI221_X1 g045(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n466), .A2(new_n464), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n473), .B2(new_n474), .ZN(new_n480));
  AND2_X1   g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n465), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n469), .A2(new_n465), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND3_X1  g069(.A1(new_n485), .A2(G126), .A3(G2105), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n465), .A2(G138), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n485), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n485), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n507), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n513), .A2(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n508), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n524));
  XOR2_X1   g099(.A(new_n524), .B(KEYINPUT69), .Z(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT70), .B(G51), .Z(new_n529));
  OAI221_X1 g104(.A(new_n527), .B1(new_n519), .B2(new_n528), .C1(new_n513), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n510), .B2(new_n511), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n534), .B1(new_n535), .B2(new_n519), .C1(new_n536), .C2(new_n507), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OR2_X1    g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(G43), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n512), .A2(new_n505), .A3(G81), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n516), .A2(new_n515), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n533), .A2(G53), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n533), .B2(G53), .ZN(new_n564));
  OAI221_X1 g139(.A(new_n559), .B1(new_n560), .B2(new_n519), .C1(new_n562), .C2(new_n564), .ZN(G299));
  OR2_X1    g140(.A1(new_n525), .A2(new_n530), .ZN(G286));
  AOI22_X1  g141(.A1(new_n540), .A2(new_n541), .B1(new_n510), .B2(new_n511), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n533), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT71), .B1(new_n556), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n505), .A2(new_n574), .A3(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n567), .A2(G86), .B1(new_n533), .B2(G48), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n507), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n513), .A2(new_n586), .B1(new_n519), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(G301), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n556), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT72), .B1(new_n519), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n512), .A2(new_n505), .A3(new_n600), .A4(G92), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n599), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n597), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT73), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT74), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n599), .A2(new_n604), .A3(new_n601), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n604), .B1(new_n599), .B2(new_n601), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n596), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT73), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n592), .B1(new_n615), .B2(new_n591), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT75), .Z(G284));
  NAND2_X1  g192(.A1(G299), .A2(new_n591), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n591), .B2(G168), .ZN(G297));
  XNOR2_X1  g194(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g200(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n626));
  XNOR2_X1  g201(.A(G323), .B(new_n626), .ZN(G282));
  NAND3_X1  g202(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n487), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n489), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n465), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT78), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT79), .Z(G156));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  INV_X1    g222(.A(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT81), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT82), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(new_n652), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n655), .B2(new_n661), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n646), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n660), .B1(new_n659), .B2(new_n652), .ZN(new_n666));
  AND4_X1   g241(.A1(new_n660), .A2(new_n652), .A3(KEYINPUT14), .A4(new_n653), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n657), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n645), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n671), .A2(G14), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n665), .B1(new_n664), .B2(new_n670), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2072), .B(G2078), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2096), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT84), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT18), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(KEYINPUT17), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n676), .A2(new_n677), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n684), .B(new_n688), .Z(G227));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1961), .B(G1966), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n692), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n701), .A3(new_n696), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n694), .A2(new_n695), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n693), .A2(new_n697), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n694), .A3(new_n695), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n691), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n710), .A2(new_n703), .A3(new_n690), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1991), .B(G1996), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  INV_X1    g290(.A(new_n713), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n709), .A2(new_n716), .A3(new_n711), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n715), .B1(new_n714), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(G229));
  OR2_X1    g295(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n721), .A2(G16), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G24), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(G16), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G1986), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(G1986), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n485), .A2(G131), .A3(new_n465), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n485), .A2(G119), .A3(G2105), .ZN(new_n731));
  OR2_X1    g306(.A1(G95), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(new_n728), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(KEYINPUT88), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n727), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n582), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G6), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT32), .B(G1981), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G22), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G166), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G1971), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n742), .A2(new_n744), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(G23), .ZN(new_n752));
  INV_X1    g327(.A(G288), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n746), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT33), .B(G1976), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT86), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n745), .A2(new_n750), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n726), .B(new_n740), .C1(new_n758), .C2(KEYINPUT34), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(KEYINPUT34), .B2(new_n758), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT88), .B1(new_n761), .B2(new_n738), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n746), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n615), .B2(new_n746), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT89), .B(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n728), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n728), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT29), .B(G2090), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G5), .A2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT94), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G171), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1961), .ZN(new_n775));
  NOR2_X1   g350(.A1(G27), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(G29), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G2078), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT30), .B(G28), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n779), .A2(new_n728), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n782), .B1(new_n728), .B2(new_n636), .C1(new_n777), .C2(G2078), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n771), .A2(new_n775), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n485), .A2(G141), .A3(new_n465), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n485), .A2(G129), .A3(G2105), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G32), .B(new_n790), .S(G29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT27), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1996), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G34), .ZN(new_n796));
  AOI21_X1  g371(.A(G29), .B1(new_n795), .B2(G34), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n483), .A2(G29), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2084), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n746), .A2(G19), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n549), .B2(new_n746), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1341), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n728), .A2(G26), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT28), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n485), .A2(G140), .A3(new_n465), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n485), .A2(G128), .A3(G2105), .ZN(new_n806));
  OR2_X1    g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(new_n728), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2067), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n784), .A2(new_n793), .A3(new_n799), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(G115), .A2(G2104), .ZN(new_n815));
  INV_X1    g390(.A(G127), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n469), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G2105), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G139), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n818), .B(new_n821), .C1(new_n822), .C2(new_n486), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  NOR2_X1   g400(.A1(G29), .A2(G33), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT90), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G2072), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT93), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n746), .A2(G21), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G168), .B2(new_n746), .ZN(new_n833));
  INV_X1    g408(.A(G1966), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n746), .A2(G20), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT23), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n562), .A2(new_n564), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n559), .B1(new_n560), .B2(new_n519), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n837), .B1(new_n840), .B2(new_n746), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1956), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n829), .B2(new_n828), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n831), .A2(new_n835), .A3(new_n843), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n767), .A2(new_n814), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n763), .A2(new_n845), .ZN(G311));
  INV_X1    g421(.A(G311), .ZN(G150));
  AOI21_X1  g422(.A(new_n621), .B1(new_n608), .B2(new_n614), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n567), .A2(G81), .B1(new_n533), .B2(G43), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n567), .A2(G93), .B1(new_n533), .B2(G55), .ZN(new_n851));
  OAI21_X1  g426(.A(G67), .B1(new_n516), .B2(new_n515), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G651), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n545), .A2(new_n850), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(G55), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n512), .A2(new_n505), .A3(G93), .ZN(new_n858));
  INV_X1    g433(.A(new_n853), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n505), .B2(G67), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n860), .C2(new_n507), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n548), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n849), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n861), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n872));
  INV_X1    g447(.A(new_n629), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n734), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n486), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n485), .A2(G130), .A3(G2105), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n489), .A2(KEYINPUT96), .A3(G130), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n629), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n874), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n874), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n872), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n874), .A2(new_n885), .ZN(new_n889));
  INV_X1    g464(.A(new_n883), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n874), .A2(new_n883), .A3(new_n885), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(KEYINPUT97), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n810), .A2(new_n790), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n788), .A2(new_n787), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n896), .A2(new_n809), .A3(new_n789), .A4(new_n786), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT95), .ZN(new_n899));
  NOR2_X1   g474(.A1(G164), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n501), .A2(new_n503), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n495), .A2(new_n497), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n898), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n503), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n502), .B1(new_n485), .B2(new_n499), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n495), .B(new_n497), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT95), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(new_n903), .A3(new_n895), .A4(new_n897), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n823), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n824), .A2(new_n905), .A3(new_n910), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n894), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n894), .A3(new_n913), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT98), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n912), .A2(new_n894), .A3(new_n913), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n483), .B(new_n636), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G162), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n871), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n912), .A2(new_n913), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT99), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n912), .A2(new_n913), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n886), .A2(new_n887), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n923), .A2(new_n929), .A3(new_n921), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(G395));
  NAND3_X1  g508(.A1(new_n611), .A2(new_n840), .A3(KEYINPUT101), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n606), .A2(G299), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT101), .B1(new_n611), .B2(new_n840), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n606), .B2(G299), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n935), .A4(new_n934), .ZN(new_n942));
  INV_X1    g517(.A(new_n863), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n615), .B2(new_n621), .ZN(new_n944));
  AOI211_X1 g519(.A(G559), .B(new_n863), .C1(new_n608), .C2(new_n614), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n938), .B(new_n942), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n623), .A2(new_n863), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n615), .A2(new_n621), .A3(new_n943), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n940), .A2(new_n935), .A3(new_n934), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  XOR2_X1   g527(.A(G288), .B(KEYINPUT102), .Z(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(new_n582), .ZN(new_n954));
  XNOR2_X1  g529(.A(G303), .B(new_n589), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n946), .A2(new_n950), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n952), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n952), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n861), .A2(new_n591), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(G295));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n963), .ZN(G331));
  NAND4_X1  g540(.A1(new_n850), .A2(new_n851), .A3(new_n545), .A4(new_n855), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n505), .A2(G56), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n507), .B1(new_n967), .B2(new_n543), .ZN(new_n968));
  INV_X1    g543(.A(G81), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n546), .B1(new_n519), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G93), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n857), .B1(new_n519), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n507), .B1(new_n852), .B2(new_n853), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n968), .A2(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n966), .A2(G301), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(G301), .B1(new_n966), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(G286), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(G171), .B1(new_n856), .B2(new_n862), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n966), .A2(G301), .A3(new_n974), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(G168), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n938), .A2(new_n981), .A3(new_n942), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n980), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n949), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT103), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n957), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n982), .A2(new_n987), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n987), .B1(new_n982), .B2(new_n984), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n956), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n992), .A3(new_n871), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  AOI21_X1  g570(.A(G37), .B1(new_n985), .B2(new_n956), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  AND4_X1   g573(.A1(new_n995), .A2(new_n989), .A3(new_n992), .A4(new_n871), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n989), .B2(new_n996), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  MUX2_X1   g576(.A(new_n998), .B(new_n1001), .S(KEYINPUT44), .Z(G397));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n909), .A2(new_n1003), .A3(new_n903), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n471), .A2(new_n477), .A3(new_n482), .A4(G40), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n809), .B(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT105), .ZN(new_n1010));
  INV_X1    g585(.A(G1996), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n790), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n734), .B(new_n736), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G290), .A2(G1986), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1018), .B2(KEYINPUT48), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1018), .A2(KEYINPUT48), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1010), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1008), .B1(new_n1022), .B2(new_n790), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(KEYINPUT46), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(KEYINPUT46), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT47), .Z(new_n1028));
  NAND2_X1  g603(.A1(new_n734), .A2(new_n736), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1013), .A2(new_n1029), .B1(G2067), .B2(new_n809), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1021), .B(new_n1028), .C1(new_n1008), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1007), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n908), .A2(new_n1036), .A3(new_n1003), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT106), .B(G2090), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1005), .A2(G1384), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n909), .A2(new_n903), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n908), .A2(new_n1003), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1005), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1044), .A3(new_n1035), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1039), .A2(new_n1040), .B1(new_n1045), .B2(new_n749), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1033), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT55), .B(G8), .C1(new_n508), .C2(new_n521), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT107), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(KEYINPUT108), .A3(new_n1050), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1045), .A2(new_n749), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1007), .B1(new_n1043), .B2(KEYINPUT50), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1048), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2084), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1034), .A2(new_n1064), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1007), .B1(new_n908), .B2(new_n1041), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1966), .B1(new_n1044), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(G286), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1061), .A2(G8), .A3(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n482), .A2(G40), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n478), .A2(new_n908), .A3(new_n1074), .A4(new_n1003), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n753), .A2(G1976), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(G8), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT109), .B(G1976), .Z(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(G288), .B2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1075), .A2(G8), .A3(new_n1076), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1075), .A2(G8), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT110), .B1(new_n577), .B2(G651), .ZN(new_n1084));
  INV_X1    g659(.A(G1981), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n579), .A2(new_n581), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n578), .A2(KEYINPUT110), .A3(G1981), .A4(new_n580), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(KEYINPUT111), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1088), .B2(KEYINPUT49), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1086), .A2(KEYINPUT111), .A3(new_n1090), .A4(new_n1087), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1082), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1071), .A2(new_n1073), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1032), .B1(new_n1063), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1073), .A2(new_n1092), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1048), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(KEYINPUT114), .A4(new_n1071), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1057), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1069), .A2(G286), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1073), .A3(new_n1099), .A4(new_n1092), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1070), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1094), .B(new_n1097), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(G1976), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1105), .A2(new_n1106), .B1(new_n1085), .B2(new_n582), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1092), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1107), .A2(new_n1083), .B1(new_n1108), .B2(new_n1073), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G286), .A2(G8), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1041), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1035), .B1(G164), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1384), .B1(new_n901), .B2(new_n902), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(KEYINPUT45), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n834), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1116), .B2(new_n1065), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G168), .A2(new_n1047), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1065), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(G8), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1118), .B2(KEYINPUT121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT51), .B1(new_n1111), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(G8), .C1(new_n1119), .C2(G286), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1110), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1069), .A2(new_n1111), .A3(new_n1122), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1117), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n1110), .A2(new_n1128), .A3(new_n1126), .A4(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1098), .A2(new_n1073), .A3(new_n1092), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1961), .B1(new_n1059), .B2(new_n1037), .ZN(new_n1134));
  INV_X1    g709(.A(G2078), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1135), .A2(KEYINPUT53), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1044), .A2(new_n1067), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1133), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1961), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1038), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1044), .A2(new_n1067), .A3(new_n1136), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT123), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1042), .A2(new_n1044), .A3(new_n1135), .A4(new_n1035), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1144));
  AOI22_X1  g719(.A1(new_n1138), .A2(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT125), .B1(new_n1145), .B2(G301), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1134), .A2(new_n1137), .A3(new_n1133), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT123), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(G171), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1132), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1109), .B1(new_n1131), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1104), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G299), .B(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1956), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1038), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(G2072), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1042), .A2(new_n1044), .A3(new_n1035), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1157), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1075), .A2(G2067), .ZN(new_n1164));
  INV_X1    g739(.A(G1348), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1038), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n607), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1159), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1163), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1166), .B1(new_n612), .B2(KEYINPUT60), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1157), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1174), .A2(KEYINPUT61), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(KEYINPUT118), .A3(new_n1168), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT61), .B1(new_n1163), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1007), .A2(G1996), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1042), .A2(new_n1044), .A3(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(KEYINPUT58), .B(G1341), .ZN(new_n1187));
  AOI211_X1 g762(.A(KEYINPUT116), .B(new_n1187), .C1(new_n1035), .C2(new_n1114), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT116), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1187), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n1075), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1186), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT117), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1186), .B(KEYINPUT117), .C1(new_n1188), .C2(new_n1191), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1184), .B1(new_n1196), .B2(new_n549), .ZN(new_n1197));
  AOI211_X1 g772(.A(KEYINPUT59), .B(new_n548), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1179), .B(new_n1183), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1172), .B1(new_n1199), .B2(KEYINPUT120), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n548), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(new_n1184), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n1178), .A2(KEYINPUT61), .A3(new_n1177), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1204), .A2(new_n1174), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1169), .B1(new_n1200), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1132), .B1(new_n1126), .B2(new_n1123), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1140), .A2(KEYINPUT126), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1006), .A2(new_n1042), .A3(new_n1035), .A4(new_n1136), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1140), .A2(KEYINPUT126), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1209), .A2(new_n1147), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1212), .A2(G171), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1213), .B(KEYINPUT54), .C1(G171), .C2(new_n1150), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1208), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g790(.A(new_n1146), .B(new_n1152), .C1(G171), .C2(new_n1212), .ZN(new_n1216));
  XNOR2_X1  g791(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1155), .B1(new_n1207), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1008), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1016), .A2(KEYINPUT104), .ZN(new_n1221));
  NAND2_X1  g796(.A1(G290), .A2(G1986), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1015), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1031), .B1(new_n1219), .B2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  NOR2_X1   g801(.A1(G227), .A2(new_n462), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n718), .B2(new_n719), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1229), .B1(new_n672), .B2(new_n674), .ZN(new_n1230));
  OAI21_X1  g804(.A(new_n1230), .B1(new_n922), .B2(new_n930), .ZN(new_n1231));
  INV_X1    g805(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g806(.A(new_n1227), .B1(new_n998), .B2(new_n1232), .ZN(new_n1233));
  AOI211_X1 g807(.A(KEYINPUT127), .B(new_n1231), .C1(new_n994), .C2(new_n997), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n1233), .A2(new_n1234), .ZN(G308));
  NAND2_X1  g809(.A1(new_n998), .A2(new_n1232), .ZN(G225));
endmodule


