//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  OAI211_X1 g005(.A(KEYINPUT73), .B(new_n202), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n208));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n205), .A2(G113gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n203), .A2(G120gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT1), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT72), .B1(new_n216), .B2(KEYINPUT73), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT74), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n220), .B(new_n210), .C1(new_n213), .C2(new_n217), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n223), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT66), .B(new_n223), .C1(new_n229), .C2(new_n236), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n243), .A2(new_n244), .A3(G183gat), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n226), .A2(new_n228), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT25), .B(new_n241), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n240), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT71), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n249), .A2(KEYINPUT26), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n249), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n250), .A2(new_n251), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  INV_X1    g052(.A(G183gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT27), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n256), .B2(G183gat), .ZN(new_n257));
  OR2_X1    g056(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n258));
  AND4_X1   g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n242), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT28), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(KEYINPUT28), .A3(new_n242), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(KEYINPUT27), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n256), .A2(G183gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n243), .A2(new_n244), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT70), .A4(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n252), .B1(new_n264), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n248), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n222), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n219), .A2(new_n248), .A3(new_n275), .A4(new_n221), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT34), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n280), .B(KEYINPUT64), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n277), .A2(new_n278), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n278), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n221), .A2(new_n219), .B1(new_n248), .B2(new_n275), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n283), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n279), .B2(new_n283), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n298), .A3(KEYINPUT75), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300));
  INV_X1    g099(.A(new_n290), .ZN(new_n301));
  INV_X1    g100(.A(new_n283), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n277), .B2(new_n278), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n303), .B2(KEYINPUT33), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n304), .B2(new_n297), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(KEYINPUT33), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n287), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n282), .A3(new_n285), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n299), .B2(new_n305), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT0), .ZN(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G85gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OR3_X1    g116(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT79), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n320), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n321), .A2(new_n322), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n319), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT80), .B1(new_n330), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT79), .A3(new_n328), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n341), .B1(new_n344), .B2(new_n320), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n218), .ZN(new_n347));
  INV_X1    g146(.A(new_n345), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n342), .A2(new_n343), .B1(new_n319), .B2(new_n318), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n331), .B2(new_n332), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n341), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n345), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n219), .A2(new_n356), .A3(KEYINPUT4), .A4(new_n221), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n218), .A2(new_n348), .A3(new_n351), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n354), .A2(new_n357), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n363));
  INV_X1    g162(.A(new_n217), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n209), .B1(new_n216), .B2(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n210), .C1(new_n340), .C2(new_n345), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n359), .ZN(new_n368));
  INV_X1    g167(.A(new_n358), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n219), .A2(new_n356), .A3(new_n221), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n360), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n359), .A2(new_n360), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n358), .A3(new_n363), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n317), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n370), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n316), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT6), .B(new_n317), .C1(new_n371), .C2(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G197gat), .B(G204gat), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  INV_X1    g190(.A(G218gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(KEYINPUT22), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n389), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n353), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n387), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n397), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n394), .A2(new_n387), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n352), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n348), .A2(new_n351), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n386), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n352), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n386), .B1(new_n406), .B2(new_n403), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n353), .A2(new_n397), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n395), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(G22gat), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT31), .B(G50gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n413), .B1(new_n405), .B2(new_n410), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n405), .A2(new_n410), .ZN(new_n423));
  NAND2_X1  g222(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n411), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n415), .A2(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  INV_X1    g228(.A(G226gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n248), .A2(new_n275), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(KEYINPUT29), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n248), .B2(new_n275), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n395), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n435), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n239), .A2(new_n240), .A3(new_n247), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n250), .A2(new_n251), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n225), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n270), .A2(new_n273), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT28), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n271), .A2(new_n255), .A3(new_n257), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n262), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n438), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n248), .A2(new_n275), .A3(new_n433), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n396), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n437), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n429), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n450), .B2(new_n454), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n437), .A2(new_n449), .A3(new_n429), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n312), .A2(new_n385), .A3(new_n428), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT35), .ZN(new_n460));
  INV_X1    g259(.A(new_n385), .ZN(new_n461));
  INV_X1    g260(.A(new_n458), .ZN(new_n462));
  NOR4_X1   g261(.A1(new_n461), .A2(new_n462), .A3(new_n427), .A4(KEYINPUT35), .ZN(new_n463));
  INV_X1    g262(.A(new_n310), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT75), .B1(new_n295), .B2(new_n298), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n304), .A2(new_n300), .A3(new_n297), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT76), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n311), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n309), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n309), .A2(new_n474), .A3(new_n311), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n306), .A2(new_n308), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n286), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n467), .A2(KEYINPUT76), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n311), .A2(new_n469), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n475), .B1(new_n480), .B2(new_n474), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n385), .A2(new_n427), .A3(new_n458), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n450), .A2(new_n454), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n434), .A2(new_n436), .A3(new_n395), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n396), .B1(new_n447), .B2(new_n448), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT37), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n437), .A2(new_n449), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n488), .A3(new_n454), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n483), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n486), .A2(new_n490), .A3(new_n488), .A4(new_n454), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n492), .A2(new_n383), .A3(new_n384), .A4(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n373), .A2(new_n375), .A3(new_n354), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n369), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n374), .B1(new_n360), .B2(new_n372), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n358), .B1(new_n499), .B2(new_n354), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT39), .B1(new_n368), .B2(new_n369), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n498), .B(new_n316), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT40), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n495), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n317), .B1(new_n500), .B2(new_n497), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n496), .B2(new_n369), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n505), .A2(KEYINPUT84), .A3(new_n507), .A4(KEYINPUT40), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n498), .A2(new_n316), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n510), .B2(new_n506), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n456), .A3(new_n379), .A4(new_n457), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n494), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n482), .B1(new_n513), .B2(new_n428), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n473), .B1(new_n481), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g315(.A1(G43gat), .A2(G50gat), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT86), .B(G43gat), .Z(new_n518));
  OAI211_X1 g317(.A(new_n516), .B(new_n517), .C1(new_n518), .C2(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT14), .B(G29gat), .Z(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(G36gat), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(G43gat), .A2(G50gat), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n516), .B1(new_n525), .B2(new_n517), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n526), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(G1gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  AOI21_X1  g333(.A(G8gat), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n532), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n535), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n527), .A2(new_n528), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n531), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n529), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n540), .B(new_n543), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n545), .B(KEYINPUT13), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G197gat), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT11), .B(G169gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT12), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n546), .A2(new_n547), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n548), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n515), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT91), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(G57gat), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(KEYINPUT90), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(KEYINPUT90), .ZN(new_n576));
  INV_X1    g375(.A(G57gat), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(G64gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n570), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n572), .B(new_n578), .C1(KEYINPUT9), .C2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT92), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(G64gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT9), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n579), .B1(new_n584), .B2(new_n569), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n583), .B(new_n585), .C1(new_n584), .C2(new_n569), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(KEYINPUT8), .A2(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G99gat), .B(G106gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n566), .B1(new_n587), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n587), .A2(new_n596), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n587), .A2(new_n596), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n597), .B1(new_n604), .B2(new_n566), .ZN(new_n605));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n600), .B2(new_n603), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT99), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n608), .B2(KEYINPUT99), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n607), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n608), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n612), .B1(new_n607), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT100), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT10), .B1(new_n600), .B2(new_n603), .ZN(new_n619));
  INV_X1    g418(.A(new_n606), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n619), .A2(new_n620), .A3(new_n597), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n613), .B1(new_n621), .B2(new_n608), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n615), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(G127gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n627), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n626), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G127gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n543), .B1(new_n587), .B2(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n635), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n334), .ZN(new_n640));
  XOR2_X1   g439(.A(G183gat), .B(G211gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n636), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n636), .B2(new_n638), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(KEYINPUT41), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G134gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G162gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n596), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n531), .A2(new_n541), .A3(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n529), .A2(new_n596), .B1(KEYINPUT41), .B2(new_n646), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G190gat), .B(G218gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT93), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n649), .B1(new_n658), .B2(KEYINPUT95), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n653), .A2(new_n655), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT94), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n661), .B(new_n658), .C1(KEYINPUT95), .C2(new_n649), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n625), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n565), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n461), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n462), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G8gat), .B1(new_n669), .B2(new_n458), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n674), .B(new_n676), .S(KEYINPUT42), .Z(G1325gat));
  NAND3_X1  g476(.A1(new_n477), .A2(KEYINPUT36), .A3(new_n467), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n471), .B2(KEYINPUT36), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n480), .A2(G15gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n669), .B2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n670), .A2(new_n427), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT101), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n481), .A2(new_n514), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n513), .A2(new_n428), .ZN(new_n689));
  INV_X1    g488(.A(new_n482), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT102), .B1(new_n691), .B2(new_n679), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n473), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n459), .A2(KEYINPUT35), .B1(new_n463), .B2(new_n471), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n687), .B1(new_n481), .B2(new_n514), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n691), .A2(new_n679), .A3(KEYINPUT102), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT103), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n666), .A2(KEYINPUT44), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n695), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n515), .A2(new_n665), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT44), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n564), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n625), .A2(new_n645), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT104), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  INV_X1    g508(.A(new_n707), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n709), .B(new_n710), .C1(new_n702), .C2(new_n704), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n385), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n515), .A2(new_n665), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n707), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(G29gat), .A3(new_n385), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT45), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(G1328gat));
  OAI21_X1  g518(.A(G36gat), .B1(new_n713), .B2(new_n458), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n716), .A2(G36gat), .A3(new_n458), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(new_n518), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n715), .A2(new_n707), .A3(new_n471), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT105), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n703), .A2(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n697), .A2(new_n698), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT103), .B1(new_n730), .B2(new_n473), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n694), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n729), .B1(new_n733), .B2(new_n701), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n709), .B1(new_n734), .B2(new_n710), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n710), .B1(new_n702), .B2(new_n704), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n481), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n728), .B1(new_n738), .B2(new_n518), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n724), .B1(new_n736), .B2(new_n481), .ZN(new_n740));
  INV_X1    g539(.A(new_n725), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT47), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT106), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n724), .B1(new_n712), .B2(new_n481), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n745), .B(new_n742), .C1(new_n746), .C2(new_n728), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1330gat));
  NOR2_X1   g547(.A1(new_n625), .A2(new_n645), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n428), .A2(G50gat), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n666), .B1(KEYINPUT107), .B2(new_n750), .ZN(new_n752));
  AND4_X1   g551(.A1(new_n565), .A2(new_n749), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n712), .A2(new_n427), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  INV_X1    g554(.A(G50gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n736), .B2(new_n427), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n755), .A2(KEYINPUT48), .B1(new_n757), .B2(new_n759), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n695), .A2(new_n700), .ZN(new_n761));
  INV_X1    g560(.A(new_n667), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n706), .A3(new_n625), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n461), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n462), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  INV_X1    g569(.A(new_n764), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n567), .B1(new_n771), .B2(new_n480), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n481), .A2(G71gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n771), .A2(KEYINPUT108), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  INV_X1    g574(.A(new_n773), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n764), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n427), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n643), .A2(new_n644), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(KEYINPUT109), .A3(new_n706), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT109), .B1(new_n782), .B2(new_n706), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n665), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n786), .A2(new_n787), .A3(new_n699), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n786), .B2(new_n699), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n591), .A3(new_n461), .A4(new_n625), .ZN(new_n792));
  INV_X1    g591(.A(new_n615), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n617), .A2(KEYINPUT100), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n622), .A2(new_n623), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n785), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n783), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n705), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n385), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n800), .ZN(G1336gat));
  NAND2_X1  g600(.A1(new_n625), .A2(new_n462), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  INV_X1    g602(.A(new_n790), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n788), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n799), .A2(new_n458), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n592), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n809), .B2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n799), .B2(new_n679), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n796), .A2(G99gat), .A3(new_n480), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n791), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1338gat));
  NOR2_X1   g618(.A1(new_n799), .A2(new_n428), .ZN(new_n820));
  INV_X1    g619(.A(G106gat), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT113), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n796), .A2(G106gat), .A3(new_n428), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n791), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n820), .B2(new_n821), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n822), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n822), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(G1339gat));
  OAI21_X1  g629(.A(new_n620), .B1(new_n619), .B2(new_n597), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n607), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n612), .B1(new_n621), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n832), .B2(new_n834), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n558), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n561), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n549), .A2(new_n551), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT114), .Z(new_n842));
  AOI21_X1  g641(.A(new_n545), .B1(new_n542), .B2(new_n544), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n557), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n665), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n663), .A2(new_n562), .A3(new_n563), .A4(new_n664), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n615), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n665), .A2(new_n845), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n838), .A2(new_n848), .B1(new_n796), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n851), .A2(new_n782), .B1(new_n668), .B2(new_n706), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n427), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n462), .A2(new_n385), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n471), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n203), .A3(new_n706), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n762), .A2(new_n706), .A3(new_n796), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n846), .A2(new_n615), .A3(new_n847), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n832), .A2(new_n834), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT55), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n858), .A2(new_n862), .B1(new_n625), .B2(new_n849), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n857), .B1(new_n863), .B2(new_n645), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n312), .A2(new_n428), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n462), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n461), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n564), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n856), .A2(new_n869), .ZN(G1340gat));
  AOI21_X1  g669(.A(G120gat), .B1(new_n868), .B2(new_n625), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n854), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n796), .A2(new_n205), .A3(new_n480), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n855), .B2(new_n782), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n632), .A3(new_n645), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1342gat));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n666), .A2(G134gat), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n867), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n879), .B1(new_n867), .B2(new_n880), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n855), .B2(new_n666), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n883), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(KEYINPUT56), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT116), .B(new_n882), .C1(new_n881), .C2(new_n883), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n679), .A2(new_n854), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n852), .B2(new_n428), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n427), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n325), .B1(new_n896), .B2(new_n564), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n481), .A2(new_n428), .ZN(new_n900));
  AND4_X1   g699(.A1(new_n461), .A2(new_n864), .A3(new_n458), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n325), .A3(new_n564), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n902), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT58), .B1(new_n897), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1344gat));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n326), .A3(new_n625), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  INV_X1    g707(.A(new_n892), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n796), .B1(KEYINPUT117), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(KEYINPUT117), .B2(new_n909), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n894), .B2(new_n895), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n326), .B1(new_n912), .B2(KEYINPUT118), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n326), .C1(new_n896), .C2(new_n625), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(new_n334), .B1(new_n896), .B2(new_n645), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n901), .A2(new_n334), .A3(new_n645), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  AOI21_X1  g719(.A(G162gat), .B1(new_n901), .B2(new_n665), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n666), .A2(new_n335), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n896), .B2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n461), .A2(new_n458), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n471), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n853), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n230), .A3(new_n706), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n852), .A2(new_n461), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n865), .A2(new_n458), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n564), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n928), .B1(new_n230), .B2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(new_n231), .B1(new_n931), .B2(new_n796), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n796), .A2(new_n231), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n927), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n853), .A2(KEYINPUT119), .A3(new_n926), .A4(new_n937), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(G1349gat));
  NAND3_X1  g742(.A1(new_n932), .A2(new_n272), .A3(new_n645), .ZN(new_n944));
  OAI21_X1  g743(.A(G183gat), .B1(new_n927), .B2(new_n782), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1350gat));
  INV_X1    g750(.A(new_n271), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n931), .A2(new_n952), .A3(new_n666), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT122), .ZN(new_n954));
  OAI21_X1  g753(.A(G190gat), .B1(new_n927), .B2(new_n666), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1351gat));
  NAND2_X1  g756(.A1(new_n894), .A2(new_n895), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n679), .A2(new_n924), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT124), .Z(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n706), .ZN(new_n962));
  XOR2_X1   g761(.A(KEYINPUT123), .B(G197gat), .Z(new_n963));
  NAND3_X1  g762(.A1(new_n929), .A2(new_n462), .A3(new_n900), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n564), .A2(new_n963), .ZN(new_n965));
  OAI22_X1  g764(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  NOR2_X1   g765(.A1(new_n802), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n929), .A2(new_n900), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT125), .ZN(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n961), .B2(new_n796), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n970), .B(new_n971), .C1(KEYINPUT62), .C2(new_n968), .ZN(G1353gat));
  NOR2_X1   g771(.A1(new_n782), .A2(new_n959), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G211gat), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT63), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(KEYINPUT63), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n645), .A2(new_n391), .ZN(new_n979));
  OR3_X1    g778(.A1(new_n964), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n978), .B1(new_n964), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n976), .A2(new_n977), .A3(new_n982), .ZN(G1354gat));
  NOR3_X1   g782(.A1(new_n961), .A2(new_n392), .A3(new_n666), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n392), .B1(new_n964), .B2(new_n666), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1355gat));
endmodule


