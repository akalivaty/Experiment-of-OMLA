//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT11), .A2(G134), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT11), .A2(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT68), .B(G131), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT67), .B(G137), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n190), .B(new_n191), .C1(new_n192), .C2(new_n188), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT69), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT67), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n188), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(new_n191), .A4(new_n190), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n194), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n196), .A2(new_n198), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT70), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n205), .B2(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n195), .A2(KEYINPUT70), .A3(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(KEYINPUT1), .A3(G146), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(new_n219), .C1(G128), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n211), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n187), .B1(new_n204), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n194), .A2(new_n203), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n201), .A2(new_n190), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n215), .A2(new_n217), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n230), .A2(new_n231), .B1(new_n215), .B2(new_n217), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n234), .ZN(new_n239));
  INV_X1    g053(.A(new_n228), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n236), .A2(new_n239), .B1(new_n220), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n227), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n211), .A2(new_n221), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n224), .A3(KEYINPUT71), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n223), .A2(new_n242), .A3(KEYINPUT30), .A4(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n251), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n194), .A2(new_n203), .B1(G131), .B2(new_n225), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n220), .A2(new_n240), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n238), .B1(new_n237), .B2(new_n234), .ZN(new_n258));
  AND4_X1   g072(.A1(new_n238), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n222), .B1(new_n203), .B2(new_n194), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n245), .A2(new_n254), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT72), .B(G953), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G237), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n254), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n223), .A2(new_n242), .A3(new_n273), .A4(new_n244), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n264), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n243), .A2(new_n224), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n242), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n280), .C1(new_n278), .C2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n275), .B1(new_n282), .B2(new_n272), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n223), .A2(new_n242), .A3(new_n244), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n254), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n274), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT29), .A3(new_n271), .A4(new_n279), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n291), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n264), .A2(new_n271), .A3(new_n274), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n281), .A2(new_n272), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n264), .A2(new_n299), .A3(new_n271), .A4(new_n274), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n301), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT32), .B1(new_n301), .B2(new_n302), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(KEYINPUT74), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n295), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n241), .A2(G125), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n221), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G224), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G953), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT90), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n312), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G122), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n318));
  OAI21_X1  g132(.A(G113), .B1(new_n247), .B2(KEYINPUT5), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n252), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G107), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G104), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  INV_X1    g137(.A(G104), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G107), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(KEYINPUT3), .A3(G104), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G101), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT85), .B1(new_n321), .B2(G104), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n324), .A3(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(G104), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G101), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n320), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n327), .B2(new_n328), .ZN(new_n339));
  INV_X1    g153(.A(new_n322), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n321), .A2(KEYINPUT3), .A3(G104), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT3), .B1(new_n321), .B2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G101), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n338), .A3(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n254), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n317), .B1(new_n337), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n337), .A2(new_n347), .A3(new_n317), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(KEYINPUT89), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n348), .B2(new_n352), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n316), .B(new_n351), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n320), .A2(new_n336), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n319), .B(KEYINPUT92), .Z(new_n359));
  OAI21_X1  g173(.A(new_n252), .B1(new_n359), .B2(new_n318), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n360), .B2(new_n336), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n317), .B(KEYINPUT91), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT8), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n314), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n309), .A2(new_n366), .A3(new_n311), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n309), .B2(new_n311), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n364), .B(new_n350), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n357), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G210), .B1(G237), .B2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n357), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G140), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT83), .ZN(new_n381));
  INV_X1    g195(.A(G953), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT72), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G953), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n386), .A2(G227), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n381), .B(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n224), .A2(KEYINPUT86), .A3(new_n226), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT86), .B1(new_n224), .B2(new_n226), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n236), .A2(new_n239), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n392), .A2(new_n345), .A3(new_n257), .A4(new_n346), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n221), .A2(new_n329), .A3(new_n335), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT10), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n221), .A2(new_n329), .A3(new_n335), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT10), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n388), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n221), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n336), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n396), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n227), .A3(KEYINPUT12), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT12), .B1(new_n403), .B2(new_n227), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n393), .A2(new_n398), .A3(new_n395), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n227), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n256), .A2(KEYINPUT86), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n399), .A2(new_n227), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n388), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n379), .B(new_n370), .C1(new_n408), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT87), .ZN(new_n418));
  INV_X1    g232(.A(new_n388), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n391), .A2(new_n399), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n399), .A2(new_n227), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n221), .B1(new_n329), .B2(new_n335), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n394), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n425), .B2(new_n256), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n404), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n427), .A3(new_n388), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n379), .A4(new_n370), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n418), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n388), .A2(KEYINPUT84), .ZN(new_n435));
  AOI211_X1 g249(.A(new_n434), .B(new_n435), .C1(new_n414), .C2(new_n427), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n414), .A2(new_n388), .A3(new_n415), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n370), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G469), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G221), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT9), .B(G234), .Z(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n370), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(KEYINPUT88), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n418), .A2(new_n431), .B1(new_n439), .B2(G469), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(new_n444), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n378), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G217), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(G234), .B2(new_n370), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n246), .A2(G128), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n454), .A2(KEYINPUT23), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n246), .A2(G128), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(KEYINPUT23), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n454), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n459), .A2(new_n456), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT24), .B(G110), .Z(new_n461));
  OAI22_X1  g275(.A1(new_n458), .A2(G110), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT16), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n310), .A2(KEYINPUT77), .A3(G140), .ZN(new_n467));
  XNOR2_X1  g281(.A(G125), .B(G140), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT77), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n471));
  OAI211_X1 g285(.A(G146), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n216), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n460), .A2(new_n461), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n310), .A2(G140), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n464), .A3(new_n469), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n310), .A2(KEYINPUT77), .A3(G140), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n465), .B1(new_n482), .B2(KEYINPUT16), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n478), .B1(new_n483), .B2(G146), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT79), .B(new_n216), .C1(new_n485), .C2(new_n465), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n472), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(KEYINPUT78), .A3(G146), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n477), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT76), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n458), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n458), .A2(new_n493), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(G110), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n475), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT82), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n442), .B1(new_n383), .B2(new_n385), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n499), .A2(new_n500), .A3(G234), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n499), .B2(G234), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT22), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n386), .A2(G221), .A3(G234), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT80), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT22), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n500), .A3(G234), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n503), .A2(G137), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(G137), .B1(new_n503), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n497), .A2(new_n498), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT22), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n195), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n503), .A2(G137), .A3(new_n508), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT81), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT79), .B1(new_n521), .B2(new_n216), .ZN(new_n522));
  INV_X1    g336(.A(new_n486), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT78), .B1(new_n483), .B2(G146), .ZN(new_n524));
  NOR4_X1   g338(.A1(new_n485), .A2(new_n488), .A3(new_n216), .A4(new_n465), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n496), .A3(new_n476), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n474), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT82), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n527), .A2(new_n474), .A3(new_n511), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n370), .B(new_n512), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND4_X1   g347(.A1(new_n498), .A2(new_n527), .A3(new_n474), .A4(new_n511), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n517), .A2(KEYINPUT81), .A3(new_n518), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n498), .B1(new_n497), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n497), .A2(new_n511), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT25), .A3(new_n370), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n453), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n452), .A2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G116), .B(G122), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n321), .ZN(new_n551));
  INV_X1    g365(.A(G122), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(new_n552), .B2(G116), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(new_n554), .B1(G116), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n554), .B2(new_n553), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n552), .A2(KEYINPUT14), .A3(G116), .ZN(new_n557));
  OAI21_X1  g371(.A(G107), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G128), .B(G143), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT95), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n205), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n205), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n551), .B(new_n558), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n550), .B(new_n321), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n212), .A2(G143), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n212), .A2(G143), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(KEYINPUT13), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(KEYINPUT13), .B2(new_n567), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n561), .B(new_n565), .C1(new_n569), .C2(new_n205), .ZN(new_n570));
  INV_X1    g384(.A(new_n443), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n571), .A2(new_n451), .A3(G953), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n564), .B2(new_n570), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n370), .B(new_n549), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n570), .ZN(new_n578));
  INV_X1    g392(.A(new_n572), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n573), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n549), .B1(new_n581), .B2(new_n370), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n191), .ZN(new_n584));
  AOI21_X1  g398(.A(G143), .B1(new_n266), .B2(G214), .ZN(new_n585));
  INV_X1    g399(.A(G237), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n386), .A2(G214), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n214), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n214), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n191), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT17), .A3(new_n584), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n594), .A2(new_n487), .A3(new_n491), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(KEYINPUT18), .A3(G131), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n473), .B1(new_n482), .B2(new_n216), .ZN(new_n599));
  NAND2_X1  g413(.A1(KEYINPUT18), .A2(G131), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n591), .A2(new_n592), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(G113), .B(G122), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT93), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(new_n324), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n597), .B2(new_n602), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n370), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT94), .B(G475), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n605), .ZN(new_n612));
  INV_X1    g426(.A(new_n602), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT19), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n468), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n482), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n472), .B1(G146), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n589), .B2(new_n593), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n612), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(G475), .B1(new_n606), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT20), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(new_n370), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n620), .B2(new_n370), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n583), .B(new_n611), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(G952), .ZN(new_n626));
  AOI211_X1 g440(.A(G953), .B(new_n626), .C1(G234), .C2(G237), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n370), .B(new_n386), .C1(G234), .C2(G237), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT21), .B(G898), .Z(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT97), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n606), .A2(new_n619), .ZN(new_n633));
  INV_X1    g447(.A(G475), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n370), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT20), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n636), .A2(new_n622), .B1(new_n609), .B2(new_n610), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n638));
  INV_X1    g452(.A(new_n631), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n583), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n308), .A2(new_n450), .A3(new_n546), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  NAND2_X1  g457(.A1(new_n446), .A2(new_n449), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n301), .A2(new_n370), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n301), .A2(new_n302), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n376), .A2(new_n639), .A3(new_n377), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n650), .A3(new_n546), .ZN(new_n651));
  INV_X1    g465(.A(new_n637), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n574), .A2(new_n575), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT33), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n581), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n654), .A2(new_n656), .A3(G478), .A4(new_n370), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n547), .B1(new_n653), .B2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT34), .B(G104), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  OR2_X1    g477(.A1(new_n577), .A2(new_n582), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n637), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n651), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT35), .B(G107), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR2_X1   g482(.A1(new_n531), .A2(new_n532), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT25), .B1(new_n540), .B2(new_n370), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n452), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n497), .B(KEYINPUT98), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n543), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n671), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n543), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n528), .B(KEYINPUT98), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(KEYINPUT36), .B2(new_n520), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n680), .B1(new_n682), .B2(new_n675), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT99), .B1(new_n542), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n648), .B1(new_n640), .B2(new_n632), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n450), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT100), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT37), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(G110), .Z(G12));
  INV_X1    g504(.A(new_n628), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n691), .A2(KEYINPUT101), .A3(G900), .ZN(new_n692));
  INV_X1    g506(.A(new_n627), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT101), .B1(new_n691), .B2(G900), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n665), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n308), .A2(new_n450), .A3(new_n685), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XNOR2_X1  g513(.A(new_n376), .B(KEYINPUT102), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n671), .A2(new_n664), .A3(new_n652), .A4(new_n678), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT32), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n647), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT74), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n301), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n306), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n370), .B1(new_n288), .B2(new_n271), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n264), .A2(new_n274), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n271), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n709), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n702), .B1(new_n708), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n701), .A2(new_n377), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n695), .B(KEYINPUT39), .Z(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n644), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT40), .Z(new_n724));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  INV_X1    g540(.A(new_n659), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n637), .A3(new_n696), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n308), .A2(new_n450), .A3(new_n685), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  NAND2_X1  g544(.A1(new_n429), .A2(new_n370), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n432), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n444), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n660), .A2(new_n649), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n308), .A2(new_n546), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT41), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G113), .ZN(G15));
  INV_X1    g552(.A(new_n649), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n308), .A2(new_n546), .A3(new_n739), .A4(new_n734), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n665), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n248), .ZN(G18));
  NOR3_X1   g556(.A1(new_n378), .A2(new_n733), .A3(new_n444), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n308), .A2(new_n685), .A3(new_n641), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  AND2_X1   g559(.A1(new_n289), .A2(new_n279), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n297), .B(new_n300), .C1(new_n746), .C2(new_n271), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT104), .B(G472), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n747), .A2(new_n302), .B1(new_n645), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n546), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n378), .A2(new_n583), .A3(new_n637), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n639), .A3(new_n734), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NAND2_X1  g567(.A1(new_n671), .A2(new_n678), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n749), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n728), .A3(new_n743), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  XNOR2_X1  g571(.A(new_n290), .B(KEYINPUT75), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n709), .B1(new_n758), .B2(new_n285), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n704), .A2(new_n706), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n546), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n374), .A2(new_n377), .A3(new_n375), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n728), .A2(new_n445), .A3(new_n441), .A4(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT42), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n696), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n441), .A2(new_n445), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n762), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n308), .A2(new_n546), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(G131), .Z(G33));
  AND4_X1   g585(.A1(new_n308), .A2(new_n546), .A3(new_n697), .A4(new_n768), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT105), .B(G134), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G36));
  NAND2_X1  g588(.A1(new_n637), .A2(new_n659), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT43), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n754), .A2(new_n648), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT44), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n779), .A2(KEYINPUT107), .A3(new_n763), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT107), .B1(new_n779), .B2(new_n763), .ZN(new_n781));
  OAI22_X1  g595(.A1(new_n780), .A2(new_n781), .B1(KEYINPUT44), .B2(new_n778), .ZN(new_n782));
  INV_X1    g596(.A(new_n434), .ZN(new_n783));
  INV_X1    g597(.A(new_n435), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n783), .B(new_n784), .C1(new_n407), .C2(new_n420), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n437), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT45), .ZN(new_n787));
  OAI21_X1  g601(.A(G469), .B1(new_n787), .B2(G902), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n432), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(KEYINPUT106), .A3(new_n432), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n792), .B(new_n793), .C1(KEYINPUT46), .C2(new_n788), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n445), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n782), .A2(new_n721), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT108), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND2_X1  g612(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n308), .A2(new_n546), .A3(new_n660), .A4(new_n696), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n801), .A3(new_n445), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n799), .A2(new_n763), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  XNOR2_X1  g621(.A(new_n664), .B(KEYINPUT110), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n660), .B1(new_n808), .B2(new_n652), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n644), .A2(new_n809), .A3(new_n650), .A4(new_n546), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n308), .A2(new_n546), .ZN(new_n811));
  INV_X1    g625(.A(new_n378), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n644), .A2(new_n641), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n687), .B(new_n810), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT111), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n642), .A2(new_n816), .A3(new_n687), .A4(new_n810), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n736), .A2(new_n744), .A3(new_n752), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n741), .A3(new_n770), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n308), .A2(new_n685), .A3(new_n808), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n644), .A2(new_n637), .A3(new_n695), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n755), .A2(new_n728), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n767), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n772), .B1(new_n824), .B2(new_n763), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n818), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT112), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n698), .A2(new_n729), .A3(new_n756), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  INV_X1    g643(.A(new_n377), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n830), .B(new_n696), .C1(new_n374), .C2(new_n375), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n445), .A3(new_n441), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n829), .B1(new_n716), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n714), .B1(new_n707), .B2(new_n306), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n835), .A2(new_n832), .A3(new_n702), .A4(KEYINPUT113), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n828), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n715), .B1(new_n305), .B2(new_n307), .ZN(new_n840));
  INV_X1    g654(.A(new_n702), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n833), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT113), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n716), .A2(new_n829), .A3(new_n833), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n698), .A2(new_n729), .A3(new_n756), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT52), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n818), .A2(new_n820), .A3(new_n849), .A4(new_n825), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n827), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n818), .A2(new_n820), .A3(new_n825), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n848), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n854), .B(new_n856), .C1(new_n852), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n818), .A2(new_n862), .A3(new_n825), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n839), .A2(new_n847), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT53), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n826), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n861), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n818), .A2(new_n862), .A3(new_n825), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n848), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n874), .A3(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(KEYINPUT116), .A3(new_n861), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n776), .A2(new_n693), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n734), .A3(new_n750), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n701), .A3(new_n377), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT50), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n733), .A2(new_n762), .A3(new_n444), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT119), .Z(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n755), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n835), .A2(new_n883), .A3(new_n546), .A4(new_n627), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n887), .A2(new_n652), .A3(new_n659), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n882), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n733), .B(KEYINPUT118), .Z(new_n890));
  AOI22_X1  g704(.A1(new_n799), .A2(new_n802), .B1(new_n444), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n879), .A2(new_n750), .A3(new_n763), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT117), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(KEYINPUT51), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n889), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n626), .A2(G953), .ZN(new_n899));
  OAI221_X1 g713(.A(new_n899), .B1(new_n660), .B2(new_n887), .C1(new_n880), .C2(new_n378), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT48), .ZN(new_n903));
  INV_X1    g717(.A(new_n761), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n885), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n901), .B2(new_n900), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n896), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n860), .A2(new_n878), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n905), .A2(new_n903), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n909), .A2(new_n910), .B1(G952), .B2(G953), .ZN(new_n911));
  INV_X1    g725(.A(new_n546), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n701), .A2(new_n912), .A3(new_n830), .A4(new_n444), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n733), .A2(KEYINPUT49), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n775), .B1(new_n733), .B2(KEYINPUT49), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n913), .A2(new_n835), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n876), .A2(new_n370), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT56), .B1(new_n918), .B2(G210), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n351), .B1(new_n354), .B2(new_n356), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n316), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n919), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n265), .A2(new_n626), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT121), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n923), .A2(new_n926), .ZN(G51));
  NAND2_X1  g741(.A1(G469), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT57), .Z(new_n929));
  INV_X1    g743(.A(new_n870), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n876), .A2(new_n861), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n429), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n918), .A2(G469), .A3(new_n787), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(G54));
  INV_X1    g749(.A(KEYINPUT58), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n876), .A2(new_n936), .A3(new_n370), .ZN(new_n937));
  AND4_X1   g751(.A1(G475), .A2(new_n937), .A3(new_n619), .A4(new_n606), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n937), .A2(G475), .B1(new_n619), .B2(new_n606), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n925), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n925), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(G60));
  AND2_X1   g758(.A1(new_n654), .A2(new_n656), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n851), .A2(new_n855), .A3(new_n852), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n855), .B1(new_n851), .B2(new_n852), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n858), .A2(new_n852), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT116), .B1(new_n876), .B2(new_n861), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n871), .B(KEYINPUT54), .C1(new_n875), .C2(new_n867), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n949), .A2(new_n861), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n945), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n945), .B(new_n955), .C1(new_n930), .C2(new_n931), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n925), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT123), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n868), .A2(new_n869), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT54), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n954), .B1(new_n962), .B2(new_n870), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n926), .B1(new_n963), .B2(new_n945), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n954), .B1(new_n860), .B2(new_n878), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n960), .B(new_n964), .C1(new_n965), .C2(new_n945), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n959), .A2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT60), .Z(new_n969));
  OAI211_X1 g783(.A(new_n961), .B(new_n969), .C1(new_n676), .C2(new_n677), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n961), .A2(new_n969), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n970), .B(new_n925), .C1(new_n971), .C2(new_n540), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n630), .B2(new_n313), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n819), .A2(new_n741), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n818), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n974), .B1(new_n977), .B2(new_n265), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n920), .B1(G898), .B2(new_n386), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  NAND2_X1  g795(.A1(new_n904), .A2(new_n751), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n795), .A2(new_n721), .A3(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n796), .A2(new_n983), .A3(new_n772), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n846), .A2(new_n770), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n806), .A2(new_n984), .A3(new_n386), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n245), .A2(new_n263), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(new_n616), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n265), .A2(G900), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n725), .A2(new_n828), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n725), .A2(KEYINPUT62), .A3(new_n828), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n796), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n809), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n811), .A2(new_n723), .A3(new_n996), .A4(new_n762), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n804), .B2(new_n805), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n265), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n990), .B1(new_n999), .B2(new_n988), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT125), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n990), .B(new_n1002), .C1(new_n999), .C2(new_n988), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n386), .B1(G227), .B2(G900), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  NAND3_X1  g822(.A1(new_n806), .A2(new_n984), .A3(new_n985), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(new_n976), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n275), .B(KEYINPUT126), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n926), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n995), .A2(new_n998), .A3(new_n977), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n713), .B1(new_n1014), .B2(new_n1008), .ZN(new_n1015));
  AND4_X1   g829(.A1(new_n275), .A2(new_n859), .A3(new_n713), .A4(new_n1008), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(G57));
endmodule


