//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G29gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n217), .A3(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(new_n212), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(new_n214), .B2(new_n215), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n224), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n213), .A2(new_n217), .A3(KEYINPUT15), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT88), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(KEYINPUT88), .A3(G1gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n229), .A2(new_n234), .B1(KEYINPUT89), .B2(G8gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n237));
  INV_X1    g036(.A(G8gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n232), .A2(new_n240), .A3(new_n233), .A4(new_n235), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n228), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n241), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(KEYINPUT90), .A3(new_n241), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n228), .A2(KEYINPUT17), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(new_n225), .B2(new_n227), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n208), .B(new_n242), .C1(new_n247), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT91), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n242), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n239), .A2(KEYINPUT90), .A3(new_n241), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT90), .B1(new_n239), .B2(new_n241), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n228), .B(KEYINPUT17), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT18), .A4(new_n208), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n208), .B(KEYINPUT13), .Z(new_n264));
  AND2_X1   g063(.A1(new_n225), .A2(new_n227), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n243), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT92), .A3(new_n242), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n243), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n264), .A2(new_n270), .B1(new_n252), .B2(new_n253), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n207), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT86), .B(new_n206), .C1(new_n263), .C2(new_n271), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278));
  INV_X1    g077(.A(G155gat), .ZN(new_n279));
  INV_X1    g078(.A(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT72), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G162gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(G162gat), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT73), .B(KEYINPUT2), .C1(new_n287), .C2(new_n279), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n280), .A2(G155gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n279), .A2(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n286), .A2(new_n288), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n293), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n291), .A2(new_n294), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT2), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  INV_X1    g101(.A(G127gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G134gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(KEYINPUT1), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G113gat), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n300), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n297), .A2(KEYINPUT4), .A3(new_n316), .A4(new_n300), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n297), .B2(new_n300), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n307), .A2(new_n315), .A3(KEYINPUT74), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT74), .B1(new_n307), .B2(new_n315), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n300), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT2), .B1(new_n287), .B2(new_n279), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n295), .B1(new_n330), .B2(new_n278), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n288), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n323), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n322), .A2(new_n334), .A3(KEYINPUT5), .A4(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT75), .B1(new_n327), .B2(new_n332), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n307), .A2(new_n315), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n307), .A2(new_n315), .A3(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n297), .A2(new_n300), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n317), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n335), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n337), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n297), .A2(new_n323), .A3(new_n300), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n350), .A2(new_n324), .A3(new_n327), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n351), .A2(new_n321), .A3(new_n348), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n336), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n359));
  INV_X1    g158(.A(new_n357), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n336), .C1(new_n349), .C2(new_n352), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT76), .B1(new_n363), .B2(KEYINPUT6), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n361), .A2(new_n365), .A3(new_n359), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT64), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n372), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n371), .A2(new_n373), .A3(new_n376), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT23), .ZN(new_n382));
  INV_X1    g181(.A(G169gat), .ZN(new_n383));
  INV_X1    g182(.A(G176gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n383), .A2(KEYINPUT23), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT65), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G176gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  OR3_X1    g192(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n394), .A2(new_n376), .A3(new_n370), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(KEYINPUT23), .B2(new_n381), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT23), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT25), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n392), .A2(new_n393), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT26), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n403), .A3(new_n381), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(KEYINPUT26), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n374), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT28), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT67), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT27), .B(G183gat), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n378), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n378), .A3(new_n408), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT69), .B1(new_n402), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n404), .A2(new_n374), .A3(new_n405), .ZN(new_n415));
  INV_X1    g214(.A(new_n412), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(new_n410), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT69), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n401), .A2(new_n396), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT65), .B(G176gat), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n420), .A2(new_n387), .B1(new_n382), .B2(new_n385), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT25), .B1(new_n421), .B2(new_n380), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n417), .B(new_n418), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n369), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G197gat), .B(G204gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT22), .ZN(new_n428));
  INV_X1    g227(.A(G211gat), .ZN(new_n429));
  INV_X1    g228(.A(G218gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G211gat), .B(G218gat), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n417), .B1(new_n419), .B2(new_n422), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n369), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT70), .B1(new_n426), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n425), .A3(new_n368), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n439), .B(new_n444), .C1(new_n424), .C2(new_n368), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT70), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT29), .B1(new_n414), .B2(new_n423), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n441), .C1(new_n447), .C2(new_n369), .ZN(new_n448));
  XNOR2_X1  g247(.A(G8gat), .B(G36gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  NAND4_X1  g250(.A1(new_n443), .A2(new_n445), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n448), .A2(new_n445), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(KEYINPUT71), .A3(new_n443), .A4(new_n451), .ZN(new_n456));
  INV_X1    g255(.A(new_n451), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n443), .A2(new_n445), .A3(new_n448), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(KEYINPUT37), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n440), .A2(new_n369), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n426), .A2(new_n438), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n444), .B1(new_n424), .B2(new_n368), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT37), .B1(new_n463), .B2(new_n439), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n454), .B(new_n456), .C1(new_n459), .C2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT85), .B1(new_n367), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n365), .B1(new_n361), .B2(new_n359), .ZN(new_n468));
  NOR4_X1   g267(.A1(new_n351), .A2(new_n321), .A3(new_n337), .A4(new_n348), .ZN(new_n469));
  INV_X1    g268(.A(new_n352), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n346), .A2(new_n317), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n345), .B1(new_n343), .B2(new_n344), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n348), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(new_n360), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n361), .A2(new_n359), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n468), .A2(new_n476), .B1(new_n477), .B2(new_n358), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n459), .A2(new_n465), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n454), .A2(new_n456), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n458), .A2(KEYINPUT37), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT38), .B1(new_n483), .B2(new_n459), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n438), .B1(new_n333), .B2(new_n425), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n438), .A2(new_n425), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n332), .B1(new_n487), .B2(new_n323), .ZN(new_n488));
  OAI211_X1 g287(.A(G228gat), .B(G233gat), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n425), .B1(new_n344), .B2(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n439), .ZN(new_n491));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n433), .A2(KEYINPUT78), .A3(new_n435), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n437), .A2(KEYINPUT79), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n432), .A2(new_n495), .A3(new_n434), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT78), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n432), .B2(new_n434), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n494), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT3), .B1(new_n499), .B2(new_n425), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n491), .B(new_n492), .C1(new_n332), .C2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G22gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n489), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n489), .B2(new_n501), .ZN(new_n505));
  XNOR2_X1  g304(.A(G78gat), .B(G106gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G50gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT80), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(KEYINPUT80), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n504), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n489), .A2(new_n501), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G22gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n511), .B1(new_n516), .B2(new_n503), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n348), .B1(new_n351), .B2(new_n321), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n520));
  OAI21_X1  g319(.A(new_n357), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n338), .A2(new_n335), .A3(new_n317), .A4(new_n346), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n519), .A2(KEYINPUT39), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n361), .B1(new_n526), .B2(KEYINPUT40), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(KEYINPUT40), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(KEYINPUT84), .A3(KEYINPUT40), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n455), .A2(KEYINPUT30), .A3(new_n443), .A4(new_n451), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n458), .A2(new_n457), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n454), .A2(new_n456), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n518), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n485), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n518), .B1(new_n538), .B2(new_n478), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT81), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n440), .A2(new_n339), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n417), .B(new_n316), .C1(new_n419), .C2(new_n422), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G227gat), .ZN(new_n549));
  INV_X1    g348(.A(G233gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n545), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G43gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(G71gat), .B(G99gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT34), .B1(new_n548), .B2(new_n551), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT34), .ZN(new_n558));
  INV_X1    g357(.A(new_n551), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n546), .A2(new_n558), .A3(new_n559), .A4(new_n547), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n548), .A2(new_n551), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT32), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n557), .B(new_n560), .C1(new_n552), .C2(new_n555), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n562), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n543), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n562), .A2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n564), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT36), .A3(new_n567), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n541), .A2(new_n542), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n518), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n535), .A2(new_n537), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n367), .ZN(new_n578));
  INV_X1    g377(.A(new_n574), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT81), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n540), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT35), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n538), .A2(new_n478), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n572), .B(new_n567), .C1(new_n514), .C2(new_n517), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR4_X1   g385(.A1(new_n478), .A2(new_n538), .A3(new_n584), .A4(KEYINPUT35), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n277), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT7), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n594));
  NOR2_X1   g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(KEYINPUT8), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n594), .B1(new_n593), .B2(new_n597), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n593), .A2(new_n597), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT97), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n600), .B1(new_n605), .B2(new_n598), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n591), .B1(new_n607), .B2(new_n265), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n259), .B2(new_n607), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n612));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G57gat), .B(G64gat), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g419(.A1(KEYINPUT93), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(G71gat), .B2(G78gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n620), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT20), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n243), .B1(new_n624), .B2(new_n623), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT96), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT94), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n630), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n623), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n603), .B2(new_n606), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n605), .A2(new_n600), .A3(new_n598), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n623), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G120gat), .B(G148gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT98), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT99), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n641), .A2(new_n654), .A3(new_n644), .ZN(new_n655));
  OAI211_X1 g454(.A(KEYINPUT10), .B(new_n640), .C1(new_n603), .C2(new_n606), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n648), .B(new_n653), .C1(new_n657), .C2(new_n647), .ZN(new_n658));
  INV_X1    g457(.A(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(new_n648), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n646), .B(KEYINPUT100), .Z(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n655), .B2(new_n656), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n639), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n589), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n367), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n231), .ZN(G1324gat));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n577), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n238), .B2(new_n669), .ZN(new_n672));
  MUX2_X1   g471(.A(new_n671), .B(new_n672), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n666), .B2(new_n574), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n568), .A2(new_n569), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(G15gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n674), .B1(new_n666), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n666), .A2(new_n576), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT101), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n638), .ZN(new_n683));
  INV_X1    g482(.A(new_n664), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n617), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n589), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n221), .A3(new_n478), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n581), .A2(new_n588), .ZN(new_n690));
  INV_X1    g489(.A(new_n617), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n541), .A2(new_n574), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n485), .B2(new_n539), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n586), .A2(new_n587), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n617), .B(KEYINPUT104), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n274), .B2(new_n275), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n252), .A2(new_n253), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n267), .A2(new_n264), .A3(new_n269), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n254), .B2(new_n262), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n206), .B1(new_n709), .B2(KEYINPUT86), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n272), .A2(new_n273), .A3(new_n207), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT102), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n685), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n703), .A2(KEYINPUT105), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n690), .B2(new_n691), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n701), .ZN(new_n721));
  INV_X1    g520(.A(new_n715), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n717), .A2(new_n724), .A3(new_n367), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n689), .B1(new_n725), .B2(new_n221), .ZN(G1328gat));
  INV_X1    g525(.A(new_n216), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n687), .A2(new_n727), .A3(new_n538), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n717), .A2(new_n724), .A3(new_n577), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n727), .ZN(G1329gat));
  NOR2_X1   g531(.A1(new_n676), .A2(G43gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n589), .A2(new_n686), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT107), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n723), .A3(new_n579), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(G43gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n703), .A2(new_n579), .A3(new_n715), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT108), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n742), .B(new_n738), .C1(new_n739), .C2(G43gat), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n737), .A2(KEYINPUT47), .B1(new_n741), .B2(new_n743), .ZN(G1330gat));
  NAND3_X1  g543(.A1(new_n703), .A2(new_n518), .A3(new_n715), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n576), .A2(G50gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n687), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(KEYINPUT48), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n716), .A2(new_n723), .A3(new_n518), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(G50gat), .B1(new_n687), .B2(new_n747), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g551(.A(new_n697), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n713), .A2(new_n639), .A3(new_n684), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n478), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n538), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n755), .B2(new_n574), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n676), .A2(G71gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g565(.A1(new_n756), .A2(new_n518), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n713), .A2(new_n638), .A3(new_n684), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n693), .B2(new_n702), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n769), .B1(new_n773), .B2(new_n367), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(KEYINPUT109), .A3(new_n478), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(G85gat), .A3(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n713), .A2(new_n638), .A3(new_n617), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n695), .B2(new_n696), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT51), .B(new_n777), .C1(new_n695), .C2(new_n696), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(KEYINPUT110), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n367), .A2(new_n684), .A3(G85gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT111), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n776), .B1(new_n785), .B2(new_n787), .ZN(G1336gat));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n538), .B(new_n770), .C1(new_n720), .C2(new_n701), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(new_n790), .B2(G92gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n577), .A2(G92gat), .A3(new_n684), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n783), .A2(new_n792), .A3(new_n784), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n783), .A2(new_n784), .A3(new_n793), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n791), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n790), .A2(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n782), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n793), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n789), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n791), .A2(new_n794), .A3(new_n796), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(KEYINPUT113), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1337gat));
  OAI21_X1  g606(.A(G99gat), .B1(new_n773), .B2(new_n574), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n676), .A2(G99gat), .A3(new_n684), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n785), .B2(new_n809), .ZN(G1338gat));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n772), .B2(new_n518), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n576), .A2(G106gat), .A3(new_n684), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT114), .Z(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n800), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  INV_X1    g615(.A(new_n813), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n785), .B2(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n815), .A2(new_n816), .B1(new_n812), .B2(new_n818), .ZN(G1339gat));
  XOR2_X1   g618(.A(new_n617), .B(KEYINPUT104), .Z(new_n820));
  INV_X1    g619(.A(new_n658), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n655), .A2(new_n656), .A3(new_n661), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT54), .B(new_n822), .C1(new_n657), .C2(new_n647), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n653), .B1(new_n662), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n705), .B2(new_n712), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n270), .A2(new_n264), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n260), .A2(new_n208), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n205), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n709), .A2(new_n207), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n664), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n820), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n829), .A2(new_n836), .A3(new_n828), .A4(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n698), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n638), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n714), .A2(new_n665), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR4_X1   g645(.A1(new_n846), .A2(new_n367), .A3(new_n538), .A4(new_n518), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n675), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n310), .A3(new_n277), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n675), .A3(new_n713), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n310), .B2(new_n850), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n675), .A3(new_n664), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n848), .A2(new_n683), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(new_n303), .ZN(G1342gat));
  NAND4_X1  g654(.A1(new_n847), .A2(new_n301), .A3(new_n675), .A4(new_n691), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n675), .A3(new_n691), .ZN(new_n857));
  AOI22_X1  g656(.A1(KEYINPUT56), .A2(new_n856), .B1(new_n857), .B2(G134gat), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n856), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(G1343gat));
  NOR3_X1   g662(.A1(new_n579), .A2(new_n367), .A3(new_n538), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n826), .A2(new_n827), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n829), .A4(new_n658), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n710), .A2(new_n869), .A3(new_n711), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n828), .B2(new_n829), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n838), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n617), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n842), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n683), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n866), .B(new_n576), .C1(new_n875), .C2(new_n844), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n846), .B2(new_n576), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n865), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n289), .B1(new_n880), .B2(new_n713), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n518), .B(new_n864), .C1(new_n843), .C2(new_n845), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n277), .A2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT58), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  INV_X1    g686(.A(new_n878), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n843), .A2(new_n845), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n518), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n276), .B(new_n864), .C1(new_n890), .C2(new_n876), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n882), .B2(new_n884), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n887), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT119), .B(new_n894), .C1(new_n891), .C2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n886), .B1(new_n896), .B2(new_n897), .ZN(G1344gat));
  AOI211_X1 g697(.A(KEYINPUT59), .B(new_n290), .C1(new_n880), .C2(new_n664), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n276), .A2(new_n639), .A3(new_n664), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n841), .A2(new_n691), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n873), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n903), .B2(new_n683), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n866), .B1(new_n904), .B2(new_n576), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n518), .B(new_n888), .C1(new_n843), .C2(new_n845), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n907), .A2(new_n664), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n900), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n664), .A2(new_n290), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n899), .A2(new_n911), .B1(new_n882), .B2(new_n912), .ZN(G1345gat));
  INV_X1    g712(.A(new_n880), .ZN(new_n914));
  OAI21_X1  g713(.A(G155gat), .B1(new_n914), .B2(new_n683), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n638), .A2(new_n279), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n882), .B2(new_n916), .ZN(G1346gat));
  NOR2_X1   g716(.A1(new_n914), .A2(new_n820), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n691), .A2(new_n287), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n918), .A2(new_n287), .B1(new_n882), .B2(new_n919), .ZN(G1347gat));
  NOR3_X1   g719(.A1(new_n577), .A2(new_n478), .A3(new_n584), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n889), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n383), .A3(new_n713), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT121), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n276), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n924), .B1(new_n383), .B2(new_n926), .ZN(G1348gat));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n664), .ZN(new_n928));
  MUX2_X1   g727(.A(new_n420), .B(G176gat), .S(new_n928), .Z(G1349gat));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n638), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(new_n409), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n377), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(G1350gat));
  AOI21_X1  g735(.A(new_n378), .B1(new_n922), .B2(new_n691), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT61), .Z(new_n938));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n378), .A3(new_n698), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n846), .A2(new_n576), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n579), .A2(new_n478), .A3(new_n577), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n713), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n942), .B(KEYINPUT122), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n905), .B2(new_n906), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(G197gat), .A3(new_n276), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n945), .A2(new_n948), .ZN(G1352gat));
  NAND2_X1  g748(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n684), .A2(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n953));
  INV_X1    g752(.A(new_n951), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n943), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n946), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n907), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(new_n684), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT124), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n958), .B2(KEYINPUT124), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n952), .B(new_n955), .C1(new_n959), .C2(new_n960), .ZN(G1353gat));
  OAI211_X1 g760(.A(KEYINPUT63), .B(G211gat), .C1(new_n957), .C2(new_n683), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n429), .B1(new_n947), .B2(new_n638), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT126), .B1(new_n964), .B2(KEYINPUT63), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n683), .B(new_n946), .C1(new_n905), .C2(new_n906), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n966), .B(new_n967), .C1(new_n968), .C2(new_n429), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n964), .A2(new_n970), .A3(KEYINPUT63), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n963), .A2(new_n965), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n944), .A2(new_n429), .A3(new_n638), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1354gat));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n617), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n698), .A2(new_n430), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n975), .A2(new_n430), .B1(new_n943), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  OAI221_X1 g778(.A(new_n979), .B1(new_n943), .B2(new_n976), .C1(new_n975), .C2(new_n430), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1355gat));
endmodule


