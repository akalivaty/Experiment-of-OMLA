

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n600, n601, n602, n603, n604, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719;

  INV_X1 U364 ( .A(n616), .ZN(n344) );
  INV_X1 U365 ( .A(n616), .ZN(n348) );
  NOR2_X1 U366 ( .A1(n715), .A2(n492), .ZN(n493) );
  XNOR2_X1 U367 ( .A(n396), .B(G469), .ZN(n502) );
  XNOR2_X1 U368 ( .A(n431), .B(n395), .ZN(n613) );
  XNOR2_X1 U369 ( .A(n416), .B(n415), .ZN(n546) );
  NOR2_X1 U370 ( .A1(G902), .A2(n607), .ZN(n416) );
  BUF_X1 U371 ( .A(G113), .Z(n352) );
  BUF_X1 U372 ( .A(G953), .Z(n342) );
  XNOR2_X1 U373 ( .A(n351), .B(n425), .ZN(n438) );
  XNOR2_X2 U374 ( .A(n525), .B(n384), .ZN(n531) );
  NOR2_X2 U375 ( .A1(n437), .A2(n436), .ZN(n518) );
  NAND2_X1 U376 ( .A1(n472), .A2(G221), .ZN(n401) );
  XNOR2_X1 U377 ( .A(n397), .B(KEYINPUT8), .ZN(n472) );
  NAND2_X1 U378 ( .A1(n546), .A2(n659), .ZN(n653) );
  XNOR2_X2 U379 ( .A(n444), .B(n389), .ZN(n431) );
  NOR2_X2 U380 ( .A1(n643), .A2(n557), .ZN(n559) );
  XNOR2_X2 U381 ( .A(n555), .B(n554), .ZN(n643) );
  NOR2_X2 U382 ( .A1(n549), .A2(n553), .ZN(n564) );
  NAND2_X2 U383 ( .A1(n564), .A2(n544), .ZN(n545) );
  INV_X1 U384 ( .A(n343), .ZN(n606) );
  NAND2_X1 U385 ( .A1(n345), .A2(n344), .ZN(n343) );
  XNOR2_X1 U386 ( .A(n604), .B(n346), .ZN(n345) );
  INV_X1 U387 ( .A(n603), .ZN(n346) );
  INV_X1 U388 ( .A(n347), .ZN(n600) );
  NAND2_X1 U389 ( .A1(n349), .A2(n348), .ZN(n347) );
  XNOR2_X1 U390 ( .A(n598), .B(n350), .ZN(n349) );
  INV_X1 U391 ( .A(n597), .ZN(n350) );
  XNOR2_X1 U392 ( .A(n424), .B(n423), .ZN(n351) );
  NOR2_X1 U393 ( .A1(n649), .A2(n510), .ZN(n367) );
  INV_X1 U394 ( .A(n571), .ZN(n657) );
  AND2_X2 U395 ( .A1(n371), .A2(n370), .ZN(n377) );
  XNOR2_X2 U396 ( .A(n448), .B(n354), .ZN(n505) );
  OR2_X2 U397 ( .A1(n595), .A2(n583), .ZN(n448) );
  XNOR2_X1 U398 ( .A(n543), .B(KEYINPUT22), .ZN(n549) );
  XNOR2_X1 U399 ( .A(G116), .B(G113), .ZN(n424) );
  NAND2_X1 U400 ( .A1(n719), .A2(n378), .ZN(n370) );
  NOR2_X1 U401 ( .A1(n379), .A2(n378), .ZN(n375) );
  XNOR2_X1 U402 ( .A(G902), .B(KEYINPUT15), .ZN(n410) );
  INV_X1 U403 ( .A(KEYINPUT71), .ZN(n362) );
  NAND2_X1 U404 ( .A1(n376), .A2(n374), .ZN(n373) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(G119), .Z(n425) );
  INV_X1 U406 ( .A(KEYINPUT3), .ZN(n423) );
  NOR2_X1 U407 ( .A1(G902), .A2(n613), .ZN(n396) );
  XNOR2_X1 U408 ( .A(n502), .B(KEYINPUT1), .ZN(n551) );
  INV_X1 U409 ( .A(n410), .ZN(n583) );
  XNOR2_X1 U410 ( .A(n438), .B(n381), .ZN(n684) );
  XNOR2_X1 U411 ( .A(KEYINPUT16), .B(G122), .ZN(n381) );
  NAND2_X1 U412 ( .A1(n357), .A2(n582), .ZN(n640) );
  XNOR2_X1 U413 ( .A(n365), .B(n413), .ZN(n414) );
  NAND2_X1 U414 ( .A1(n542), .A2(n386), .ZN(n543) );
  BUF_X1 U415 ( .A(n551), .Z(n654) );
  XOR2_X1 U416 ( .A(G104), .B(G107), .Z(n391) );
  INV_X1 U417 ( .A(KEYINPUT44), .ZN(n378) );
  NAND2_X1 U418 ( .A1(n368), .A2(n367), .ZN(n513) );
  NOR2_X1 U419 ( .A1(n513), .A2(KEYINPUT73), .ZN(n512) );
  XNOR2_X1 U420 ( .A(n411), .B(n366), .ZN(n417) );
  XNOR2_X1 U421 ( .A(n412), .B(KEYINPUT95), .ZN(n366) );
  NOR2_X1 U422 ( .A1(G237), .A2(G953), .ZN(n451) );
  NAND2_X1 U423 ( .A1(n417), .A2(G217), .ZN(n365) );
  INV_X1 U424 ( .A(G902), .ZN(n475) );
  AND2_X1 U425 ( .A1(n705), .A2(G234), .ZN(n397) );
  XNOR2_X1 U426 ( .A(G116), .B(G107), .ZN(n468) );
  XNOR2_X1 U427 ( .A(n439), .B(n403), .ZN(n462) );
  XNOR2_X1 U428 ( .A(n402), .B(KEYINPUT68), .ZN(n403) );
  INV_X1 U429 ( .A(KEYINPUT10), .ZN(n402) );
  NOR2_X1 U430 ( .A1(n647), .A2(n648), .ZN(n482) );
  BUF_X1 U431 ( .A(n538), .Z(n510) );
  NOR2_X1 U432 ( .A1(n502), .A2(n653), .ZN(n572) );
  AND2_X2 U433 ( .A1(n640), .A2(n583), .ZN(n356) );
  XNOR2_X1 U434 ( .A(n684), .B(n361), .ZN(n360) );
  XNOR2_X1 U435 ( .A(n364), .B(n444), .ZN(n363) );
  XOR2_X1 U436 ( .A(KEYINPUT89), .B(n587), .Z(n616) );
  INV_X1 U437 ( .A(n342), .ZN(n692) );
  INV_X1 U438 ( .A(KEYINPUT84), .ZN(n562) );
  INV_X1 U439 ( .A(n654), .ZN(n567) );
  AND2_X1 U440 ( .A1(n531), .A2(n387), .ZN(n353) );
  XOR2_X1 U441 ( .A(n447), .B(n446), .Z(n354) );
  AND2_X1 U442 ( .A1(n387), .A2(KEYINPUT2), .ZN(n355) );
  XNOR2_X1 U443 ( .A(n363), .B(n360), .ZN(n595) );
  NAND2_X1 U444 ( .A1(n691), .A2(n353), .ZN(n357) );
  XNOR2_X2 U445 ( .A(n580), .B(n579), .ZN(n691) );
  AND2_X4 U446 ( .A1(n641), .A2(n356), .ZN(n601) );
  XNOR2_X2 U447 ( .A(n358), .B(KEYINPUT76), .ZN(n641) );
  NAND2_X1 U448 ( .A1(n581), .A2(n691), .ZN(n358) );
  XNOR2_X2 U449 ( .A(n359), .B(G143), .ZN(n470) );
  XNOR2_X2 U450 ( .A(G128), .B(KEYINPUT81), .ZN(n359) );
  INV_X1 U451 ( .A(n443), .ZN(n361) );
  XNOR2_X1 U452 ( .A(n688), .B(n362), .ZN(n443) );
  XNOR2_X2 U453 ( .A(n701), .B(n388), .ZN(n444) );
  XNOR2_X1 U454 ( .A(n442), .B(n385), .ZN(n364) );
  XNOR2_X1 U455 ( .A(n409), .B(n408), .ZN(n607) );
  NAND2_X1 U456 ( .A1(n531), .A2(n355), .ZN(n532) );
  XNOR2_X1 U457 ( .A(n353), .B(n704), .ZN(n706) );
  XNOR2_X2 U458 ( .A(n470), .B(KEYINPUT4), .ZN(n701) );
  INV_X1 U459 ( .A(n511), .ZN(n368) );
  NOR2_X1 U460 ( .A1(n511), .A2(n510), .ZN(n369) );
  NAND2_X1 U461 ( .A1(n369), .A2(n635), .ZN(n627) );
  NAND2_X1 U462 ( .A1(n369), .A2(n633), .ZN(n632) );
  INV_X1 U463 ( .A(n626), .ZN(n379) );
  NAND2_X1 U464 ( .A1(n718), .A2(n626), .ZN(n372) );
  XNOR2_X2 U465 ( .A(n545), .B(KEYINPUT32), .ZN(n718) );
  XNOR2_X2 U466 ( .A(n380), .B(n563), .ZN(n719) );
  NAND2_X1 U467 ( .A1(n372), .A2(n378), .ZN(n371) );
  NAND2_X1 U468 ( .A1(n377), .A2(n373), .ZN(n578) );
  AND2_X1 U469 ( .A1(n718), .A2(n375), .ZN(n374) );
  INV_X1 U470 ( .A(n719), .ZN(n376) );
  NOR2_X2 U471 ( .A1(n561), .A2(n560), .ZN(n380) );
  NAND2_X1 U472 ( .A1(n518), .A2(n644), .ZN(n450) );
  NOR2_X1 U473 ( .A1(n486), .A2(n571), .ZN(n487) );
  XNOR2_X1 U474 ( .A(n400), .B(KEYINPUT78), .ZN(n383) );
  XNOR2_X1 U475 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n384) );
  AND2_X1 U476 ( .A1(G224), .A2(n705), .ZN(n385) );
  NOR2_X1 U477 ( .A1(n647), .A2(n541), .ZN(n386) );
  AND2_X1 U478 ( .A1(n639), .A2(n530), .ZN(n387) );
  BUF_X1 U479 ( .A(n643), .Z(n676) );
  XNOR2_X1 U480 ( .A(n401), .B(n383), .ZN(n409) );
  XNOR2_X1 U481 ( .A(n562), .B(KEYINPUT35), .ZN(n563) );
  XNOR2_X1 U482 ( .A(KEYINPUT67), .B(G101), .ZN(n388) );
  XNOR2_X1 U483 ( .A(G134), .B(G131), .ZN(n700) );
  XNOR2_X1 U484 ( .A(n700), .B(G146), .ZN(n389) );
  XNOR2_X1 U485 ( .A(KEYINPUT75), .B(G110), .ZN(n390) );
  XNOR2_X1 U486 ( .A(n391), .B(n390), .ZN(n688) );
  XOR2_X1 U487 ( .A(G137), .B(G140), .Z(n404) );
  XOR2_X1 U488 ( .A(n404), .B(KEYINPUT79), .Z(n393) );
  XOR2_X2 U489 ( .A(KEYINPUT64), .B(G953), .Z(n705) );
  NAND2_X1 U490 ( .A1(G227), .A2(n705), .ZN(n392) );
  XNOR2_X1 U491 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U492 ( .A(n443), .B(n394), .ZN(n395) );
  XOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n399) );
  XNOR2_X1 U494 ( .A(G128), .B(G110), .ZN(n398) );
  XNOR2_X1 U495 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X2 U496 ( .A(G146), .B(G125), .Z(n439) );
  XNOR2_X1 U497 ( .A(n462), .B(n404), .ZN(n703) );
  XOR2_X1 U498 ( .A(KEYINPUT93), .B(KEYINPUT82), .Z(n406) );
  XNOR2_X1 U499 ( .A(G119), .B(KEYINPUT92), .ZN(n405) );
  XNOR2_X1 U500 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n703), .B(n407), .ZN(n408) );
  XOR2_X1 U502 ( .A(KEYINPUT94), .B(KEYINPUT97), .Z(n413) );
  XOR2_X1 U503 ( .A(KEYINPUT96), .B(KEYINPUT20), .Z(n412) );
  NAND2_X1 U504 ( .A1(G234), .A2(n410), .ZN(n411) );
  XNOR2_X1 U505 ( .A(KEYINPUT25), .B(n414), .ZN(n415) );
  NAND2_X1 U506 ( .A1(n417), .A2(G221), .ZN(n418) );
  XOR2_X1 U507 ( .A(KEYINPUT21), .B(n418), .Z(n659) );
  NOR2_X1 U508 ( .A1(n705), .A2(G900), .ZN(n419) );
  NAND2_X1 U509 ( .A1(G902), .A2(n419), .ZN(n420) );
  NAND2_X1 U510 ( .A1(G952), .A2(n692), .ZN(n534) );
  NAND2_X1 U511 ( .A1(n420), .A2(n534), .ZN(n495) );
  NAND2_X1 U512 ( .A1(G237), .A2(G234), .ZN(n421) );
  XNOR2_X1 U513 ( .A(n421), .B(KEYINPUT14), .ZN(n642) );
  AND2_X1 U514 ( .A1(n495), .A2(n642), .ZN(n422) );
  NAND2_X1 U515 ( .A1(n572), .A2(n422), .ZN(n437) );
  NAND2_X1 U516 ( .A1(n451), .A2(G210), .ZN(n426) );
  XNOR2_X1 U517 ( .A(n426), .B(G137), .ZN(n428) );
  XNOR2_X1 U518 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n427) );
  XNOR2_X1 U519 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U520 ( .A(n438), .B(n429), .ZN(n430) );
  XNOR2_X1 U521 ( .A(n431), .B(n430), .ZN(n589) );
  OR2_X1 U522 ( .A1(n589), .A2(G902), .ZN(n433) );
  INV_X1 U523 ( .A(G472), .ZN(n432) );
  XNOR2_X2 U524 ( .A(n433), .B(n432), .ZN(n571) );
  INV_X1 U525 ( .A(G237), .ZN(n434) );
  NAND2_X1 U526 ( .A1(n475), .A2(n434), .ZN(n445) );
  NAND2_X1 U527 ( .A1(n445), .A2(G214), .ZN(n645) );
  NAND2_X1 U528 ( .A1(n657), .A2(n645), .ZN(n435) );
  XNOR2_X1 U529 ( .A(n435), .B(KEYINPUT30), .ZN(n436) );
  XOR2_X1 U530 ( .A(KEYINPUT18), .B(KEYINPUT80), .Z(n441) );
  XNOR2_X1 U531 ( .A(KEYINPUT17), .B(n439), .ZN(n440) );
  XNOR2_X1 U532 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U533 ( .A1(G210), .A2(n445), .ZN(n447) );
  INV_X1 U534 ( .A(KEYINPUT90), .ZN(n446) );
  XNOR2_X1 U535 ( .A(n505), .B(KEYINPUT38), .ZN(n644) );
  XOR2_X1 U536 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n449) );
  XNOR2_X2 U537 ( .A(n450), .B(n449), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n453) );
  NAND2_X1 U539 ( .A1(G214), .A2(n451), .ZN(n452) );
  XNOR2_X1 U540 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U541 ( .A(n454), .B(KEYINPUT12), .Z(n460) );
  XOR2_X1 U542 ( .A(G122), .B(G140), .Z(n456) );
  XNOR2_X1 U543 ( .A(n352), .B(G104), .ZN(n455) );
  XNOR2_X1 U544 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U545 ( .A(G143), .B(G131), .ZN(n457) );
  XNOR2_X1 U546 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U548 ( .A(n462), .B(n461), .ZN(n602) );
  NAND2_X1 U549 ( .A1(n602), .A2(n475), .ZN(n464) );
  XNOR2_X1 U550 ( .A(KEYINPUT13), .B(G475), .ZN(n463) );
  XNOR2_X1 U551 ( .A(n464), .B(n463), .ZN(n481) );
  INV_X1 U552 ( .A(n481), .ZN(n515) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n466) );
  XNOR2_X1 U554 ( .A(G134), .B(G122), .ZN(n465) );
  XNOR2_X1 U555 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U556 ( .A(n467), .B(KEYINPUT7), .Z(n469) );
  XNOR2_X1 U557 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U558 ( .A(n470), .B(n471), .ZN(n474) );
  NAND2_X1 U559 ( .A1(n472), .A2(G217), .ZN(n473) );
  XNOR2_X1 U560 ( .A(n474), .B(n473), .ZN(n584) );
  NAND2_X1 U561 ( .A1(n584), .A2(n475), .ZN(n477) );
  INV_X1 U562 ( .A(G478), .ZN(n476) );
  XNOR2_X1 U563 ( .A(n477), .B(n476), .ZN(n514) );
  NOR2_X1 U564 ( .A1(n515), .A2(n514), .ZN(n635) );
  NAND2_X1 U565 ( .A1(n478), .A2(n635), .ZN(n530) );
  XNOR2_X1 U566 ( .A(n530), .B(G134), .ZN(G36) );
  AND2_X1 U567 ( .A1(n515), .A2(n514), .ZN(n633) );
  NAND2_X1 U568 ( .A1(n478), .A2(n633), .ZN(n480) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U570 ( .A(n480), .B(n479), .ZN(n492) );
  XOR2_X1 U571 ( .A(G131), .B(n492), .Z(G33) );
  NAND2_X1 U572 ( .A1(n514), .A2(n481), .ZN(n647) );
  NAND2_X1 U573 ( .A1(n645), .A2(n644), .ZN(n648) );
  XNOR2_X1 U574 ( .A(KEYINPUT41), .B(n482), .ZN(n675) );
  INV_X1 U575 ( .A(n642), .ZN(n483) );
  NOR2_X1 U576 ( .A1(n546), .A2(n483), .ZN(n484) );
  NAND2_X1 U577 ( .A1(n484), .A2(n659), .ZN(n497) );
  INV_X1 U578 ( .A(n497), .ZN(n485) );
  NAND2_X1 U579 ( .A1(n485), .A2(n495), .ZN(n486) );
  XNOR2_X1 U580 ( .A(n487), .B(KEYINPUT28), .ZN(n489) );
  INV_X1 U581 ( .A(n502), .ZN(n488) );
  NAND2_X1 U582 ( .A1(n489), .A2(n488), .ZN(n511) );
  NOR2_X1 U583 ( .A1(n675), .A2(n511), .ZN(n491) );
  XNOR2_X1 U584 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n490) );
  XNOR2_X1 U585 ( .A(n491), .B(n490), .ZN(n715) );
  XNOR2_X1 U586 ( .A(n493), .B(KEYINPUT46), .ZN(n524) );
  BUF_X1 U587 ( .A(n505), .Z(n494) );
  NAND2_X1 U588 ( .A1(n495), .A2(n645), .ZN(n496) );
  NOR2_X1 U589 ( .A1(n497), .A2(n496), .ZN(n499) );
  XNOR2_X1 U590 ( .A(n571), .B(KEYINPUT6), .ZN(n553) );
  AND2_X1 U591 ( .A1(n553), .A2(n633), .ZN(n498) );
  NAND2_X1 U592 ( .A1(n499), .A2(n498), .ZN(n526) );
  NOR2_X1 U593 ( .A1(n494), .A2(n526), .ZN(n501) );
  XNOR2_X1 U594 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n500) );
  XNOR2_X1 U595 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U596 ( .A1(n503), .A2(n654), .ZN(n504) );
  XNOR2_X1 U597 ( .A(n504), .B(KEYINPUT107), .ZN(n717) );
  INV_X1 U598 ( .A(n505), .ZN(n506) );
  NAND2_X1 U599 ( .A1(n506), .A2(n645), .ZN(n509) );
  XNOR2_X1 U600 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n507) );
  XNOR2_X1 U601 ( .A(n507), .B(KEYINPUT77), .ZN(n508) );
  XNOR2_X1 U602 ( .A(n509), .B(n508), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n633), .A2(n635), .ZN(n649) );
  XOR2_X1 U604 ( .A(KEYINPUT47), .B(n512), .Z(n521) );
  NAND2_X1 U605 ( .A1(n513), .A2(KEYINPUT73), .ZN(n519) );
  INV_X1 U606 ( .A(n514), .ZN(n516) );
  NAND2_X1 U607 ( .A1(n516), .A2(n515), .ZN(n560) );
  NOR2_X1 U608 ( .A1(n494), .A2(n560), .ZN(n517) );
  NAND2_X1 U609 ( .A1(n518), .A2(n517), .ZN(n631) );
  NAND2_X1 U610 ( .A1(n519), .A2(n631), .ZN(n520) );
  NOR2_X1 U611 ( .A1(n521), .A2(n520), .ZN(n522) );
  AND2_X1 U612 ( .A1(n717), .A2(n522), .ZN(n523) );
  NAND2_X1 U613 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U614 ( .A(n526), .B(KEYINPUT104), .Z(n527) );
  NAND2_X1 U615 ( .A1(n527), .A2(n654), .ZN(n528) );
  XNOR2_X1 U616 ( .A(KEYINPUT43), .B(n528), .ZN(n529) );
  NAND2_X1 U617 ( .A1(n529), .A2(n494), .ZN(n639) );
  XNOR2_X1 U618 ( .A(n532), .B(KEYINPUT83), .ZN(n581) );
  NOR2_X1 U619 ( .A1(G898), .A2(n692), .ZN(n533) );
  XOR2_X1 U620 ( .A(KEYINPUT91), .B(n533), .Z(n689) );
  NAND2_X1 U621 ( .A1(n689), .A2(G902), .ZN(n535) );
  NAND2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n536), .A2(n642), .ZN(n537) );
  NOR2_X1 U624 ( .A1(n538), .A2(n537), .ZN(n540) );
  INV_X1 U625 ( .A(KEYINPUT0), .ZN(n539) );
  XNOR2_X1 U626 ( .A(n540), .B(n539), .ZN(n556) );
  INV_X1 U627 ( .A(n556), .ZN(n542) );
  INV_X1 U628 ( .A(n659), .ZN(n541) );
  XOR2_X1 U629 ( .A(n546), .B(KEYINPUT103), .Z(n660) );
  NOR2_X1 U630 ( .A1(n654), .A2(n660), .ZN(n544) );
  INV_X1 U631 ( .A(n546), .ZN(n547) );
  NAND2_X1 U632 ( .A1(n547), .A2(n571), .ZN(n548) );
  NOR2_X1 U633 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U634 ( .A1(n654), .A2(n550), .ZN(n626) );
  NOR2_X1 U635 ( .A1(n551), .A2(n653), .ZN(n552) );
  XNOR2_X1 U636 ( .A(n552), .B(KEYINPUT74), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n568), .A2(n553), .ZN(n555) );
  XOR2_X1 U638 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n554) );
  BUF_X1 U639 ( .A(n556), .Z(n557) );
  INV_X1 U640 ( .A(KEYINPUT34), .ZN(n558) );
  XNOR2_X1 U641 ( .A(n559), .B(n558), .ZN(n561) );
  XNOR2_X1 U642 ( .A(n564), .B(KEYINPUT86), .ZN(n565) );
  NAND2_X1 U643 ( .A1(n565), .A2(n660), .ZN(n566) );
  NOR2_X1 U644 ( .A1(n567), .A2(n566), .ZN(n618) );
  NAND2_X1 U645 ( .A1(n568), .A2(n657), .ZN(n665) );
  NOR2_X1 U646 ( .A1(n557), .A2(n665), .ZN(n570) );
  XOR2_X1 U647 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n569) );
  XNOR2_X1 U648 ( .A(n570), .B(n569), .ZN(n636) );
  NAND2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n573) );
  OR2_X1 U650 ( .A1(n557), .A2(n573), .ZN(n574) );
  XNOR2_X1 U651 ( .A(KEYINPUT99), .B(n574), .ZN(n623) );
  NOR2_X1 U652 ( .A1(n636), .A2(n623), .ZN(n575) );
  NOR2_X1 U653 ( .A1(n649), .A2(n575), .ZN(n576) );
  NOR2_X1 U654 ( .A1(n618), .A2(n576), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U656 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n579) );
  INV_X1 U657 ( .A(KEYINPUT2), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n601), .A2(G478), .ZN(n586) );
  XOR2_X1 U659 ( .A(KEYINPUT118), .B(n584), .Z(n585) );
  XNOR2_X1 U660 ( .A(n586), .B(n585), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n705), .A2(G952), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n588), .A2(n616), .ZN(G63) );
  NAND2_X1 U663 ( .A1(n601), .A2(G472), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n589), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n591), .B(n590), .ZN(n592) );
  NOR2_X2 U666 ( .A1(n592), .A2(n616), .ZN(n594) );
  XOR2_X1 U667 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n593) );
  XNOR2_X1 U668 ( .A(n594), .B(n593), .ZN(G57) );
  NAND2_X1 U669 ( .A1(n601), .A2(G210), .ZN(n598) );
  XOR2_X1 U670 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n596) );
  XNOR2_X1 U671 ( .A(n595), .B(n596), .ZN(n597) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U673 ( .A1(n601), .A2(G475), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT59), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U676 ( .A1(n601), .A2(G217), .ZN(n609) );
  XOR2_X1 U677 ( .A(KEYINPUT119), .B(n607), .Z(n608) );
  XNOR2_X1 U678 ( .A(n609), .B(n608), .ZN(n610) );
  NOR2_X1 U679 ( .A1(n610), .A2(n616), .ZN(G66) );
  NAND2_X1 U680 ( .A1(n601), .A2(G469), .ZN(n615) );
  XNOR2_X1 U681 ( .A(KEYINPUT117), .B(KEYINPUT57), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT58), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(n617) );
  NOR2_X1 U685 ( .A1(n617), .A2(n616), .ZN(G54) );
  XOR2_X1 U686 ( .A(G101), .B(n618), .Z(G3) );
  NAND2_X1 U687 ( .A1(n623), .A2(n633), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n619), .B(G104), .ZN(G6) );
  XOR2_X1 U689 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n621) );
  XNOR2_X1 U690 ( .A(G107), .B(KEYINPUT26), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(n622) );
  XOR2_X1 U692 ( .A(KEYINPUT108), .B(n622), .Z(n625) );
  NAND2_X1 U693 ( .A1(n623), .A2(n635), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(G9) );
  XNOR2_X1 U695 ( .A(G110), .B(n626), .ZN(G12) );
  XOR2_X1 U696 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n628) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(n630) );
  XOR2_X1 U698 ( .A(G128), .B(KEYINPUT110), .Z(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G30) );
  XNOR2_X1 U700 ( .A(G143), .B(n631), .ZN(G45) );
  XNOR2_X1 U701 ( .A(n632), .B(G146), .ZN(G48) );
  NAND2_X1 U702 ( .A1(n636), .A2(n633), .ZN(n634) );
  XNOR2_X1 U703 ( .A(n634), .B(n352), .ZN(G15) );
  NAND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n637), .B(KEYINPUT112), .ZN(n638) );
  XNOR2_X1 U706 ( .A(G116), .B(n638), .ZN(G18) );
  XNOR2_X1 U707 ( .A(G140), .B(n639), .ZN(G42) );
  AND2_X1 U708 ( .A1(n641), .A2(n640), .ZN(n681) );
  NAND2_X1 U709 ( .A1(G952), .A2(n642), .ZN(n674) );
  NOR2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U711 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U712 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U713 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U714 ( .A1(n676), .A2(n652), .ZN(n670) );
  XOR2_X1 U715 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n656) );
  NAND2_X1 U716 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U717 ( .A(n656), .B(n655), .ZN(n658) );
  NOR2_X1 U718 ( .A1(n658), .A2(n657), .ZN(n664) );
  NOR2_X1 U719 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U720 ( .A(KEYINPUT113), .B(n661), .Z(n662) );
  XNOR2_X1 U721 ( .A(KEYINPUT49), .B(n662), .ZN(n663) );
  NAND2_X1 U722 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U723 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U724 ( .A(KEYINPUT51), .B(n667), .ZN(n668) );
  NOR2_X1 U725 ( .A1(n668), .A2(n675), .ZN(n669) );
  NOR2_X1 U726 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U727 ( .A(KEYINPUT115), .B(n671), .Z(n672) );
  XNOR2_X1 U728 ( .A(KEYINPUT52), .B(n672), .ZN(n673) );
  NOR2_X1 U729 ( .A1(n674), .A2(n673), .ZN(n678) );
  NOR2_X1 U730 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U731 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U732 ( .A1(n679), .A2(n692), .ZN(n680) );
  NOR2_X1 U733 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U734 ( .A(KEYINPUT53), .B(KEYINPUT116), .ZN(n682) );
  XNOR2_X1 U735 ( .A(n683), .B(n682), .ZN(G75) );
  XOR2_X1 U736 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n686) );
  XNOR2_X1 U737 ( .A(G101), .B(n684), .ZN(n685) );
  XNOR2_X1 U738 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U739 ( .A(n688), .B(n687), .ZN(n690) );
  NOR2_X1 U740 ( .A1(n690), .A2(n689), .ZN(n699) );
  NAND2_X1 U741 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U742 ( .A1(n342), .A2(G224), .ZN(n693) );
  XNOR2_X1 U743 ( .A(KEYINPUT61), .B(n693), .ZN(n694) );
  NAND2_X1 U744 ( .A1(n694), .A2(G898), .ZN(n695) );
  NAND2_X1 U745 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U746 ( .A(n697), .B(KEYINPUT120), .ZN(n698) );
  XNOR2_X1 U747 ( .A(n699), .B(n698), .ZN(G69) );
  XOR2_X1 U748 ( .A(n701), .B(n700), .Z(n702) );
  XNOR2_X1 U749 ( .A(n703), .B(n702), .ZN(n708) );
  XNOR2_X1 U750 ( .A(n708), .B(KEYINPUT123), .ZN(n704) );
  NAND2_X1 U751 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U752 ( .A(n707), .B(KEYINPUT124), .ZN(n713) );
  XNOR2_X1 U753 ( .A(G227), .B(n708), .ZN(n709) );
  NAND2_X1 U754 ( .A1(n709), .A2(G900), .ZN(n710) );
  NAND2_X1 U755 ( .A1(n342), .A2(n710), .ZN(n711) );
  XOR2_X1 U756 ( .A(KEYINPUT125), .B(n711), .Z(n712) );
  NAND2_X1 U757 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U758 ( .A(n714), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U759 ( .A(G137), .B(n715), .Z(G39) );
  XOR2_X1 U760 ( .A(G125), .B(KEYINPUT37), .Z(n716) );
  XNOR2_X1 U761 ( .A(n717), .B(n716), .ZN(G27) );
  XNOR2_X1 U762 ( .A(n718), .B(G119), .ZN(G21) );
  XOR2_X1 U763 ( .A(n719), .B(G122), .Z(G24) );
endmodule

