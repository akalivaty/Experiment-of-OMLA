//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178, new_n1179,
    new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI21_X1  g032(.A(KEYINPUT68), .B1(new_n453), .B2(G2106), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(G567), .B2(new_n455), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n453), .A2(KEYINPUT68), .A3(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n463), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT71), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT69), .Z(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n464), .A2(new_n479), .A3(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n472), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND3_X1  g058(.A1(new_n467), .A2(G2105), .A3(new_n469), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n471), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n467), .A2(G138), .A3(new_n468), .A4(new_n469), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n464), .A2(new_n479), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n468), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n484), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n497), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .A3(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n508), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(G543), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n508), .A2(KEYINPUT72), .A3(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT72), .B1(new_n508), .B2(G651), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n516), .B(new_n512), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n506), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n515), .A2(new_n521), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n520), .B2(G89), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n511), .B1(new_n507), .B2(new_n509), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT73), .B(G51), .Z(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(G543), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n528), .B1(new_n534), .B2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(new_n514), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n506), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT5), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n514), .A2(G43), .B1(G651), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n563));
  AND4_X1   g138(.A1(new_n563), .A2(new_n510), .A3(new_n512), .A4(new_n516), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n563), .B1(new_n529), .B2(new_n516), .ZN(new_n565));
  OAI21_X1  g140(.A(G91), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n510), .A2(G53), .A3(G543), .A4(new_n512), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n529), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n516), .A2(G65), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n506), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n566), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n529), .A2(new_n563), .A3(new_n516), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n574), .B1(new_n581), .B2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n582), .A2(KEYINPUT76), .A3(new_n571), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(G299));
  AND2_X1   g159(.A1(new_n581), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n513), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n585), .A2(new_n588), .ZN(G288));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n579), .B2(new_n580), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n550), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n513), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n506), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT77), .Z(new_n602));
  AOI22_X1  g177(.A1(G47), .A2(new_n514), .B1(new_n520), .B2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n513), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n529), .A2(KEYINPUT78), .A3(G543), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n607), .A2(G54), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n550), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(G92), .B1(new_n564), .B2(new_n565), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n581), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n605), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n605), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT76), .B1(new_n582), .B2(new_n571), .ZN(new_n623));
  AND4_X1   g198(.A1(KEYINPUT76), .A2(new_n566), .A3(new_n571), .A4(new_n575), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n622), .B1(new_n625), .B2(G868), .ZN(G297));
  XNOR2_X1  g201(.A(G297), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n619), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n619), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n485), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n471), .A2(G135), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n636), .A2(new_n468), .A3(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n468), .B2(G111), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n634), .B(new_n635), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n474), .A2(new_n494), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT80), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2443), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT83), .ZN(new_n662));
  INV_X1    g237(.A(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(new_n660), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n673), .A2(KEYINPUT17), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n670), .B1(new_n673), .B2(KEYINPUT17), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n674), .A2(new_n675), .A3(new_n669), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  INV_X1    g267(.A(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n697));
  INV_X1    g272(.A(new_n686), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  INV_X1    g274(.A(new_n692), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(KEYINPUT86), .A3(new_n686), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n701), .A3(new_n688), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n691), .A2(new_n696), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT21), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT87), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(KEYINPUT22), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n709), .B1(new_n706), .B2(new_n710), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n681), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n715), .A2(new_n711), .A3(new_n680), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G23), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n585), .A2(new_n588), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n719), .A2(G6), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n598), .B2(new_n719), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT32), .B(G1981), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n723), .A2(new_n725), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G22), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G166), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT91), .B(G1971), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n728), .A2(new_n730), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n726), .A2(new_n731), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT34), .Z(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  INV_X1    g315(.A(G131), .ZN(new_n741));
  OR3_X1    g316(.A1(new_n470), .A2(KEYINPUT88), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n485), .A2(G119), .ZN(new_n743));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n470), .B2(new_n741), .ZN(new_n744));
  OR2_X1    g319(.A1(G95), .A2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n740), .B1(new_n748), .B2(new_n739), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT35), .B(G1991), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G24), .B(G290), .S(G16), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT89), .B(G1986), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n749), .A2(new_n750), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n738), .A2(new_n751), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT36), .Z(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT24), .B(G34), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(new_n739), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT95), .Z(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n482), .B2(new_n739), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT96), .Z(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n739), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n739), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT29), .B(G2090), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G27), .A2(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G164), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT101), .B(G2078), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n764), .B(new_n772), .C1(new_n770), .C2(new_n771), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n739), .A2(G26), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n485), .A2(G128), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n471), .A2(G140), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n468), .A2(G116), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(G29), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n774), .B(new_n780), .S(KEYINPUT28), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT93), .B(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n719), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n619), .B2(new_n719), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n773), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n719), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n556), .B2(new_n719), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT92), .Z(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G1341), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n471), .A2(G141), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n485), .A2(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT26), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n474), .A2(G105), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G32), .B(new_n802), .S(G29), .Z(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n792), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT31), .B(G11), .Z(new_n808));
  NOR2_X1   g383(.A1(new_n640), .A2(new_n739), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT30), .B(G28), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n808), .B(new_n809), .C1(new_n739), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G33), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT94), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n471), .A2(G139), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n473), .A2(G103), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT25), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n816), .C1(new_n468), .C2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(new_n739), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2072), .ZN(new_n820));
  INV_X1    g395(.A(G1961), .ZN(new_n821));
  NAND2_X1  g396(.A1(G171), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G5), .B2(G16), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n811), .B(new_n820), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G1341), .B2(new_n791), .ZN(new_n825));
  INV_X1    g400(.A(G1966), .ZN(new_n826));
  NAND2_X1  g401(.A1(G168), .A2(G16), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(G16), .B2(G21), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n807), .B(new_n825), .C1(new_n826), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n826), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT99), .Z(new_n833));
  NOR3_X1   g408(.A1(new_n788), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT23), .ZN(new_n835));
  INV_X1    g410(.A(G20), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(G16), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n835), .B(new_n837), .C1(G299), .C2(G16), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT102), .B(G1956), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n762), .A2(new_n763), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n823), .A2(new_n821), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(new_n804), .C2(new_n806), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n839), .A2(new_n840), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n834), .A2(new_n841), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n757), .A2(new_n847), .ZN(G311));
  INV_X1    g423(.A(G311), .ZN(G150));
  NAND2_X1  g424(.A1(new_n514), .A2(G55), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n520), .A2(G93), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n506), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n556), .A2(KEYINPUT103), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n851), .A2(new_n850), .A3(new_n853), .A4(KEYINPUT103), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n555), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G54), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n513), .B2(new_n606), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n863), .A2(new_n608), .B1(G651), .B2(new_n612), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n581), .B2(G92), .ZN(new_n865));
  INV_X1    g440(.A(G92), .ZN(new_n866));
  AOI211_X1 g441(.A(new_n616), .B(new_n866), .C1(new_n579), .C2(new_n580), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n628), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n861), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n871));
  AOI21_X1  g446(.A(G860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n854), .A2(G860), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT37), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(G145));
  NOR2_X1   g451(.A1(new_n818), .A2(KEYINPUT105), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n643), .Z(new_n878));
  INV_X1    g453(.A(new_n503), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n494), .A2(new_n496), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n879), .B(KEYINPUT104), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n497), .B2(new_n503), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n747), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n640), .B(new_n482), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n471), .A2(G142), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n468), .A2(G118), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(G130), .B2(new_n485), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n802), .B(new_n898), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n779), .B(new_n490), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n891), .A2(new_n904), .A3(new_n892), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT106), .B1(new_n625), .B2(new_n868), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n868), .A2(new_n578), .A3(new_n583), .A4(KEYINPUT106), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n908), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(G299), .B2(new_n619), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n911), .A4(new_n910), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n861), .B(new_n630), .Z(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n911), .A3(new_n910), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(KEYINPUT107), .A3(new_n908), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n919), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(new_n721), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n598), .B(G303), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n925), .A2(new_n926), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G868), .B2(new_n855), .ZN(G295));
  OAI21_X1  g510(.A(new_n934), .B1(G868), .B2(new_n855), .ZN(G331));
  XNOR2_X1  g511(.A(new_n533), .B(KEYINPUT74), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(G171), .A3(KEYINPUT108), .A4(new_n528), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g514(.A1(G301), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n540), .A2(new_n539), .A3(new_n542), .A4(KEYINPUT108), .ZN(new_n941));
  NAND3_X1  g516(.A1(G286), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n861), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n938), .A2(new_n942), .A3(new_n856), .A4(new_n860), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n918), .A2(new_n921), .A3(new_n946), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n943), .A2(new_n861), .A3(KEYINPUT109), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(KEYINPUT109), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n920), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n947), .A2(new_n930), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n948), .A2(new_n949), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT111), .B(new_n908), .C1(new_n909), .C2(new_n912), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n917), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT111), .B1(new_n920), .B2(new_n908), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n923), .A2(new_n946), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n930), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT112), .B1(new_n952), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n913), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n917), .A3(new_n954), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n958), .B1(new_n966), .B2(new_n953), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n967), .B2(new_n930), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n961), .A2(new_n962), .A3(new_n903), .A4(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n947), .A2(new_n930), .A3(new_n951), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n903), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n930), .B1(new_n947), .B2(new_n951), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n947), .A2(new_n951), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n932), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n903), .A3(new_n970), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n969), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND4_X1   g557(.A1(KEYINPUT43), .A2(new_n961), .A3(new_n903), .A4(new_n968), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n978), .A2(new_n962), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(G397));
  XOR2_X1   g561(.A(KEYINPUT113), .B(G1384), .Z(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n882), .B2(new_n884), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n472), .A2(G40), .A3(new_n475), .A4(new_n481), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n747), .A2(new_n750), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n802), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G2067), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n779), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(new_n992), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n779), .A2(G2067), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n993), .B1(new_n1003), .B2(KEYINPUT125), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(KEYINPUT125), .B2(new_n1003), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n993), .B2(G1996), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n992), .A2(KEYINPUT46), .A3(new_n995), .ZN(new_n1008));
  INV_X1    g583(.A(new_n998), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n992), .B1(new_n802), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1012));
  XNOR2_X1  g587(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n747), .A2(new_n750), .ZN(new_n1014));
  AND4_X1   g589(.A1(new_n998), .A2(new_n996), .A3(new_n1014), .A4(new_n994), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n993), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT48), .ZN(new_n1017));
  OR3_X1    g592(.A1(new_n993), .A2(G1986), .A3(G290), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1005), .A2(new_n1013), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1384), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n497), .B2(new_n503), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n991), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT117), .B(G8), .Z(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT118), .Z(new_n1028));
  INV_X1    g603(.A(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n598), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n519), .A2(new_n590), .ZN(new_n1031));
  OAI21_X1  g606(.A(G1981), .B1(new_n597), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1030), .A2(KEYINPUT49), .A3(new_n1032), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1027), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n721), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1030), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1028), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1027), .C1(new_n1038), .C2(G288), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1027), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G288), .A2(new_n1038), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1043), .A2(new_n1046), .A3(new_n1037), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  AOI22_X1  g624(.A1(G303), .A2(G8), .B1(new_n1049), .B2(KEYINPUT55), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(KEYINPUT55), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n991), .B1(new_n988), .B2(KEYINPUT45), .ZN(new_n1053));
  INV_X1    g628(.A(new_n989), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1023), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1971), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n1022), .C1(new_n497), .C2(new_n503), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n991), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G2090), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1052), .C1(new_n1056), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1041), .B1(new_n1048), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1058), .B1(new_n1061), .B2(new_n1070), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1053), .A2(new_n1055), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n576), .B(KEYINPUT57), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1068), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1077), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1079), .A3(KEYINPUT61), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1064), .A2(new_n786), .B1(new_n997), .B2(new_n1024), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1088), .A2(new_n1089), .B1(KEYINPUT60), .B2(new_n619), .ZN(new_n1090));
  INV_X1    g665(.A(new_n987), .ZN(new_n1091));
  INV_X1    g666(.A(new_n884), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n497), .A2(new_n503), .A3(new_n883), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT45), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n991), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(new_n995), .A3(new_n1095), .A4(new_n1055), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT58), .B(G1341), .Z(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1023), .B2(new_n991), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n555), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1082), .A2(new_n1085), .A3(new_n1090), .A4(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1086), .A2(new_n868), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1081), .B1(new_n1079), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT45), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n991), .B1(new_n1023), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1054), .B2(new_n1023), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n826), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1060), .A2(new_n763), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1025), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G168), .A2(new_n1026), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT51), .B1(new_n1117), .B2(new_n1113), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1115), .A2(new_n1118), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1023), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1095), .B1(new_n1120), .B2(new_n1057), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1059), .B1(new_n1121), .B2(KEYINPUT119), .ZN(new_n1122));
  INV_X1    g697(.A(G2090), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1071), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1094), .A2(new_n1095), .A3(new_n1055), .ZN(new_n1125));
  INV_X1    g700(.A(G1971), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1026), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1066), .B(new_n1047), .C1(new_n1128), .C2(new_n1052), .ZN(new_n1129));
  INV_X1    g704(.A(G2078), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n990), .A2(new_n1053), .A3(KEYINPUT53), .A4(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(G301), .B(KEYINPUT54), .Z(new_n1132));
  NAND4_X1  g707(.A1(new_n1094), .A2(new_n1130), .A3(new_n1095), .A4(new_n1055), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT122), .B(G1961), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1064), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1131), .A2(new_n1132), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1130), .A2(KEYINPUT53), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1108), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1135), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n1141), .B2(new_n1132), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1119), .A2(new_n1129), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1067), .B1(new_n1105), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1111), .A2(G168), .A3(new_n1025), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1129), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT121), .B(new_n1145), .C1(new_n1129), .C2(new_n1146), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1066), .A2(new_n1047), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n1116), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1151), .B(new_n1153), .C1(new_n1052), .C2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1149), .A2(new_n1150), .A3(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1144), .A2(KEYINPUT123), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT123), .B1(new_n1144), .B2(new_n1157), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1119), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1129), .A2(G301), .A3(new_n1141), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1119), .A2(new_n1161), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1119), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1158), .A2(new_n1159), .A3(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(G290), .B(G1986), .Z(new_n1169));
  AOI21_X1  g744(.A(new_n993), .B1(new_n1015), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1021), .B1(new_n1168), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g746(.A(new_n461), .B(G227), .C1(new_n662), .C2(new_n664), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n717), .A2(new_n906), .A3(new_n1173), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n980), .A2(KEYINPUT127), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g749(.A(KEYINPUT127), .B1(new_n980), .B2(new_n1174), .ZN(new_n1176));
  NOR2_X1   g750(.A1(new_n1175), .A2(new_n1176), .ZN(G308));
  NAND2_X1  g751(.A1(new_n980), .A2(new_n1174), .ZN(new_n1178));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n980), .A2(new_n1174), .A3(KEYINPUT127), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1181), .ZN(G225));
endmodule


