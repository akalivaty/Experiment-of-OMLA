

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U320 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n465) );
  XOR2_X1 U321 ( .A(KEYINPUT38), .B(n447), .Z(n494) );
  XOR2_X1 U322 ( .A(n413), .B(n412), .Z(n511) );
  NOR2_X1 U323 ( .A1(n532), .A2(n417), .ZN(n418) );
  XNOR2_X1 U324 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U325 ( .A(n337), .B(n336), .ZN(n340) );
  XNOR2_X1 U326 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U327 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U328 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U329 ( .A(n349), .B(n394), .Z(n570) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n472) );
  INV_X1 U331 ( .A(G29GAT), .ZN(n448) );
  XNOR2_X1 U332 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U333 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(G1328GAT) );
  XOR2_X1 U336 ( .A(G127GAT), .B(KEYINPUT0), .Z(n289) );
  XNOR2_X1 U337 ( .A(G113GAT), .B(KEYINPUT77), .ZN(n288) );
  XNOR2_X1 U338 ( .A(n289), .B(n288), .ZN(n380) );
  XOR2_X1 U339 ( .A(n380), .B(KEYINPUT90), .Z(n291) );
  NAND2_X1 U340 ( .A1(G225GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n291), .B(n290), .ZN(n310) );
  XOR2_X1 U342 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n293) );
  XNOR2_X1 U343 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U345 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n295) );
  XNOR2_X1 U346 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U348 ( .A(n297), .B(n296), .Z(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(G141GAT), .B(n300), .Z(n391) );
  XOR2_X1 U353 ( .A(G148GAT), .B(G134GAT), .Z(n302) );
  XNOR2_X1 U354 ( .A(G1GAT), .B(G120GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(G85GAT), .B(G57GAT), .Z(n331) );
  XOR2_X1 U357 ( .A(n303), .B(n331), .Z(n305) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(G162GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n391), .B(n306), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(n310), .B(n309), .Z(n533) );
  XOR2_X1 U363 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n316) );
  XOR2_X1 U364 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n312) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(KEYINPUT65), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n314) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n313), .B(KEYINPUT7), .ZN(n428) );
  XNOR2_X1 U369 ( .A(n314), .B(n428), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n322) );
  XOR2_X1 U371 ( .A(G1GAT), .B(G8GAT), .Z(n318) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G15GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n350) );
  XOR2_X1 U374 ( .A(G50GAT), .B(n350), .Z(n320) );
  NAND2_X1 U375 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U377 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U378 ( .A(G113GAT), .B(G141GAT), .Z(n324) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G197GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n325), .B(G36GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n548) );
  XOR2_X1 U383 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n329) );
  XNOR2_X1 U384 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U386 ( .A(n331), .B(n330), .Z(n337) );
  XOR2_X1 U387 ( .A(KEYINPUT33), .B(KEYINPUT68), .Z(n333) );
  XNOR2_X1 U388 ( .A(KEYINPUT32), .B(KEYINPUT69), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n335) );
  NAND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G71GAT), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n338), .B(G120GAT), .ZN(n381) );
  XNOR2_X1 U393 ( .A(G204GAT), .B(G92GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n339), .B(G64GAT), .ZN(n405) );
  XOR2_X1 U395 ( .A(n381), .B(n405), .Z(n341) );
  NAND2_X1 U396 ( .A1(n340), .A2(n341), .ZN(n345) );
  INV_X1 U397 ( .A(n340), .ZN(n343) );
  INV_X1 U398 ( .A(n341), .ZN(n342) );
  NAND2_X1 U399 ( .A1(n343), .A2(n342), .ZN(n344) );
  NAND2_X1 U400 ( .A1(n345), .A2(n344), .ZN(n349) );
  XOR2_X1 U401 ( .A(G148GAT), .B(G106GAT), .Z(n347) );
  XNOR2_X1 U402 ( .A(KEYINPUT71), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U404 ( .A(KEYINPUT70), .B(n348), .Z(n394) );
  NOR2_X1 U405 ( .A1(n548), .A2(n570), .ZN(n481) );
  XOR2_X1 U406 ( .A(n350), .B(KEYINPUT14), .Z(n352) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U409 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n354) );
  XNOR2_X1 U410 ( .A(KEYINPUT13), .B(KEYINPUT75), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U412 ( .A(n356), .B(n355), .Z(n364) );
  XOR2_X1 U413 ( .A(G78GAT), .B(G211GAT), .Z(n358) );
  XNOR2_X1 U414 ( .A(G71GAT), .B(G155GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U416 ( .A(G57GAT), .B(G64GAT), .Z(n360) );
  XNOR2_X1 U417 ( .A(G183GAT), .B(G127GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n574) );
  INV_X1 U421 ( .A(KEYINPUT99), .ZN(n419) );
  XOR2_X1 U422 ( .A(G176GAT), .B(G183GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U425 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n368) );
  XNOR2_X1 U426 ( .A(G190GAT), .B(KEYINPUT82), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U428 ( .A(n370), .B(n369), .Z(n409) );
  XOR2_X1 U429 ( .A(G43GAT), .B(G134GAT), .Z(n434) );
  XOR2_X1 U430 ( .A(KEYINPUT83), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U431 ( .A(KEYINPUT84), .B(KEYINPUT80), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(n434), .B(n373), .Z(n375) );
  NAND2_X1 U434 ( .A1(G227GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U436 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n377) );
  XNOR2_X1 U437 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U439 ( .A(n379), .B(n378), .Z(n383) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n409), .B(n384), .ZN(n520) );
  XOR2_X1 U443 ( .A(G211GAT), .B(KEYINPUT87), .Z(n386) );
  XNOR2_X1 U444 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n407) );
  XOR2_X1 U446 ( .A(KEYINPUT86), .B(n407), .Z(n388) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U449 ( .A(G218GAT), .B(n389), .ZN(n401) );
  XOR2_X1 U450 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n393) );
  XNOR2_X1 U451 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n390), .B(G162GAT), .ZN(n433) );
  XNOR2_X1 U453 ( .A(n391), .B(n433), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n396) );
  XNOR2_X1 U456 ( .A(n394), .B(G204GAT), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U458 ( .A(G22GAT), .B(n397), .Z(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n468) );
  NOR2_X1 U461 ( .A1(n520), .A2(n468), .ZN(n402) );
  XOR2_X1 U462 ( .A(KEYINPUT26), .B(n402), .Z(n563) );
  XOR2_X1 U463 ( .A(G36GAT), .B(G218GAT), .Z(n432) );
  XOR2_X1 U464 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n404) );
  XNOR2_X1 U465 ( .A(G8GAT), .B(KEYINPUT96), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U467 ( .A(n406), .B(n405), .Z(n408) );
  XOR2_X1 U468 ( .A(n432), .B(n411), .Z(n413) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n412) );
  XOR2_X1 U470 ( .A(n511), .B(KEYINPUT27), .Z(n422) );
  NOR2_X1 U471 ( .A1(n563), .A2(n422), .ZN(n532) );
  NAND2_X1 U472 ( .A1(n520), .A2(n511), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n414), .B(KEYINPUT98), .ZN(n415) );
  NAND2_X1 U474 ( .A1(n415), .A2(n468), .ZN(n416) );
  XNOR2_X1 U475 ( .A(KEYINPUT25), .B(n416), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  NOR2_X1 U477 ( .A1(n533), .A2(n420), .ZN(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT28), .B(KEYINPUT64), .Z(n421) );
  XNOR2_X1 U479 ( .A(n468), .B(n421), .ZN(n514) );
  NOR2_X1 U480 ( .A1(n514), .A2(n422), .ZN(n423) );
  NAND2_X1 U481 ( .A1(n533), .A2(n423), .ZN(n518) );
  XOR2_X1 U482 ( .A(KEYINPUT85), .B(n520), .Z(n424) );
  NOR2_X1 U483 ( .A1(n518), .A2(n424), .ZN(n425) );
  NOR2_X1 U484 ( .A1(n426), .A2(n425), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n427), .B(KEYINPUT100), .ZN(n480) );
  NOR2_X1 U486 ( .A1(n574), .A2(n480), .ZN(n445) );
  XOR2_X1 U487 ( .A(G85GAT), .B(n428), .Z(n430) );
  NAND2_X1 U488 ( .A1(G232GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n444) );
  XOR2_X1 U493 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n438) );
  XNOR2_X1 U494 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U496 ( .A(G92GAT), .B(G106GAT), .Z(n440) );
  XNOR2_X1 U497 ( .A(G190GAT), .B(G99GAT), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n476) );
  INV_X1 U501 ( .A(n476), .ZN(n546) );
  XNOR2_X1 U502 ( .A(KEYINPUT36), .B(n546), .ZN(n576) );
  NAND2_X1 U503 ( .A1(n445), .A2(n576), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n446), .B(KEYINPUT37), .ZN(n508) );
  NAND2_X1 U505 ( .A1(n481), .A2(n508), .ZN(n447) );
  NAND2_X1 U506 ( .A1(n533), .A2(n494), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n449) );
  XNOR2_X1 U508 ( .A(n570), .B(KEYINPUT41), .ZN(n553) );
  NOR2_X1 U509 ( .A1(n548), .A2(n553), .ZN(n453) );
  XNOR2_X1 U510 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n455) );
  INV_X1 U512 ( .A(n574), .ZN(n558) );
  NAND2_X1 U513 ( .A1(n558), .A2(n476), .ZN(n454) );
  OR2_X1 U514 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(KEYINPUT47), .ZN(n462) );
  NAND2_X1 U516 ( .A1(n574), .A2(n576), .ZN(n458) );
  XNOR2_X1 U517 ( .A(KEYINPUT45), .B(KEYINPUT109), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n458), .B(n457), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n459), .A2(n548), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n460), .A2(n570), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT48), .ZN(n535) );
  XOR2_X1 U523 ( .A(n511), .B(KEYINPUT116), .Z(n464) );
  NOR2_X1 U524 ( .A1(n535), .A2(n464), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n533), .A2(n467), .ZN(n562) );
  NAND2_X1 U526 ( .A1(n562), .A2(n468), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT55), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(n520), .ZN(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT118), .B(n471), .ZN(n559) );
  NOR2_X1 U530 ( .A1(n559), .A2(n476), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n574), .A2(n476), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(KEYINPUT16), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT76), .ZN(n479) );
  NOR2_X1 U535 ( .A1(n480), .A2(n479), .ZN(n496) );
  AND2_X1 U536 ( .A1(n481), .A2(n496), .ZN(n487) );
  NAND2_X1 U537 ( .A1(n533), .A2(n487), .ZN(n482) );
  XNOR2_X1 U538 ( .A(KEYINPUT34), .B(n482), .ZN(n483) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n511), .A2(n487), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U543 ( .A1(n487), .A2(n520), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n487), .A2(n514), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U547 ( .A1(n494), .A2(n511), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT102), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G36GAT), .B(n490), .ZN(G1329GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n492) );
  NAND2_X1 U551 ( .A1(n494), .A2(n520), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n494), .A2(n514), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n499) );
  INV_X1 U557 ( .A(n548), .ZN(n565) );
  NOR2_X1 U558 ( .A1(n565), .A2(n553), .ZN(n507) );
  NAND2_X1 U559 ( .A1(n496), .A2(n507), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT105), .ZN(n504) );
  NAND2_X1 U561 ( .A1(n504), .A2(n533), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U563 ( .A(G57GAT), .B(n500), .Z(G1332GAT) );
  NAND2_X1 U564 ( .A1(n511), .A2(n504), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n520), .A2(n504), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U570 ( .A1(n504), .A2(n514), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  AND2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n533), .A2(n515), .ZN(n509) );
  XOR2_X1 U574 ( .A(KEYINPUT107), .B(n509), .Z(n510) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n515), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n520), .A2(n515), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT44), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n517), .ZN(G1339GAT) );
  XOR2_X1 U583 ( .A(G113GAT), .B(KEYINPUT111), .Z(n523) );
  NOR2_X1 U584 ( .A1(n535), .A2(n518), .ZN(n519) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n521), .Z(n529) );
  NAND2_X1 U587 ( .A1(n529), .A2(n565), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n525) );
  INV_X1 U590 ( .A(n553), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n541), .A2(n529), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n526), .ZN(G1341GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n574), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(KEYINPUT50), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U598 ( .A1(n529), .A2(n546), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(n536), .Z(n545) );
  NAND2_X1 U603 ( .A1(n565), .A2(n545), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n539) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(n540), .Z(n543) );
  NAND2_X1 U609 ( .A1(n545), .A2(n541), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n574), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U615 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n548), .A2(n559), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n559), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  INV_X1 U628 ( .A(n562), .ZN(n564) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n577) );
  AND2_X1 U630 ( .A1(n577), .A2(n565), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

