//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G116), .A2(G270), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  AND3_X1   g0029(.A1(new_n218), .A2(new_n228), .A3(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n254), .B1(new_n255), .B2(new_n252), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT69), .B1(new_n269), .B2(new_n206), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n259), .B2(new_n260), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n206), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G226), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n261), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n263), .B(new_n277), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n281), .A2(G179), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n283), .A2(new_n214), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n207), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G50), .A2(G58), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n207), .B1(new_n294), .B2(new_n220), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT71), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n285), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n207), .A3(G1), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G50), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n206), .B2(G20), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n300), .A2(new_n302), .B1(new_n301), .B2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n281), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n282), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n304), .B(KEYINPUT9), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n281), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n281), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  INV_X1    g0120(.A(new_n309), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n311), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n322), .A2(new_n317), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n308), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n206), .A2(G20), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n300), .A2(G77), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT73), .B1(new_n299), .B2(new_n255), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n299), .A2(KEYINPUT73), .A3(new_n255), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n286), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(G20), .B2(G77), .ZN(new_n336));
  INV_X1    g0136(.A(new_n289), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n291), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n284), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n341), .B1(new_n203), .B2(new_n252), .C1(new_n256), .C2(new_n219), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n262), .ZN(new_n343));
  INV_X1    g0143(.A(G244), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n277), .C1(new_n344), .C2(new_n280), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT72), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(KEYINPUT72), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(KEYINPUT72), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n310), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n252), .A2(new_n253), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n278), .ZN(new_n357));
  INV_X1    g0157(.A(new_n280), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n262), .B1(G238), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n359), .A2(new_n277), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n359), .B2(new_n277), .ZN(new_n363));
  OAI21_X1  g0163(.A(G190), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(new_n277), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n360), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(KEYINPUT13), .A3(new_n277), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(G200), .A3(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n288), .B2(new_n255), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n300), .A2(G68), .A3(new_n328), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT12), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n299), .B2(new_n220), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n298), .A2(G1), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G20), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n376), .A2(KEYINPUT12), .A3(G68), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n371), .B(new_n372), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT11), .B1(new_n370), .B2(new_n285), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n364), .A2(new_n368), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n366), .A2(G169), .A3(new_n367), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n366), .A2(new_n385), .A3(G169), .A4(new_n367), .ZN(new_n386));
  OAI21_X1  g0186(.A(G179), .B1(new_n362), .B2(new_n363), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n380), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G179), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n340), .B1(new_n346), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n350), .A2(new_n305), .A3(new_n351), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n353), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  INV_X1    g0196(.A(new_n300), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n337), .A2(new_n328), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n397), .A2(new_n398), .B1(new_n376), .B2(new_n337), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n250), .A2(new_n207), .A3(new_n251), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(KEYINPUT3), .A2(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(KEYINPUT3), .A2(G33), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n406), .B2(new_n207), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G58), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n220), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n291), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n284), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT78), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n401), .A2(new_n402), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n220), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n417), .B1(new_n423), .B2(new_n414), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n419), .A2(new_n424), .A3(KEYINPUT78), .A4(new_n285), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n400), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n275), .A2(new_n270), .A3(new_n273), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n358), .A2(G232), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n432), .B1(new_n356), .B2(new_n257), .C1(new_n278), .C2(new_n256), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n262), .ZN(new_n434));
  AOI21_X1  g0234(.A(G200), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n428), .B2(new_n430), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n277), .A2(KEYINPUT79), .A3(new_n429), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G190), .B1(new_n433), .B2(new_n262), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n396), .B1(new_n427), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n434), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n305), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n437), .A2(new_n438), .A3(new_n391), .A4(new_n434), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n427), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n419), .A2(new_n424), .A3(new_n285), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n399), .B1(new_n451), .B2(new_n425), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n444), .A2(new_n445), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT18), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n435), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n440), .A2(new_n437), .A3(new_n438), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n457), .A3(KEYINPUT17), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n442), .A2(new_n448), .A3(new_n454), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n327), .A2(new_n395), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT5), .B1(new_n265), .B2(new_n267), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n206), .B(G45), .C1(new_n464), .C2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n262), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n467), .A2(G270), .B1(new_n272), .B2(new_n466), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(new_n253), .C1(new_n404), .C2(new_n405), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(KEYINPUT85), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G264), .B(G1698), .C1(new_n404), .C2(new_n405), .ZN(new_n474));
  INV_X1    g0274(.A(G303), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n252), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT86), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n261), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n479), .B(new_n476), .C1(new_n471), .C2(new_n472), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n469), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G116), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n299), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n206), .A2(G33), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n284), .A2(new_n376), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n486), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(G20), .B1(G33), .B2(G283), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n249), .A2(G97), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n494), .A2(new_n495), .B1(new_n283), .B2(new_n214), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n484), .A2(G116), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(G20), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT20), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n496), .A2(KEYINPUT20), .A3(new_n499), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n493), .B(KEYINPUT87), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT87), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n501), .A2(new_n500), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n492), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n483), .A2(G179), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n305), .B1(new_n502), .B2(new_n505), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n476), .B1(new_n471), .B2(new_n472), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n262), .B1(new_n509), .B2(KEYINPUT86), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n468), .B1(new_n510), .B2(new_n481), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT21), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n508), .B2(new_n511), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(G200), .ZN(new_n516));
  INV_X1    g0316(.A(new_n506), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(new_n310), .C2(new_n511), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OR3_X1    g0319(.A1(new_n491), .A2(KEYINPUT84), .A3(new_n333), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT84), .B1(new_n491), .B2(new_n333), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n207), .B1(new_n355), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G87), .B2(new_n204), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n286), .B2(new_n202), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n207), .B(G68), .C1(new_n404), .C2(new_n405), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(new_n285), .B1(new_n299), .B2(new_n333), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G33), .B1(new_n485), .B2(new_n487), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(G1698), .C1(new_n404), .C2(new_n405), .ZN(new_n532));
  OAI211_X1 g0332(.A(G238), .B(new_n253), .C1(new_n404), .C2(new_n405), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n262), .ZN(new_n535));
  INV_X1    g0335(.A(G250), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n268), .B2(G1), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n206), .A2(new_n271), .A3(G45), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n261), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(G179), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n534), .B2(new_n262), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n305), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n535), .A2(new_n540), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(G190), .ZN(new_n547));
  INV_X1    g0347(.A(new_n491), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G87), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n546), .A2(new_n529), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n515), .A2(new_n519), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n299), .A2(new_n203), .ZN(new_n553));
  NOR2_X1   g0353(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n555), .A2(new_n557), .B1(new_n548), .B2(G107), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n207), .B(G87), .C1(new_n404), .C2(new_n405), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT22), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT22), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n252), .A2(new_n561), .A3(new_n207), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n249), .B1(new_n497), .B2(new_n498), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n207), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n564), .A2(new_n207), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(KEYINPUT88), .A3(new_n568), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(KEYINPUT24), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT88), .B1(new_n563), .B2(new_n568), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT24), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n284), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n573), .A2(KEYINPUT89), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT89), .B1(new_n573), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n558), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n467), .A2(G264), .ZN(new_n580));
  INV_X1    g0380(.A(new_n465), .ZN(new_n581));
  XNOR2_X1  g0381(.A(KEYINPUT68), .B(G41), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n272), .C1(KEYINPUT5), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n536), .A2(new_n253), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G257), .B2(new_n253), .ZN(new_n585));
  INV_X1    g0385(.A(G294), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n585), .A2(new_n406), .B1(new_n249), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n262), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n580), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n305), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G179), .B2(new_n589), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n579), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n589), .A2(new_n310), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(G200), .B2(new_n589), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(new_n558), .C1(new_n578), .C2(new_n577), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT6), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n203), .A2(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G97), .A2(G107), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n204), .A2(new_n600), .A3(new_n602), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(G20), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n291), .A2(G77), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n203), .B1(new_n421), .B2(new_n422), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n285), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n376), .A2(G97), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n548), .B2(G97), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(new_n261), .C1(new_n463), .C2(new_n465), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n583), .ZN(new_n617));
  AND2_X1   g0417(.A1(KEYINPUT4), .A2(G244), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n253), .B(new_n618), .C1(new_n404), .C2(new_n405), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G283), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n344), .B1(new_n250), .B2(new_n251), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(KEYINPUT4), .ZN(new_n622));
  OAI21_X1  g0422(.A(G250), .B1(new_n404), .B2(new_n405), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n253), .B1(new_n623), .B2(KEYINPUT4), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n262), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n615), .B1(G200), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n626), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G190), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n617), .A2(new_n625), .A3(new_n391), .ZN(new_n630));
  AOI21_X1  g0430(.A(G169), .B1(new_n617), .B2(new_n625), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT81), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n617), .A2(new_n625), .A3(new_n391), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT81), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n612), .B2(new_n614), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n627), .A2(new_n629), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT82), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n462), .A2(new_n552), .A3(new_n598), .A4(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n388), .A2(new_n389), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n394), .B2(new_n382), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n442), .A3(new_n458), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n448), .A2(new_n454), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n320), .A2(new_n326), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n308), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n515), .ZN(new_n648));
  INV_X1    g0448(.A(new_n558), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n573), .A2(new_n576), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n573), .A2(KEYINPUT89), .A3(new_n576), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(KEYINPUT92), .A3(new_n591), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n579), .B2(new_n592), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n648), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT91), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n305), .B1(new_n535), .B2(new_n540), .ZN(new_n660));
  AOI211_X1 g0460(.A(new_n391), .B(new_n539), .C1(new_n534), .C2(new_n262), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n541), .B(KEYINPUT91), .C1(new_n305), .C2(new_n542), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n529), .B2(new_n522), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n596), .A2(new_n550), .A3(new_n636), .A4(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n632), .A2(new_n544), .A3(new_n550), .A4(new_n635), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n668), .B2(KEYINPUT26), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n545), .A2(new_n310), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n542), .A2(new_n347), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n528), .A2(new_n285), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n333), .A2(new_n299), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n549), .A3(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n662), .A2(new_n663), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n530), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n626), .A2(new_n305), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n634), .B1(new_n678), .B2(new_n633), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n615), .B1(new_n630), .B2(KEYINPUT81), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n669), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT93), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT93), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n669), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n658), .A2(new_n667), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n647), .B1(new_n461), .B2(new_n688), .ZN(G369));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n375), .A2(new_n207), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n648), .B(new_n518), .C1(new_n517), .C2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n515), .A2(new_n506), .A3(new_n696), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n690), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n654), .A2(new_n697), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n597), .A2(new_n701), .B1(new_n593), .B2(new_n697), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT92), .B1(new_n654), .B2(new_n591), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n579), .A2(new_n656), .A3(new_n592), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n697), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n515), .A2(new_n593), .A3(new_n596), .A4(new_n697), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(G399));
  NAND2_X1  g0508(.A1(new_n210), .A2(new_n582), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n216), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  OR3_X1    g0513(.A1(new_n688), .A2(KEYINPUT29), .A3(new_n696), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n552), .A2(new_n598), .A3(new_n638), .A4(new_n697), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n628), .A2(new_n661), .A3(new_n580), .A4(new_n588), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n511), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n589), .A2(new_n391), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n542), .B(KEYINPUT94), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n511), .A3(new_n626), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n717), .A2(new_n511), .A3(new_n716), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n696), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n715), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n596), .A2(new_n550), .A3(new_n636), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n648), .B2(new_n593), .ZN(new_n729));
  INV_X1    g0529(.A(new_n677), .ZN(new_n730));
  INV_X1    g0530(.A(new_n681), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT26), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n665), .C1(KEYINPUT26), .C2(new_n668), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n697), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n714), .A2(new_n727), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n713), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(new_n709), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n298), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n206), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n700), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n698), .A2(new_n699), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(G330), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n210), .A2(new_n252), .ZN(new_n747));
  INV_X1    g0547(.A(G355), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n747), .A2(new_n748), .B1(G116), .B2(new_n210), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n246), .A2(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n210), .A2(new_n406), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n268), .B2(new_n217), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n214), .B1(G20), .B2(new_n305), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n743), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT95), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(new_n310), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(new_n391), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n310), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n409), .B1(new_n768), .B2(new_n301), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n771), .A2(new_n391), .A3(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT96), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n772), .A2(KEYINPUT96), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n769), .B1(new_n777), .B2(G77), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  OR3_X1    g0582(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT32), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n766), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n783), .B(new_n784), .C1(new_n220), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n207), .B1(new_n780), .B2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n406), .B1(new_n789), .B2(G97), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n391), .A2(G200), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT98), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n771), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G87), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n763), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n790), .B1(new_n795), .B2(new_n203), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  OR3_X1    g0599(.A1(new_n779), .A2(new_n787), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n781), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G329), .ZN(new_n802));
  INV_X1    g0602(.A(new_n772), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n252), .B(new_n805), .C1(G322), .C2(new_n764), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n788), .A2(new_n586), .ZN(new_n807));
  OR2_X1    g0607(.A1(KEYINPUT33), .A2(G317), .ZN(new_n808));
  NAND2_X1  g0608(.A1(KEYINPUT33), .A2(G317), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n786), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n807), .B(new_n810), .C1(G326), .C2(new_n767), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n797), .A2(G303), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n794), .A2(G283), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n806), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n800), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n757), .ZN(new_n816));
  INV_X1    g0616(.A(new_n756), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n761), .B1(new_n815), .B2(new_n816), .C1(new_n745), .C2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n746), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  OAI21_X1  g0620(.A(new_n696), .B1(new_n339), .B2(new_n332), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n353), .A2(new_n394), .A3(new_n697), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT101), .B1(new_n688), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n515), .B1(new_n704), .B2(new_n705), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n669), .A2(new_n683), .A3(new_n686), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n686), .B1(new_n669), .B2(new_n683), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n824), .A2(new_n666), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n394), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n821), .B1(new_n348), .B2(new_n352), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n828), .A2(new_n829), .A3(new_n696), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT101), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n394), .A2(new_n696), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n829), .A2(new_n394), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n688), .B2(new_n696), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n743), .B1(new_n839), .B2(new_n727), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n727), .B2(new_n839), .ZN(new_n841));
  INV_X1    g0641(.A(new_n743), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n757), .A2(new_n754), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n255), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n252), .B1(new_n781), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n795), .A2(new_n220), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(G58), .C2(new_n789), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n301), .B2(new_n798), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT100), .Z(new_n850));
  AOI22_X1  g0650(.A1(new_n764), .A2(G143), .B1(G137), .B2(new_n767), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n851), .B1(new_n290), .B2(new_n786), .C1(new_n776), .C2(new_n782), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT34), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n252), .B1(new_n797), .B2(G107), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT99), .Z(new_n855));
  OAI22_X1  g0655(.A1(new_n776), .A2(new_n488), .B1(new_n796), .B2(new_n795), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n789), .A2(G97), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n857), .B1(new_n804), .B2(new_n781), .C1(new_n765), .C2(new_n586), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n786), .A2(new_n859), .B1(new_n768), .B2(new_n475), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n850), .A2(new_n853), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n837), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n844), .B1(new_n816), .B2(new_n862), .C1(new_n863), .C2(new_n755), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n841), .A2(new_n864), .ZN(G384));
  NAND2_X1  g0665(.A1(new_n605), .A2(new_n607), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT35), .ZN(new_n867));
  OAI211_X1 g0667(.A(G116), .B(new_n215), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OAI21_X1  g0670(.A(G77), .B1(new_n409), .B2(new_n220), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n871), .A2(new_n216), .B1(G50), .B2(new_n220), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(G1), .A3(new_n298), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT102), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n688), .A2(KEYINPUT101), .A3(new_n822), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n831), .B1(new_n827), .B2(new_n830), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n835), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n399), .B1(new_n418), .B2(new_n419), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n694), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  INV_X1    g0682(.A(new_n694), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n427), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT104), .B1(new_n452), .B2(new_n694), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n427), .A2(new_n446), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n452), .A2(new_n457), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n889), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n880), .B1(new_n453), .B2(new_n694), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI221_X4 g0693(.A(new_n879), .B1(new_n459), .B2(new_n881), .C1(new_n890), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n459), .A2(new_n881), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n389), .A2(new_n696), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n390), .A2(KEYINPUT103), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT103), .B1(new_n390), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n388), .A2(new_n382), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n901), .A2(new_n902), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n878), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n897), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT39), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n640), .A2(new_n696), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n884), .A2(new_n885), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n888), .A2(new_n889), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n890), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT105), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n459), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n459), .A2(new_n910), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT105), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n894), .B1(new_n918), .B2(new_n879), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n908), .B(new_n909), .C1(new_n919), .C2(KEYINPUT39), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n644), .A2(new_n883), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n905), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n461), .B1(new_n714), .B2(new_n735), .ZN(new_n924));
  INV_X1    g0724(.A(new_n647), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n923), .B(new_n926), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n918), .A2(new_n879), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n907), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n904), .A2(new_n726), .A3(new_n863), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT40), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n930), .B2(new_n898), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n462), .A2(new_n726), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(G330), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n927), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n206), .B2(new_n740), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n927), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n875), .B1(new_n941), .B2(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n674), .A2(new_n696), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n677), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(new_n665), .C2(new_n944), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n615), .A2(new_n696), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n636), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n681), .A2(new_n696), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n515), .A2(new_n697), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n959), .A2(KEYINPUT42), .A3(new_n598), .A4(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT42), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n952), .A2(new_n953), .B1(new_n957), .B2(new_n956), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(new_n707), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n731), .B1(new_n964), .B2(new_n593), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n697), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n949), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n968), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n969), .B2(new_n970), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n972), .A2(new_n975), .B1(new_n703), .B2(new_n964), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n969), .A2(new_n970), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n703), .A2(new_n964), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n977), .A2(new_n978), .A3(new_n971), .A4(new_n974), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n709), .B(KEYINPUT41), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n959), .A2(new_n982), .A3(new_n706), .A4(new_n707), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n706), .A2(new_n707), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT110), .B1(new_n964), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n964), .A2(new_n984), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n983), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(new_n700), .A3(new_n702), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n707), .B1(new_n702), .B2(new_n961), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n700), .A2(KEYINPUT111), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n700), .A2(KEYINPUT111), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n736), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n988), .A2(new_n991), .A3(new_n703), .A4(new_n992), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n994), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n981), .B1(new_n1003), .B2(new_n737), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n980), .B1(new_n1004), .B2(new_n742), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT112), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n980), .B(KEYINPUT112), .C1(new_n1004), .C2(new_n742), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n238), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n758), .B1(new_n210), .B2(new_n333), .C1(new_n1010), .C2(new_n751), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n743), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n406), .B1(new_n765), .B2(new_n475), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT46), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n798), .A2(new_n1015), .A3(new_n486), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(G317), .C2(new_n801), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n777), .A2(G283), .B1(new_n794), .B2(G97), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1015), .B1(new_n798), .B2(new_n488), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n768), .A2(new_n804), .B1(new_n788), .B2(new_n203), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G294), .B2(new_n785), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n788), .A2(new_n220), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G143), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n768), .B2(new_n1025), .C1(new_n782), .C2(new_n786), .ZN(new_n1026));
  INV_X1    g0826(.A(G137), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n252), .B1(new_n781), .B2(new_n1027), .C1(new_n765), .C2(new_n290), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G58), .B2(new_n797), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n301), .B2(new_n776), .C1(new_n255), .C2(new_n795), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1022), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT47), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n757), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1013), .B1(new_n1034), .B2(new_n1035), .C1(new_n948), .C2(new_n817), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1009), .A2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n1000), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n702), .A2(new_n817), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n747), .A2(new_n710), .B1(G107), .B2(new_n210), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n235), .A2(G45), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n710), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n289), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n751), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1040), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n743), .B1(new_n1048), .B2(new_n759), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n252), .B1(new_n801), .B2(G326), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n798), .A2(new_n586), .B1(new_n859), .B2(new_n788), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n764), .A2(G317), .B1(G311), .B2(new_n785), .ZN(new_n1052));
  INV_X1    g0852(.A(G322), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n768), .C1(new_n776), .C2(new_n475), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1050), .B1(new_n488), .B2(new_n795), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n789), .A2(new_n334), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n768), .B2(new_n782), .C1(new_n289), .C2(new_n786), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n803), .A2(new_n220), .B1(new_n781), .B2(new_n290), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n406), .B(new_n1063), .C1(G50), .C2(new_n764), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n797), .A2(G77), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n202), .C2(new_n795), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1059), .A2(new_n1060), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1049), .B1(new_n1067), .B2(new_n757), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1038), .A2(new_n742), .B1(new_n1039), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n739), .B1(new_n1000), .B2(new_n736), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT115), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1070), .A2(new_n1071), .B1(new_n737), .B2(new_n1038), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(G393));
  NAND2_X1  g0874(.A1(new_n994), .A2(new_n1002), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1001), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n739), .A3(new_n1003), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n994), .A2(new_n742), .A3(new_n1002), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n243), .A2(new_n751), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n758), .B1(new_n202), .B2(new_n210), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n743), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n203), .A2(new_n795), .B1(new_n798), .B2(new_n859), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n406), .B1(new_n1053), .B2(new_n781), .C1(new_n803), .C2(new_n586), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n475), .A2(new_n786), .B1(new_n488), .B2(new_n788), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n764), .A2(G311), .B1(G317), .B2(new_n767), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n764), .A2(G159), .B1(G150), .B2(new_n767), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n788), .A2(new_n255), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n252), .B1(new_n781), .B2(new_n1025), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G50), .C2(new_n785), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G68), .A2(new_n797), .B1(new_n794), .B2(G87), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n776), .C2(new_n289), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1086), .A2(new_n1088), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1082), .B1(new_n1096), .B2(new_n757), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n959), .B2(new_n817), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1079), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1078), .A2(KEYINPUT116), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT116), .B1(new_n1078), .B2(new_n1099), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(G390));
  OAI21_X1  g0903(.A(new_n908), .B1(new_n919), .B2(KEYINPUT39), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n904), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n833), .B2(new_n835), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1106), .B2(new_n909), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n690), .B1(new_n715), .B2(new_n725), .ZN(new_n1108));
  AND4_X1   g0908(.A1(KEYINPUT117), .A2(new_n1108), .A3(new_n904), .A4(new_n863), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n835), .B1(new_n734), .B2(new_n837), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n909), .B1(new_n1110), .B2(new_n904), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n929), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n904), .A3(new_n863), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1107), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n461), .A2(new_n727), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n924), .A2(new_n925), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1105), .B1(new_n727), .B2(new_n837), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1113), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1122), .A2(new_n878), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1110), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n709), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1119), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n714), .A2(new_n735), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n647), .B(new_n1127), .C1(new_n1128), .C2(new_n461), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1122), .A2(new_n1110), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1122), .A2(new_n878), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1126), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n843), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n781), .A2(new_n586), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1091), .B(new_n1136), .C1(G116), .C2(new_n764), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n203), .B2(new_n786), .C1(new_n859), .C2(new_n768), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n847), .B(new_n1138), .C1(G97), .C2(new_n777), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n252), .B1(new_n797), .B2(G87), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT120), .Z(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT118), .Z(new_n1143));
  OAI22_X1  g0943(.A1(new_n776), .A2(new_n1143), .B1(new_n1027), .B2(new_n786), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n797), .A2(G150), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT53), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n795), .A2(new_n301), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n801), .A2(G125), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n252), .B(new_n1149), .C1(new_n765), .C2(new_n845), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n768), .A2(new_n1151), .B1(new_n788), .B2(new_n782), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1139), .A2(new_n1141), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n743), .B1(new_n337), .B2(new_n1135), .C1(new_n1154), .C2(new_n816), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1104), .B2(new_n754), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1118), .B2(new_n741), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1134), .A2(new_n1159), .ZN(G378));
  OAI21_X1  g0960(.A(new_n1024), .B1(new_n768), .B2(new_n486), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n794), .A2(G58), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G107), .A2(new_n764), .B1(new_n772), .B2(new_n334), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n406), .A2(new_n582), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G283), .B2(new_n801), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1065), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1161), .B(new_n1166), .C1(G97), .C2(new_n785), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT58), .Z(new_n1168));
  OAI211_X1 g0968(.A(new_n1164), .B(new_n301), .C1(G33), .C2(G41), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n765), .A2(new_n1151), .B1(new_n803), .B2(new_n1027), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G150), .B2(new_n789), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G125), .A2(new_n767), .B1(new_n785), .B2(G132), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n798), .C2(new_n1143), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n794), .A2(G159), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n801), .C2(G124), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1168), .B(new_n1169), .C1(new_n1174), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT121), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n816), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1180), .B2(new_n1179), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n743), .C1(G50), .C2(new_n1135), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n304), .A2(new_n883), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n327), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n316), .B1(KEYINPUT76), .B2(new_n312), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n324), .B1(new_n1188), .B2(new_n313), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n326), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n307), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1186), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1185), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n327), .A2(new_n1186), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1184), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1183), .B1(new_n1199), .B2(new_n754), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n932), .A2(G330), .A3(new_n934), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n921), .B1(new_n1106), .B2(new_n899), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1198), .B1(new_n1202), .B2(new_n920), .ZN(new_n1203));
  AND4_X1   g1003(.A1(new_n920), .A2(new_n905), .A3(new_n1198), .A4(new_n922), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n923), .A2(new_n1199), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n920), .A3(new_n1198), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1201), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1200), .B1(new_n1210), .B2(new_n742), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1133), .A2(new_n1120), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n739), .B1(new_n1212), .B2(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1115), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1107), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1125), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1129), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1210), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1211), .B1(new_n1213), .B2(new_n1221), .ZN(G375));
  NOR2_X1   g1022(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1129), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(new_n1132), .A3(new_n981), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n743), .B1(G68), .B2(new_n1135), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n406), .B1(new_n781), .B2(new_n475), .C1(new_n765), .C2(new_n859), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G77), .B2(new_n794), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n202), .B2(new_n798), .C1(new_n203), .C2(new_n776), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1061), .B1(new_n768), .B2(new_n586), .C1(new_n488), .C2(new_n786), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n406), .B1(new_n764), .B2(G137), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n772), .A2(G150), .B1(G128), .B2(new_n801), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n789), .A2(G50), .B1(G132), .B2(new_n767), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1162), .B1(new_n1143), .B2(new_n786), .C1(new_n798), .C2(new_n782), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1230), .A2(new_n1231), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1227), .B1(new_n1237), .B2(new_n757), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n904), .B2(new_n755), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n741), .B(KEYINPUT122), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1239), .B1(new_n1223), .B2(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1226), .A2(new_n1241), .ZN(G381));
  OAI211_X1 g1042(.A(new_n819), .B(new_n1069), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1243));
  OR3_X1    g1043(.A1(G381), .A2(G384), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1102), .A2(new_n1009), .A3(new_n1036), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G378), .A2(new_n1244), .A3(G375), .A4(new_n1245), .ZN(G407));
  AOI21_X1  g1046(.A(new_n1158), .B1(new_n1133), .B2(new_n1126), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n695), .A2(G213), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G375), .C2(new_n1250), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1243), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1253), .A2(new_n1245), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1254), .A3(new_n1243), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1253), .A2(new_n1245), .B1(new_n1259), .B2(new_n1257), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1211), .C1(new_n1213), .C2(new_n1221), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n981), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1218), .B2(new_n1129), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1220), .B1(new_n1264), .B2(new_n1240), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1247), .B1(new_n1265), .B2(new_n1200), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1249), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n709), .B1(new_n1269), .B2(new_n1225), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1224), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1241), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G384), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G384), .B(new_n1273), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1272), .A2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1261), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1262), .A2(new_n1266), .A3(KEYINPUT123), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1248), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1249), .A2(G2897), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1276), .B(new_n1289), .C1(new_n1272), .C2(new_n1279), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G2897), .B(new_n1249), .C1(new_n1277), .C2(new_n1280), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1286), .A2(new_n1248), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1283), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1290), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(new_n1267), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1267), .A2(KEYINPUT62), .A3(new_n1281), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1296), .B1(new_n1303), .B2(new_n1305), .ZN(G405));
  AND2_X1   g1106(.A1(G375), .A2(new_n1247), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1262), .ZN(new_n1308));
  OR3_X1    g1108(.A1(new_n1307), .A2(new_n1281), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1281), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1304), .ZN(G402));
endmodule


