//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G116), .A2(G270), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OAI21_X1  g0046(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G150), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT8), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(new_n202), .B2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(KEYINPUT8), .A3(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n209), .A2(G33), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n247), .B1(new_n248), .B2(new_n250), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n217), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n261), .A3(new_n217), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n257), .A2(new_n263), .B1(new_n201), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n263), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n208), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G50), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  OAI211_X1 g0072(.A(G1), .B(G13), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n275), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n273), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G222), .ZN(new_n286));
  INV_X1    g0086(.A(G77), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(G1698), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n286), .B1(new_n287), .B2(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n280), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n270), .B1(new_n293), .B2(G169), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n270), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT72), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(G190), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n266), .A2(KEYINPUT9), .A3(new_n269), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n293), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n299), .B2(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n296), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n288), .A2(new_n312), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n310), .B1(new_n290), .B2(new_n311), .C1(new_n279), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n292), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(new_n276), .ZN(new_n317));
  INV_X1    g0117(.A(new_n278), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(G238), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n315), .B2(new_n319), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n315), .A2(new_n319), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n303), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n265), .A2(new_n221), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n221), .A2(G20), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(new_n256), .B2(new_n287), .C1(new_n250), .C2(new_n201), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n263), .A3(KEYINPUT11), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n265), .A2(new_n259), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G68), .A3(new_n268), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT11), .B1(new_n331), .B2(new_n263), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n324), .A2(new_n327), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(G169), .B1(new_n321), .B2(new_n322), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(G169), .C1(new_n321), .C2(new_n322), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n326), .A2(G179), .A3(new_n320), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n345), .B2(new_n338), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n347), .A2(new_n256), .B1(new_n209), .B2(new_n287), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT8), .B(G58), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n250), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n259), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT70), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n333), .A2(G77), .A3(new_n268), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G77), .B2(new_n264), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n285), .A2(G232), .B1(G107), .B2(new_n284), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n220), .B2(new_n290), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n273), .B1(new_n357), .B2(KEYINPUT69), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT69), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n356), .B(new_n359), .C1(new_n220), .C2(new_n290), .ZN(new_n360));
  INV_X1    g0160(.A(G244), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n276), .B1(new_n278), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT68), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n358), .A2(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n355), .B1(new_n366), .B2(new_n303), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT71), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(G190), .ZN(new_n370));
  OAI211_X1 g0170(.A(KEYINPUT71), .B(new_n355), .C1(new_n366), .C2(new_n303), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n358), .A2(new_n360), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(new_n364), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n295), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n355), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(G169), .C2(new_n366), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n309), .A2(new_n346), .A3(new_n372), .A4(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT7), .B1(new_n288), .B2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n284), .A2(new_n209), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n379), .B(G68), .C1(new_n380), .C2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(G58), .B(G68), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n259), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT76), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n385), .B1(new_n209), .B2(new_n284), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n281), .A2(new_n283), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT7), .B(new_n209), .C1(new_n283), .C2(new_n393), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT75), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(KEYINPUT74), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n281), .A2(new_n283), .A3(new_n393), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n392), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n391), .B1(new_n403), .B2(new_n221), .ZN(new_n404));
  INV_X1    g0204(.A(new_n392), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT76), .A3(G68), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n409), .A3(new_n388), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n390), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n289), .A2(new_n312), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n279), .A2(G1698), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n288), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n273), .B1(new_n417), .B2(KEYINPUT77), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT77), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n276), .B1(new_n278), .B2(new_n311), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(G200), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI211_X1 g0224(.A(G190), .B(new_n422), .C1(new_n418), .C2(new_n420), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n255), .B1(new_n208), .B2(G20), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n267), .A2(new_n428), .B1(new_n265), .B2(new_n255), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n412), .A2(new_n426), .A3(new_n427), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n424), .A2(new_n425), .ZN(new_n433));
  INV_X1    g0233(.A(new_n388), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n408), .A2(G68), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n391), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT16), .B1(new_n436), .B2(new_n409), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n429), .B(new_n433), .C1(new_n437), .C2(new_n390), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n427), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n422), .B1(new_n418), .B2(new_n420), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G179), .ZN(new_n441));
  INV_X1    g0241(.A(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n412), .B2(new_n430), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n443), .C1(new_n412), .C2(new_n430), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n432), .A2(new_n439), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n378), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n281), .A2(new_n283), .A3(G257), .A4(G1698), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n281), .A2(new_n283), .A3(G250), .A4(new_n312), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G294), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n292), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n274), .A2(G1), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n292), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G264), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n456), .A2(new_n273), .A3(G274), .A4(new_n455), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n292), .A2(new_n453), .B1(new_n457), .B2(G264), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(KEYINPUT87), .A3(new_n459), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G169), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n454), .A2(new_n458), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT88), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(KEYINPUT88), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(G179), .A4(new_n459), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n281), .A2(new_n283), .A3(new_n209), .A4(G87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n288), .A2(new_n475), .A3(new_n209), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G20), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n209), .B2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT23), .A3(G20), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n472), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n477), .A2(new_n472), .A3(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT24), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n259), .C1(new_n489), .C2(new_n485), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n264), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT25), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n208), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n260), .A2(new_n264), .A3(new_n262), .A4(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n492), .B(KEYINPUT86), .C1(new_n482), .C2(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n466), .A2(new_n471), .B1(new_n490), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n490), .A2(new_n499), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n462), .A2(new_n464), .A3(new_n323), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT89), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT89), .A4(new_n323), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n469), .A2(new_n470), .A3(new_n459), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n303), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n500), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n281), .A2(new_n283), .A3(G238), .A4(new_n312), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n281), .A2(new_n283), .A3(G244), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n478), .C1(new_n512), .C2(new_n312), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n292), .ZN(new_n514));
  INV_X1    g0314(.A(G274), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n208), .A2(new_n515), .A3(G45), .ZN(new_n516));
  INV_X1    g0316(.A(G250), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n274), .B2(G1), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n273), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT79), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n273), .A2(KEYINPUT79), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT80), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n514), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n514), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n442), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n514), .A2(new_n523), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n514), .A2(new_n523), .A3(new_n524), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n295), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n288), .A2(new_n209), .A3(G68), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n209), .B1(new_n310), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G87), .B2(new_n206), .ZN(new_n535));
  INV_X1    g0335(.A(G97), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n256), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n259), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n347), .A2(new_n265), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(new_n540), .C1(new_n347), .C2(new_n494), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n527), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(G200), .B1(new_n525), .B2(new_n526), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n529), .A2(G190), .A3(new_n530), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n540), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT81), .ZN(new_n546));
  INV_X1    g0346(.A(G87), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n494), .B2(new_n547), .ZN(new_n548));
  OR3_X1    g0348(.A1(new_n494), .A2(new_n546), .A3(new_n547), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n543), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n542), .A2(new_n551), .A3(KEYINPUT82), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT82), .B1(new_n542), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n281), .A2(new_n283), .A3(G264), .A4(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n281), .A2(new_n283), .A3(G257), .A4(new_n312), .ZN(new_n556));
  INV_X1    g0356(.A(G303), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n288), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT83), .B1(new_n558), .B2(new_n292), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n456), .A2(new_n455), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(G270), .A3(new_n273), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n459), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(KEYINPUT83), .A3(new_n292), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n303), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G283), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n566), .B(new_n209), .C1(G33), .C2(new_n536), .ZN(new_n567));
  INV_X1    g0367(.A(G116), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G20), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n259), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT20), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n208), .A2(G13), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n569), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n568), .B1(new_n208), .B2(G33), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n333), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT84), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  INV_X1    g0379(.A(new_n577), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n558), .A2(KEYINPUT83), .A3(new_n292), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n581), .A2(new_n559), .A3(new_n562), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n579), .B(new_n580), .C1(new_n582), .C2(new_n303), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(G190), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n578), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n570), .B(KEYINPUT20), .ZN(new_n587));
  INV_X1    g0387(.A(new_n576), .ZN(new_n588));
  OAI21_X1  g0388(.A(G169), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n582), .A2(G179), .A3(new_n577), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n558), .A2(new_n292), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT83), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n562), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n564), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT21), .A3(G169), .A4(new_n577), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n590), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n459), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n560), .A2(G257), .A3(new_n273), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n457), .A2(KEYINPUT78), .A3(G257), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n312), .ZN(new_n605));
  INV_X1    g0405(.A(new_n512), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n566), .C1(new_n606), .C2(KEYINPUT4), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n288), .A2(G250), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n312), .B1(new_n608), .B2(KEYINPUT4), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n292), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n442), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n604), .A2(new_n610), .A3(new_n295), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n408), .A2(G107), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n482), .A2(KEYINPUT6), .A3(G97), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n536), .A2(new_n482), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n205), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n617), .B2(KEYINPUT6), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n614), .A2(new_n619), .B1(new_n217), .B2(new_n258), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n264), .A2(G97), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n494), .B2(new_n536), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n612), .B(new_n613), .C1(new_n620), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n611), .A2(G200), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n619), .B1(new_n403), .B2(new_n482), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n259), .ZN(new_n627));
  INV_X1    g0427(.A(new_n623), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n604), .A2(new_n610), .A3(G190), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n625), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n585), .A2(new_n598), .A3(new_n624), .A4(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n449), .A2(new_n510), .A3(new_n554), .A4(new_n631), .ZN(G372));
  NOR2_X1   g0432(.A1(new_n412), .A2(new_n430), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT17), .B1(new_n633), .B2(new_n433), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n431), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n339), .A2(new_n377), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n338), .B2(new_n345), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n445), .A2(KEYINPUT91), .A3(new_n447), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT91), .B1(new_n445), .B2(new_n447), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n636), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n307), .A2(new_n308), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n296), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n542), .A2(new_n551), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT82), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n542), .A2(new_n551), .A3(KEYINPUT82), .ZN(new_n647));
  INV_X1    g0447(.A(new_n624), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n646), .A2(KEYINPUT26), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n528), .A2(new_n442), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n531), .A2(new_n541), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n528), .A2(G200), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n544), .A2(new_n550), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n650), .B1(new_n655), .B2(new_n624), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n612), .A2(new_n613), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n627), .A2(new_n628), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n659), .A2(new_n652), .A3(new_n654), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(KEYINPUT90), .A3(new_n650), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n649), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n624), .A2(new_n630), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n509), .A2(new_n502), .ZN(new_n666));
  INV_X1    g0466(.A(new_n655), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n590), .A2(new_n591), .A3(new_n597), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n500), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n652), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n449), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n643), .A2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  INV_X1    g0476(.A(G213), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n585), .B(new_n598), .C1(new_n580), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n669), .A2(new_n577), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n501), .A2(new_n681), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n510), .A2(new_n687), .B1(new_n500), .B2(new_n681), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n598), .A2(new_n681), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n510), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n500), .A2(new_n682), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  INV_X1    g0497(.A(new_n212), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(G41), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n212), .A2(KEYINPUT93), .A3(new_n272), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n215), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT96), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n594), .A2(G179), .A3(new_n595), .A4(new_n564), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT94), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n563), .A2(KEYINPUT94), .A3(G179), .A4(new_n564), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n469), .A2(new_n470), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n525), .A2(new_n526), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(new_n610), .A4(new_n604), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n707), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n710), .A2(new_n711), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n611), .A2(new_n526), .A3(new_n525), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n718), .A4(new_n713), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n596), .A2(new_n295), .A3(new_n528), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT95), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n507), .A2(new_n721), .A3(new_n611), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n507), .B2(new_n611), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n716), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n681), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n706), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n681), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(KEYINPUT96), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n631), .A2(new_n554), .A3(new_n510), .A4(new_n682), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n646), .A2(new_n650), .A3(new_n647), .A4(new_n648), .ZN(new_n737));
  INV_X1    g0537(.A(new_n652), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n466), .A2(new_n471), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n501), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n598), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT97), .B1(new_n500), .B2(new_n669), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n737), .B(new_n739), .C1(new_n745), .C2(new_n668), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT29), .A3(new_n682), .ZN(new_n747));
  INV_X1    g0547(.A(new_n671), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n681), .B1(new_n748), .B2(new_n663), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n749), .B2(KEYINPUT29), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n736), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n705), .B1(new_n751), .B2(G1), .ZN(G364));
  XNOR2_X1  g0552(.A(new_n686), .B(KEYINPUT98), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n701), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n209), .A2(G13), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G45), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n208), .B1(new_n757), .B2(KEYINPUT99), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n754), .B(new_n762), .C1(G330), .C2(new_n685), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n212), .A2(new_n288), .ZN(new_n764));
  INV_X1    g0564(.A(G355), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n765), .B1(G116), .B2(new_n212), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n288), .B(new_n698), .C1(new_n274), .C2(new_n216), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n242), .A2(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT100), .Z(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n217), .B1(G20), .B2(new_n442), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n761), .B1(new_n769), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n209), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n323), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n482), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n209), .A2(new_n295), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n221), .B1(new_n786), .B2(new_n547), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n783), .A2(new_n323), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n781), .B(new_n787), .C1(G50), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n303), .A2(G190), .ZN(new_n790));
  OAI21_X1  g0590(.A(G20), .B1(new_n790), .B2(G179), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT101), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G97), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G190), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n779), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n782), .A2(new_n798), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n288), .B1(new_n803), .B2(new_n287), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n790), .A2(new_n209), .A3(new_n295), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G58), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n789), .A2(new_n797), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n795), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n788), .ZN(new_n810));
  INV_X1    g0610(.A(G326), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(new_n786), .B2(new_n557), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n785), .A2(new_n813), .B1(new_n780), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n288), .B1(new_n805), .B2(G322), .ZN(new_n817));
  INV_X1    g0617(.A(new_n803), .ZN(new_n818));
  INV_X1    g0618(.A(new_n799), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G311), .A2(new_n818), .B1(new_n819), .B2(G329), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n807), .B1(new_n809), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n778), .B1(new_n822), .B2(new_n775), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n685), .B2(new_n773), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n763), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n377), .A2(KEYINPUT105), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n373), .A2(new_n374), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n442), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT105), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n829), .A2(new_n830), .A3(new_n376), .A4(new_n375), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n372), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n682), .B(new_n832), .C1(new_n664), .C2(new_n671), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n376), .A2(new_n681), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n372), .A2(new_n834), .A3(new_n827), .A4(new_n831), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n377), .A2(new_n682), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n749), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n761), .B1(new_n736), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n736), .B2(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(new_n775), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n771), .ZN(new_n842));
  INV_X1    g0642(.A(new_n805), .ZN(new_n843));
  INV_X1    g0643(.A(G311), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n843), .A2(new_n808), .B1(new_n799), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n780), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G87), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n810), .B2(new_n557), .C1(new_n814), .C2(new_n785), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n845), .B(new_n848), .C1(G116), .C2(new_n818), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n284), .B1(new_n786), .B2(new_n482), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT102), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n849), .A2(new_n797), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n818), .A2(G159), .B1(new_n805), .B2(G143), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n810), .B2(new_n854), .C1(new_n248), .C2(new_n785), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT34), .Z(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n780), .A2(new_n221), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n288), .B1(new_n799), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n786), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n859), .B(new_n861), .C1(G50), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n202), .B2(new_n795), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n856), .B2(new_n857), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n852), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n761), .B1(G77), .B2(new_n842), .C1(new_n866), .C2(new_n841), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT104), .Z(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n771), .B2(new_n837), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n840), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  NAND2_X1  g0671(.A1(new_n389), .A2(new_n263), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n386), .B2(new_n388), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n429), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n679), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT107), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n448), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n443), .A2(new_n874), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n438), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT108), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n438), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n875), .B1(new_n412), .B2(new_n430), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n444), .A2(new_n438), .A3(new_n887), .A4(new_n880), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n879), .C1(new_n886), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n438), .A2(new_n444), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n888), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n894));
  INV_X1    g0694(.A(new_n887), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n890), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT109), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n338), .A2(new_n681), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n346), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n338), .B(new_n681), .C1(new_n345), .C2(new_n339), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND4_X1   g0703(.A1(KEYINPUT40), .A2(new_n899), .A3(new_n837), .A4(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n898), .B1(new_n897), .B2(new_n904), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n412), .A2(new_n430), .A3(new_n426), .ZN(new_n908));
  INV_X1    g0708(.A(new_n881), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n883), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n876), .B(KEYINPUT107), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n885), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n889), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n445), .A2(new_n447), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n911), .B1(new_n914), .B2(new_n635), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n907), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n890), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n899), .A2(new_n837), .A3(new_n903), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT40), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n905), .A2(new_n906), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n449), .A2(new_n899), .ZN(new_n922));
  OAI21_X1  g0722(.A(G330), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n921), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n897), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n345), .A2(new_n338), .A3(new_n682), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n916), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n903), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n827), .A2(new_n831), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT106), .B1(new_n932), .B2(new_n682), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n934), .B(new_n681), .C1(new_n827), .C2(new_n831), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n931), .B1(new_n833), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n639), .A2(new_n640), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n937), .A2(new_n917), .B1(new_n938), .B2(new_n679), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n449), .B(new_n747), .C1(new_n749), .C2(KEYINPUT29), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(new_n643), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n924), .A2(new_n943), .B1(new_n208), .B2(new_n756), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n924), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n618), .A2(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n618), .A2(KEYINPUT35), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(G116), .A3(new_n218), .A4(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT36), .Z(new_n949));
  OAI211_X1 g0749(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n221), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n201), .A2(G68), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n208), .B(G13), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n945), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT110), .Z(G367));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n624), .A2(new_n682), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT111), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n660), .A2(new_n681), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n665), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n955), .B1(new_n962), .B2(new_n694), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n695), .A2(new_n961), .A3(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n694), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT44), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n695), .B2(new_n961), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n689), .ZN(new_n971));
  INV_X1    g0771(.A(new_n688), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n692), .B1(new_n972), .B2(new_n691), .ZN(new_n973));
  MUX2_X1   g0773(.A(new_n686), .B(new_n753), .S(new_n973), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n751), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n751), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n701), .B(KEYINPUT41), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n760), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT112), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n961), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n741), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n682), .B1(new_n985), .B2(new_n648), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n962), .A2(new_n692), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n550), .A2(new_n682), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n655), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n738), .A2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT113), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n982), .A2(new_n984), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n690), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n986), .A2(new_n988), .A3(new_n995), .A4(new_n994), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n998), .A2(new_n1002), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n981), .A2(new_n1003), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n347), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n777), .B1(new_n698), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n698), .A2(new_n288), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n238), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n762), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n819), .A2(G317), .B1(new_n805), .B2(G303), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n284), .C1(new_n814), .C2(new_n803), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n788), .A2(G311), .B1(new_n846), .B2(G97), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n808), .B2(new_n785), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT46), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n862), .A2(G116), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1016), .B(new_n1018), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1019), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT114), .Z(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n482), .C2(new_n795), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT115), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n803), .A2(new_n201), .B1(new_n799), .B2(new_n854), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n284), .B(new_n1026), .C1(G150), .C2(new_n805), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n796), .A2(G68), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n780), .A2(new_n287), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G159), .B2(new_n784), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n788), .A2(G143), .B1(new_n862), .B2(G58), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT47), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n1014), .B1(new_n773), .B2(new_n993), .C1(new_n1034), .C2(new_n841), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1009), .A2(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n975), .A2(new_n755), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(KEYINPUT117), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n751), .A2(new_n974), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT118), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n284), .B1(new_n799), .B2(new_n811), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n818), .A2(G303), .B1(new_n805), .B2(G317), .ZN(new_n1045));
  INV_X1    g0845(.A(G322), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1045), .B1(new_n810), .B2(new_n1046), .C1(new_n844), .C2(new_n785), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n796), .A2(G283), .B1(G294), .B2(new_n862), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT49), .Z(new_n1053));
  AOI211_X1 g0853(.A(new_n1044), .B(new_n1053), .C1(G116), .C2(new_n846), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n795), .A2(new_n347), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n284), .B1(new_n805), .B2(G50), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n221), .B2(new_n803), .C1(new_n248), .C2(new_n799), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n810), .A2(new_n800), .B1(new_n780), .B2(new_n536), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n785), .A2(new_n255), .B1(new_n786), .B2(new_n287), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n775), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n235), .A2(G45), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n349), .A2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n274), .B1(new_n221), .B2(new_n287), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n702), .B2(KEYINPUT116), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(KEYINPUT116), .C2(new_n702), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1062), .A2(new_n1012), .A3(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(G107), .B2(new_n212), .C1(new_n702), .C2(new_n764), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n762), .B1(new_n1069), .B2(new_n776), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n688), .B2(new_n774), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n974), .B2(new_n760), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1043), .A2(new_n1073), .ZN(G393));
  AND3_X1   g0874(.A1(new_n971), .A2(KEYINPUT120), .A3(new_n975), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT120), .B1(new_n971), .B2(new_n975), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n755), .B1(new_n975), .B2(new_n971), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n971), .A2(new_n980), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1012), .A2(new_n245), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n776), .B1(new_n536), .B2(new_n212), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n788), .A2(G150), .B1(G159), .B2(new_n805), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT51), .Z(new_n1082));
  INV_X1    g0882(.A(G143), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n288), .B1(new_n799), .B2(new_n1083), .C1(new_n349), .C2(new_n803), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n847), .B1(new_n221), .B2(new_n786), .C1(new_n785), .C2(new_n201), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G77), .C2(new_n796), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n788), .A2(G317), .B1(G311), .B2(new_n805), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G116), .B2(new_n796), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n284), .B1(new_n799), .B2(new_n1046), .C1(new_n808), .C2(new_n803), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n785), .A2(new_n557), .B1(new_n780), .B2(new_n482), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G283), .C2(new_n862), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1082), .A2(new_n1086), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n761), .B1(new_n1079), .B2(new_n1080), .C1(new_n1094), .C2(new_n841), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1000), .B2(new_n774), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1078), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1077), .A2(new_n1097), .ZN(G390));
  AND4_X1   g0898(.A1(G330), .A2(new_n899), .A3(new_n837), .A4(new_n903), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n937), .A2(new_n928), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n926), .B2(new_n929), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n746), .A2(new_n682), .A3(new_n832), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n936), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n903), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n897), .A2(new_n927), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1099), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n903), .A2(new_n837), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n735), .A2(new_n1108), .A3(G330), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n916), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n925), .B2(new_n897), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1105), .C1(new_n1111), .C2(new_n1100), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n449), .A2(G330), .A3(new_n899), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n941), .A2(new_n643), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n899), .A2(G330), .A3(new_n837), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1103), .B1(new_n931), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1109), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT121), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1117), .A2(KEYINPUT121), .A3(new_n1109), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n833), .A2(new_n936), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n735), .A2(G330), .A3(new_n837), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n931), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1099), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1115), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1113), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1099), .B1(new_n1125), .B2(new_n931), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1120), .B(new_n1121), .C1(new_n1124), .C2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1107), .A2(new_n1132), .A3(new_n1112), .A4(new_n1115), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n755), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1107), .A2(new_n760), .A3(new_n1112), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n255), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n761), .B1(new_n1136), .B2(new_n842), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n482), .A2(new_n785), .B1(new_n810), .B2(new_n814), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n859), .B(new_n1138), .C1(G87), .C2(new_n862), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n803), .A2(new_n536), .B1(new_n799), .B2(new_n808), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n288), .B(new_n1140), .C1(G116), .C2(new_n805), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n287), .C2(new_n795), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n284), .B1(new_n819), .B2(G125), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n201), .B2(new_n780), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT122), .Z(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n818), .A2(new_n1147), .B1(new_n805), .B2(G132), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n810), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G137), .B2(new_n784), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n786), .A2(new_n248), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n800), .C2(new_n795), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1142), .B1(new_n1145), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1137), .B1(new_n1155), .B2(new_n775), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1111), .B2(new_n771), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1134), .A2(new_n1135), .A3(new_n1157), .ZN(G378));
  NAND3_X1  g0958(.A1(new_n920), .A2(G330), .A3(new_n940), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n937), .A2(new_n917), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n938), .A2(new_n679), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1111), .B2(new_n928), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n897), .A2(new_n904), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT109), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n917), .A2(new_n918), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT40), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1165), .A2(G330), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1163), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n270), .A2(new_n875), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n309), .B(new_n1172), .Z(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1173), .B(new_n1174), .Z(new_n1175));
  AND3_X1   g0975(.A1(new_n1159), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1159), .B2(new_n1171), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n760), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n761), .B1(G50), .B2(new_n842), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n284), .B2(new_n272), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n843), .A2(new_n482), .B1(new_n347), .B2(new_n803), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n272), .B(new_n284), .C1(new_n799), .C2(new_n814), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n780), .A2(new_n202), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G77), .B2(new_n862), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n784), .A2(G97), .B1(new_n788), .B2(G116), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1028), .A2(new_n1184), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n843), .A2(new_n1149), .B1(new_n803), .B2(new_n854), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n862), .B2(new_n1147), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n784), .A2(G132), .B1(new_n788), .B2(G125), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n248), .C2(new_n795), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n846), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n819), .C2(G124), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1190), .B1(new_n1189), .B2(new_n1188), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1179), .B1(new_n1200), .B2(new_n775), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1175), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n771), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1178), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n940), .B1(new_n920), .B2(G330), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1163), .A2(new_n1170), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1159), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1207), .A2(new_n1208), .B1(new_n1115), .B2(new_n1133), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n755), .B1(new_n1209), .B2(KEYINPUT57), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1133), .A2(new_n1115), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(KEYINPUT57), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1204), .B1(new_n1210), .B2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n931), .A2(new_n770), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n761), .B1(G68), .B2(new_n842), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n810), .A2(new_n860), .B1(new_n786), .B2(new_n800), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1185), .B(new_n1217), .C1(new_n784), .C2(new_n1147), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n843), .A2(new_n854), .B1(new_n799), .B2(new_n1149), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n284), .B(new_n1219), .C1(G150), .C2(new_n818), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n201), .C2(new_n795), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n843), .A2(new_n814), .B1(new_n799), .B2(new_n557), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n288), .B(new_n1222), .C1(G107), .C2(new_n818), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1029), .B1(G294), .B2(new_n788), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n784), .A2(G116), .B1(new_n862), .B2(G97), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1221), .B1(new_n1055), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1216), .B1(new_n1227), .B2(new_n775), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1132), .A2(new_n760), .B1(new_n1215), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1129), .A2(new_n978), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1117), .A2(KEYINPUT121), .A3(new_n1109), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT121), .B1(new_n1117), .B2(new_n1109), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1128), .A2(new_n1231), .A3(new_n1232), .A4(new_n1115), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1230), .B2(new_n1233), .ZN(G381));
  NAND4_X1  g1034(.A1(new_n1009), .A2(new_n1035), .A3(new_n1077), .A4(new_n1097), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1043), .A2(new_n825), .A3(new_n870), .A4(new_n1073), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1235), .A2(G381), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1178), .A2(new_n1203), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1211), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT57), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n701), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1238), .B1(new_n1241), .B2(new_n1212), .ZN(new_n1242));
  INV_X1    g1042(.A(G378), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1237), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1237), .A2(new_n1242), .A3(KEYINPUT123), .A4(new_n1243), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(G407));
  NOR2_X1   g1048(.A1(G375), .A2(G378), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n677), .A2(G343), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT124), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n677), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G407), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(KEYINPUT125), .A3(new_n1252), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(G409));
  OAI211_X1 g1057(.A(G378), .B(new_n1204), .C1(new_n1210), .C2(new_n1213), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1178), .B(new_n1203), .C1(new_n1239), .C2(new_n977), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1243), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1250), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1132), .B2(new_n1115), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n701), .B1(new_n1132), .B2(new_n1115), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1123), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1115), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(KEYINPUT60), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT126), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1128), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(KEYINPUT60), .A4(new_n1270), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1266), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1277), .B2(new_n1229), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1229), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n870), .B(new_n1279), .C1(new_n1266), .C2(new_n1276), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1261), .A2(new_n1262), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1251), .A2(G2897), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n755), .B(new_n1129), .C1(new_n1233), .C2(KEYINPUT60), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1275), .B2(new_n1272), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n870), .B1(new_n1288), .B2(new_n1279), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1277), .A2(G384), .A3(new_n1229), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1286), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1250), .A2(G2897), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1278), .A2(new_n1280), .A3(new_n1292), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1285), .A2(new_n1250), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1235), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(new_n825), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(G396), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1295), .A3(new_n1235), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(KEYINPUT61), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1251), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1281), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1284), .A2(new_n1294), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1293), .A2(new_n1291), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1303), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1282), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1303), .A2(KEYINPUT62), .A3(new_n1281), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1301), .B(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1305), .B1(new_n1312), .B2(new_n1314), .ZN(G405));
  NOR2_X1   g1115(.A1(new_n1242), .A2(G378), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1258), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1281), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G375), .A2(new_n1243), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1319), .B(new_n1258), .C1(new_n1278), .C2(new_n1280), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(new_n1301), .ZN(G402));
endmodule


