//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n202), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n201), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G68), .A2(G238), .ZN(new_n222));
  NOR4_X1   g0022(.A1(new_n217), .A2(new_n219), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT64), .B(G77), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n223), .A2(new_n225), .B1(G1), .B2(G20), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n208), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n211), .B(new_n227), .C1(new_n229), .C2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(new_n207), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n201), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(new_n228), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n228), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n208), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n261), .A2(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(G20), .B2(new_n204), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n256), .A2(new_n269), .A3(new_n259), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n250), .A3(new_n270), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n253), .B1(new_n260), .B2(new_n267), .C1(new_n271), .C2(new_n201), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G223), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G222), .B2(G1698), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n224), .B2(new_n280), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT66), .A3(G274), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n207), .B(G274), .C1(G41), .C2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(new_n284), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n282), .B(new_n289), .C1(new_n220), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT73), .A3(G200), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n292), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT73), .B1(new_n292), .B2(G200), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT10), .B1(new_n297), .B2(KEYINPUT72), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n289), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n280), .A2(G232), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n305), .B(new_n306), .C1(new_n215), .C2(new_n280), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n303), .B1(new_n307), .B2(new_n290), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n290), .A2(new_n284), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G244), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n255), .A2(G77), .A3(new_n250), .ZN(new_n314));
  INV_X1    g0114(.A(new_n261), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n264), .B1(new_n224), .B2(G20), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n262), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n314), .B1(new_n319), .B2(new_n257), .ZN(new_n320));
  INV_X1    g0120(.A(new_n224), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n252), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n308), .A2(new_n324), .A3(new_n310), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n313), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n302), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n280), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT7), .A2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT80), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G33), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n337));
  AOI21_X1  g0137(.A(G20), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  OAI211_X1 g0139(.A(G68), .B(new_n331), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(G58), .B(G68), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(G20), .B1(G159), .B2(new_n264), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n255), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n335), .B1(new_n332), .B2(new_n334), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n335), .A2(G33), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT81), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT81), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT80), .B(G33), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n347), .C1(new_n351), .C2(new_n335), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n330), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n332), .A2(new_n334), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n354), .B2(KEYINPUT3), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT7), .B1(new_n355), .B2(G20), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(G68), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT16), .A3(new_n342), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n345), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n271), .A2(new_n315), .ZN(new_n360));
  INV_X1    g0160(.A(new_n252), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n261), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n277), .A2(new_n304), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n347), .B(new_n366), .C1(new_n351), .C2(new_n335), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n304), .A2(G226), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n290), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n291), .A2(new_n218), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n372), .A3(new_n289), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n324), .B2(new_n373), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n364), .A2(KEYINPUT18), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n345), .A2(new_n358), .B1(new_n362), .B2(new_n360), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n303), .B1(new_n369), .B2(new_n290), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n312), .B1(new_n379), .B2(new_n372), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n333), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT3), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n368), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(new_n347), .A3(new_n366), .A4(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n276), .B1(new_n385), .B2(new_n365), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n386), .A2(new_n324), .A3(new_n371), .A4(new_n303), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n377), .B1(new_n378), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n376), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(G190), .A3(new_n372), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n373), .A2(G200), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n359), .A2(new_n363), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT17), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n378), .A2(KEYINPUT17), .A3(new_n391), .A4(new_n392), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n292), .A2(G179), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT69), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n292), .A2(new_n312), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n272), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT70), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT70), .B1(new_n399), .B2(new_n402), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n390), .A2(new_n397), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n220), .A2(new_n304), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n218), .A2(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n347), .A2(new_n407), .A3(new_n337), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT74), .B1(new_n411), .B2(new_n290), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n413), .B(new_n276), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n309), .A2(G238), .B1(new_n285), .B2(new_n288), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n406), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G226), .A2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n218), .B2(G1698), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n280), .B1(G33), .B2(G97), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n413), .B1(new_n420), .B2(new_n276), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n411), .A2(KEYINPUT74), .A3(new_n290), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n416), .A4(new_n406), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G200), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n416), .A3(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT13), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(G190), .A3(new_n423), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n250), .A2(new_n254), .A3(G68), .A4(new_n228), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT75), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n255), .A2(new_n431), .A3(G68), .A4(new_n250), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n207), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT12), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT12), .B1(new_n433), .B2(new_n434), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n430), .B(new_n432), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT77), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n435), .B(new_n436), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n429), .B(new_n431), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n208), .A2(G33), .A3(G77), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n446), .B1(new_n208), .B2(G68), .C1(new_n265), .C2(new_n201), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n256), .A3(new_n259), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT11), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n445), .B2(new_n449), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n425), .B(new_n428), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n445), .A2(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n428), .A4(new_n425), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT14), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n427), .A2(new_n423), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G169), .ZN(new_n463));
  AOI211_X1 g0263(.A(KEYINPUT14), .B(new_n312), .C1(new_n427), .C2(new_n423), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n324), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n454), .B(new_n460), .C1(new_n466), .C2(new_n458), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n311), .A2(G200), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT71), .A3(new_n322), .A4(new_n320), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT71), .ZN(new_n471));
  INV_X1    g0271(.A(G200), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n308), .B2(new_n310), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n323), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n470), .B(new_n474), .C1(new_n294), .C2(new_n311), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n328), .A2(new_n405), .A3(new_n468), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  INV_X1    g0277(.A(G87), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G20), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n347), .B(new_n479), .C1(new_n351), .C2(new_n335), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT86), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n383), .A2(KEYINPUT86), .A3(new_n347), .A4(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(KEYINPUT22), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n280), .A2(new_n485), .A3(new_n479), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n354), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n208), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT87), .B1(new_n215), .B2(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n477), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  AOI211_X1 g0296(.A(KEYINPUT24), .B(new_n494), .C1(new_n484), .C2(new_n486), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n257), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT88), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(KEYINPUT88), .B(new_n257), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n252), .A2(new_n215), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT25), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n207), .A2(G33), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n260), .A2(new_n361), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n507), .B2(G107), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n214), .A2(G1698), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n355), .B(new_n510), .C1(G250), .C2(G1698), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n351), .A2(G294), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n276), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G41), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n515), .A2(new_n517), .A3(new_n207), .A4(G45), .ZN(new_n518));
  INV_X1    g0318(.A(G274), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n276), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(KEYINPUT90), .A3(G264), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT90), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n521), .B2(new_n216), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n520), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n514), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n513), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n526), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(G169), .B1(new_n531), .B2(G179), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n509), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n252), .A2(new_n213), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n507), .A2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  OAI211_X1 g0337(.A(G107), .B(new_n331), .C1(new_n338), .C2(new_n339), .ZN(new_n538));
  INV_X1    g0338(.A(G77), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n265), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n213), .A2(new_n215), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n546), .B2(G20), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n537), .B1(new_n548), .B2(new_n257), .ZN(new_n549));
  AOI211_X1 g0349(.A(KEYINPUT82), .B(new_n255), .C1(new_n538), .C2(new_n547), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n535), .B(new_n536), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n383), .A2(G244), .A3(new_n304), .A4(new_n347), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n347), .A2(new_n337), .A3(G250), .A4(G1698), .ZN(new_n555));
  AND2_X1   g0355(.A1(KEYINPUT4), .A2(G244), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n347), .A2(new_n337), .A3(new_n556), .A4(new_n304), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n290), .ZN(new_n562));
  INV_X1    g0362(.A(new_n520), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n522), .A2(G257), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n562), .A2(new_n324), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n559), .B1(new_n552), .B2(new_n553), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n563), .B(new_n564), .C1(new_n566), .C2(new_n276), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n312), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n551), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n562), .A2(new_n294), .A3(new_n563), .A4(new_n564), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n472), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n255), .B1(new_n538), .B2(new_n547), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(new_n537), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n572), .A2(new_n574), .A3(new_n535), .A4(new_n536), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n207), .A2(G45), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n276), .A2(G250), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT83), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n276), .A2(new_n579), .A3(G250), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n576), .A2(new_n519), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G238), .A2(G1698), .ZN(new_n584));
  INV_X1    g0384(.A(G244), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(G1698), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n489), .B1(new_n355), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n581), .B(new_n583), .C1(new_n587), .C2(new_n276), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n203), .A2(G20), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n347), .B(new_n589), .C1(new_n351), .C2(new_n335), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n208), .B1(new_n410), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n543), .A2(new_n478), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n262), .B2(new_n213), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT84), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT84), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n591), .C1(new_n262), .C2(new_n213), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n590), .A2(new_n594), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n257), .B1(new_n252), .B2(new_n318), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n260), .A2(new_n361), .A3(new_n317), .A4(new_n505), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n312), .A2(new_n588), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n588), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n324), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n351), .A2(G116), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n347), .B1(new_n351), .B2(new_n335), .ZN(new_n607));
  INV_X1    g0407(.A(new_n586), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n582), .B1(new_n609), .B2(new_n290), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n472), .B1(new_n610), .B2(new_n581), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n260), .A2(G87), .A3(new_n361), .A4(new_n505), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n600), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT85), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n603), .A2(G190), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n588), .A2(G200), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n600), .A4(new_n612), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n569), .A2(new_n575), .A3(new_n605), .A4(new_n619), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n528), .A2(G190), .B1(new_n531), .B2(G200), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n502), .A2(new_n508), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n214), .A2(new_n304), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n355), .B(new_n623), .C1(G264), .C2(new_n304), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n329), .A2(G303), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n276), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n522), .A2(G270), .ZN(new_n627));
  OR3_X1    g0427(.A1(new_n626), .A2(new_n520), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n361), .A2(G116), .A3(new_n255), .A4(new_n505), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n558), .B(new_n208), .C1(G33), .C2(new_n213), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n257), .C1(new_n208), .C2(G116), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT20), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI221_X1 g0434(.A(new_n629), .B1(G116), .B2(new_n361), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(G169), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n626), .A2(new_n520), .A3(new_n627), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(G179), .A3(new_n635), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n628), .A2(KEYINPUT21), .A3(G169), .A4(new_n635), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(G190), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n472), .B2(new_n639), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n635), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n534), .A2(new_n620), .A3(new_n622), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n476), .A2(new_n647), .ZN(G372));
  NOR2_X1   g0448(.A1(new_n403), .A2(new_n404), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n453), .A2(new_n327), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n466), .B2(new_n458), .ZN(new_n651));
  INV_X1    g0451(.A(new_n397), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n390), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(new_n302), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n565), .A2(new_n568), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n619), .A2(new_n551), .A3(new_n656), .A4(new_n605), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n611), .A2(new_n613), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(new_n615), .B1(new_n602), .B2(new_n604), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n551), .A4(new_n656), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n605), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n642), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n534), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n575), .A2(new_n569), .A3(new_n660), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n622), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n655), .B1(new_n476), .B2(new_n668), .ZN(G369));
  AND2_X1   g0469(.A1(new_n534), .A2(new_n622), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n251), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n207), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n509), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n532), .B1(new_n502), .B2(new_n508), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT91), .B(G330), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n635), .A2(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n646), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n664), .B2(new_n684), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n682), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n664), .A2(new_n677), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n670), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n677), .B(KEYINPUT92), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n209), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G1), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n543), .A2(new_n478), .A3(new_n488), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n231), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n668), .B2(new_n690), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n642), .B1(new_n509), .B2(new_n533), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n622), .A2(new_n666), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(KEYINPUT93), .B(new_n691), .C1(new_n707), .C2(new_n663), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n628), .A2(new_n530), .A3(new_n324), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n603), .A2(new_n564), .A3(new_n562), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n710), .B2(new_n712), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n530), .A2(new_n324), .A3(new_n567), .A4(new_n588), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n714), .A2(new_n715), .B1(new_n639), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n716), .A2(new_n639), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n710), .A2(new_n712), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n722), .B2(new_n713), .ZN(new_n723));
  INV_X1    g0523(.A(new_n677), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n718), .B(new_n725), .C1(new_n647), .C2(new_n690), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n683), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n657), .A2(new_n661), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT94), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT94), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n657), .A2(new_n730), .A3(new_n661), .ZN(new_n731));
  INV_X1    g0531(.A(new_n569), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT26), .A3(new_n660), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n622), .B(new_n666), .C1(new_n680), .C2(new_n642), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n605), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n724), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n709), .A2(new_n727), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n701), .B1(new_n740), .B2(G1), .ZN(G364));
  OR2_X1    g0541(.A1(new_n686), .A2(new_n683), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n686), .A2(new_n683), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n698), .B1(G45), .B2(new_n671), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n208), .B1(new_n747), .B2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(G20), .A2(G179), .A3(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n472), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n749), .A2(G294), .B1(G326), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n208), .A2(G190), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G179), .A3(G200), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT33), .B(G317), .Z(new_n755));
  OAI211_X1 g0555(.A(new_n752), .B(new_n329), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n472), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G20), .A3(new_n294), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n753), .A2(new_n747), .ZN(new_n760));
  INV_X1    g0560(.A(G329), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT96), .Z(new_n763));
  NOR2_X1   g0563(.A1(new_n750), .A2(G200), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n756), .B(new_n763), .C1(G322), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G303), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n757), .A2(G20), .A3(G190), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n753), .A2(G179), .A3(new_n472), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(G311), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT97), .Z(new_n772));
  INV_X1    g0572(.A(new_n751), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n201), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n764), .B(KEYINPUT95), .ZN(new_n775));
  INV_X1    g0575(.A(new_n758), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n775), .A2(G58), .B1(G107), .B2(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n777), .B1(new_n203), .B2(new_n754), .C1(new_n321), .C2(new_n769), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n760), .A2(KEYINPUT32), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n778), .A2(new_n329), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n767), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G87), .B1(new_n749), .B2(G97), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT32), .B1(new_n760), .B2(new_n779), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n772), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n228), .B1(G20), .B2(new_n312), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n787), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n280), .A2(new_n209), .A3(G355), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n349), .A2(new_n352), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n695), .ZN(new_n794));
  INV_X1    g0594(.A(new_n245), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n283), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n231), .A2(G45), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n792), .B1(G116), .B2(new_n209), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n786), .A2(new_n787), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n790), .B(KEYINPUT98), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n686), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n746), .B1(new_n802), .B2(new_n745), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n323), .A2(new_n677), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n475), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n326), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n327), .A2(new_n724), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n658), .A2(new_n605), .A3(new_n662), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n690), .B(new_n808), .C1(new_n735), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n703), .A2(new_n708), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n808), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(new_n727), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n745), .ZN(new_n814));
  INV_X1    g0614(.A(new_n754), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G150), .B1(new_n770), .B2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  INV_X1    g0617(.A(new_n775), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n816), .B1(new_n817), .B2(new_n773), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT100), .Z(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  INV_X1    g0622(.A(new_n793), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n767), .A2(new_n201), .B1(new_n748), .B2(new_n202), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n758), .A2(new_n203), .B1(new_n760), .B2(new_n825), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n815), .A2(G283), .B1(new_n770), .B2(G116), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n766), .B2(new_n773), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT99), .Z(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G294), .B2(new_n764), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n776), .A2(G87), .B1(new_n749), .B2(G97), .ZN(new_n832));
  INV_X1    g0632(.A(new_n760), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n280), .B1(new_n833), .B2(G311), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G107), .B2(new_n782), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n787), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n787), .A2(new_n788), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n539), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n744), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT101), .ZN(new_n841));
  INV_X1    g0641(.A(new_n808), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n789), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n814), .A2(new_n843), .ZN(G384));
  INV_X1    g0644(.A(KEYINPUT40), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n725), .C1(new_n647), .C2(new_n690), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n458), .A2(new_n724), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT103), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n463), .A2(new_n464), .ZN(new_n851));
  INV_X1    g0651(.A(new_n465), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n458), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n466), .A2(KEYINPUT103), .A3(new_n458), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n453), .B(new_n849), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n467), .A2(new_n858), .A3(new_n848), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n467), .B2(new_n848), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n847), .A2(new_n861), .A3(new_n842), .ZN(new_n862));
  INV_X1    g0662(.A(new_n675), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n357), .A2(new_n342), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n260), .B1(new_n864), .B2(new_n344), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n358), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n363), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n863), .B(new_n867), .C1(new_n390), .C2(new_n397), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n866), .A2(new_n363), .B1(new_n388), .B2(new_n675), .ZN(new_n869));
  INV_X1    g0669(.A(new_n393), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n364), .B1(new_n375), .B2(new_n863), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n393), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n845), .B1(new_n862), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n364), .B(new_n863), .C1(new_n390), .C2(new_n397), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n872), .A2(new_n393), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n874), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n845), .B1(new_n888), .B2(new_n879), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n889), .A2(new_n842), .A3(new_n847), .A4(new_n861), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n847), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n476), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n891), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n683), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n709), .A2(new_n738), .ZN(new_n896));
  INV_X1    g0696(.A(new_n476), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n654), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n895), .B(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n390), .A2(new_n675), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n849), .A2(new_n453), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n458), .B1(new_n851), .B2(new_n852), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n850), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT103), .B1(new_n466), .B2(new_n458), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n454), .A2(new_n460), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n848), .B1(new_n908), .B2(new_n904), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n467), .A2(new_n858), .A3(new_n848), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n691), .B(new_n842), .C1(new_n707), .C2(new_n663), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(new_n807), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n902), .B1(new_n914), .B2(new_n880), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n887), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n855), .A2(new_n856), .A3(new_n677), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n900), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n807), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n880), .B(new_n861), .C1(new_n810), .C2(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n924), .A2(new_n921), .A3(new_n900), .A4(new_n901), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT106), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n899), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n207), .B2(new_n671), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n488), .B1(new_n546), .B2(KEYINPUT35), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n229), .C1(KEYINPUT35), .C2(new_n546), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n232), .B1(new_n202), .B2(new_n203), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(new_n321), .B1(G50), .B2(new_n203), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n251), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT102), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n933), .A3(new_n937), .ZN(G367));
  NAND2_X1  g0738(.A1(new_n689), .A2(new_n692), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n732), .A2(new_n690), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n551), .A2(new_n690), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n575), .A2(new_n569), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n939), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT42), .B1(new_n689), .B2(new_n943), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(new_n569), .C2(new_n690), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n613), .A2(new_n677), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n660), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n605), .A2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT107), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n948), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT108), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n956), .A2(new_n959), .B1(new_n687), .B2(new_n943), .ZN(new_n960));
  INV_X1    g0760(.A(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(new_n687), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n961), .A2(new_n962), .A3(new_n944), .A4(new_n955), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n696), .B(new_n965), .Z(new_n966));
  NOR2_X1   g0766(.A1(new_n693), .A2(new_n944), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT44), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n939), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n693), .A2(new_n944), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT45), .B1(new_n693), .B2(new_n944), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n968), .A2(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n962), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n967), .B(KEYINPUT44), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n970), .B(new_n971), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n687), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT110), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n962), .A2(new_n980), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n743), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT111), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n687), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n985), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n739), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n981), .A2(new_n983), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n966), .B1(new_n991), .B2(new_n740), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n207), .B1(new_n671), .B2(G45), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n964), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n280), .B1(new_n321), .B2(new_n758), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n996), .A2(KEYINPUT113), .B1(G50), .B2(new_n770), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(KEYINPUT113), .B2(new_n996), .C1(new_n202), .C2(new_n767), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n754), .A2(new_n779), .B1(new_n760), .B2(new_n817), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n749), .A2(G68), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n773), .B2(new_n819), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n764), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n263), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n775), .A2(G303), .B1(G311), .B2(new_n751), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n793), .B(new_n1006), .C1(G107), .C2(new_n749), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n815), .A2(G294), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n770), .A2(G283), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n776), .A2(G97), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1007), .B(new_n1011), .C1(new_n1012), .C2(new_n760), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n767), .A2(new_n488), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT46), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1004), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT114), .Z(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT47), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT47), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n1019), .A3(new_n787), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n950), .A2(new_n800), .A3(new_n951), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n794), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n791), .B1(new_n209), .B2(new_n318), .C1(new_n1022), .C2(new_n241), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n744), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT115), .Z(new_n1025));
  NAND2_X1  g0825(.A1(new_n995), .A2(new_n1025), .ZN(G387));
  AOI22_X1  g0826(.A1(new_n815), .A2(G311), .B1(new_n770), .B2(G303), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n818), .B2(new_n1012), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G322), .B2(new_n751), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(G294), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1031), .B1(new_n759), .B2(new_n748), .C1(new_n1032), .C2(new_n767), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT117), .B(KEYINPUT49), .Z(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1033), .A2(new_n1034), .B1(G326), .B2(new_n833), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n776), .A2(G116), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n823), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n318), .A2(new_n748), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n321), .A2(new_n767), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n263), .B2(new_n760), .C1(new_n773), .C2(new_n779), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1003), .A2(new_n201), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n754), .A2(new_n261), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n770), .A2(G68), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1045), .A2(new_n793), .A3(new_n1010), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1038), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n787), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n679), .A2(new_n681), .A3(new_n800), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n238), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n794), .B1(new_n1051), .B2(new_n283), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n280), .A2(new_n209), .A3(new_n699), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n261), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1052), .A2(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n209), .A2(G107), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n791), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1049), .A2(new_n744), .A3(new_n1050), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n989), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n696), .B1(new_n1061), .B2(new_n740), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1060), .B1(new_n993), .B2(new_n989), .C1(new_n1062), .C2(new_n990), .ZN(G393));
  INV_X1    g0863(.A(new_n979), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n994), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n943), .A2(new_n790), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n751), .B1(new_n764), .B2(G159), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(new_n782), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n815), .A2(G50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n823), .B1(G87), .B2(new_n776), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n769), .A2(new_n261), .B1(new_n760), .B2(new_n819), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G77), .B2(new_n749), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n764), .B1(new_n751), .B2(G317), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G322), .B2(new_n833), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n815), .A2(G303), .B1(new_n749), .B2(G116), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G107), .B2(new_n776), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n329), .B1(new_n767), .B2(new_n759), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1078), .B2(KEYINPUT118), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n769), .A2(new_n1032), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1074), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n787), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n791), .B1(new_n213), .B2(new_n209), .C1(new_n1022), .C2(new_n248), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1066), .A2(new_n744), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1065), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT110), .B1(new_n975), .B2(new_n978), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n990), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n982), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1064), .A2(new_n990), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1089), .B1(new_n1094), .B2(new_n696), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G390));
  NAND4_X1  g0896(.A1(new_n847), .A2(new_n861), .A3(G330), .A4(new_n842), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n861), .B1(new_n810), .B2(new_n923), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n920), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n918), .B2(new_n919), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n736), .A2(new_n724), .A3(new_n806), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n912), .B1(new_n1102), .B2(new_n807), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1100), .B1(new_n917), .B2(new_n887), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1098), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n918), .A2(new_n919), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n914), .B2(new_n920), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n726), .A2(new_n861), .A3(new_n683), .A4(new_n842), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n994), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1107), .A2(new_n788), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n280), .B1(new_n760), .B2(new_n1115), .C1(new_n201), .C2(new_n758), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT120), .Z(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  AOI22_X1  g0918(.A1(new_n815), .A2(G137), .B1(new_n770), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1003), .A2(new_n825), .B1(new_n748), .B2(new_n779), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n782), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n767), .B2(new_n263), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1117), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G128), .B2(new_n751), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G87), .A2(new_n782), .B1(new_n815), .B2(G107), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n213), .B2(new_n769), .C1(new_n1032), .C2(new_n760), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n773), .A2(new_n759), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n758), .A2(new_n203), .B1(new_n748), .B2(new_n539), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n329), .B1(new_n1003), .B2(new_n488), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n787), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n838), .A2(new_n261), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1114), .A2(new_n744), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n847), .A2(G330), .A3(new_n842), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n912), .ZN(new_n1137));
  AND4_X1   g0937(.A1(new_n807), .A2(new_n1137), .A3(new_n1109), .A4(new_n1102), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n912), .B1(new_n727), .B2(new_n808), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n1097), .B1(new_n807), .B2(new_n913), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n896), .A2(new_n897), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n897), .A2(G330), .A3(new_n847), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1145), .A3(new_n655), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n1145), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1142), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(new_n1112), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n696), .B1(new_n1150), .B2(new_n1111), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1113), .B(new_n1135), .C1(new_n1152), .C2(new_n1153), .ZN(G378));
  NAND3_X1  g0954(.A1(new_n924), .A2(new_n921), .A3(new_n901), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT105), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n882), .A2(G330), .A3(new_n890), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1156), .A2(new_n925), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1156), .B2(new_n925), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n302), .B1(new_n402), .B2(new_n399), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n272), .A2(new_n863), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1158), .A2(new_n1159), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1157), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n922), .B2(new_n926), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1156), .A2(new_n925), .A3(new_n1157), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1164), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n994), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n788), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n815), .A2(G132), .B1(new_n749), .B2(G150), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n770), .A2(G137), .B1(G128), .B2(new_n764), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n782), .A2(new_n1118), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G125), .B2(new_n751), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G41), .B1(new_n833), .B2(G124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n274), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G159), .B2(new_n776), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1178), .B2(new_n1177), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1000), .B1(new_n213), .B2(new_n754), .C1(new_n1003), .C2(new_n215), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G116), .B2(new_n751), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n793), .B1(G58), .B2(new_n776), .ZN(new_n1186));
  AND4_X1   g0986(.A1(new_n275), .A2(new_n1185), .A3(new_n1041), .A4(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n759), .B2(new_n760), .C1(new_n318), .C2(new_n769), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G41), .B1(new_n793), .B2(G33), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1183), .B(new_n1190), .C1(G50), .C2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n787), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n838), .A2(new_n201), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1172), .A2(new_n744), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1171), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1148), .B(new_n1149), .C1(new_n1111), .C2(new_n1141), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n697), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(KEYINPUT57), .B(new_n1198), .C1(new_n1166), .C2(new_n1170), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(G375));
  AOI21_X1  g1004(.A(KEYINPUT119), .B1(new_n898), .B2(new_n1145), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n476), .B1(new_n709), .B2(new_n738), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1206), .A2(new_n1144), .A3(new_n1147), .A4(new_n654), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1141), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n966), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1150), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT121), .Z(new_n1211));
  NAND2_X1  g1011(.A1(new_n912), .A2(new_n788), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n818), .A2(new_n817), .B1(new_n825), .B2(new_n773), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n815), .B2(new_n1118), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n833), .A2(G128), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n769), .A2(new_n263), .B1(new_n748), .B2(new_n201), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n823), .A2(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n782), .A2(G159), .B1(new_n776), .B2(G58), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n767), .A2(new_n213), .B1(new_n760), .B2(new_n766), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT122), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1003), .A2(new_n759), .B1(new_n769), .B2(new_n215), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1039), .A2(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n773), .A2(new_n1032), .B1(new_n758), .B2(new_n539), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G116), .B2(new_n815), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1221), .A2(new_n329), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n787), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n838), .A2(new_n203), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1212), .A2(new_n744), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1141), .B2(new_n993), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1211), .A2(new_n1232), .ZN(G381));
  NOR2_X1   g1033(.A1(G375), .A2(G378), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n995), .A2(new_n1025), .A3(new_n1095), .ZN(new_n1235));
  INV_X1    g1035(.A(G381), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(G407));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1234), .B2(new_n676), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G407), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT127), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1197), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1199), .A2(new_n966), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G378), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n696), .A3(new_n1202), .ZN(new_n1248));
  AND4_X1   g1048(.A1(KEYINPUT123), .A2(new_n1248), .A3(G378), .A4(new_n1243), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT123), .B1(new_n1203), .B2(G378), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1246), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1150), .B2(new_n1208), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT60), .B1(new_n1254), .B2(new_n1141), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n1255), .A3(new_n697), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n814), .B(new_n843), .C1(new_n1256), .C2(new_n1231), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1253), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1255), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n696), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(G384), .A3(new_n1232), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1239), .A2(G343), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1251), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT124), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1248), .A2(G378), .A3(new_n1243), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1203), .A2(KEYINPUT123), .A3(G378), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1264), .B1(new_n1273), .B2(new_n1246), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(KEYINPUT124), .A3(new_n1263), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT63), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(G393), .B(G396), .Z(new_n1277));
  AOI21_X1  g1077(.A(new_n1095), .B1(new_n995), .B2(new_n1025), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1235), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(G390), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n995), .A2(new_n1095), .A3(new_n1025), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1277), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1279), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1279), .A2(new_n1283), .A3(KEYINPUT126), .A4(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1263), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1264), .A2(G2897), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT125), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1257), .A2(new_n1261), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1245), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1296), .B2(new_n1264), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1290), .A2(new_n1297), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1276), .A2(new_n1289), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1284), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1274), .B2(new_n1263), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1268), .A2(new_n1275), .A3(new_n1303), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1301), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1242), .B1(new_n1299), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT124), .B1(new_n1274), .B2(new_n1263), .ZN(new_n1309));
  NOR4_X1   g1109(.A1(new_n1296), .A2(new_n1267), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1309), .A2(new_n1310), .A3(KEYINPUT62), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1284), .A3(new_n1297), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1300), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1290), .A2(new_n1297), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(new_n1318), .A3(KEYINPUT127), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1308), .A2(new_n1319), .ZN(G405));
  OAI21_X1  g1120(.A(new_n1273), .B1(G378), .B2(new_n1203), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1300), .B(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1263), .ZN(G402));
endmodule


