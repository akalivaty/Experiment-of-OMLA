//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n191));
  OAI211_X1 g005(.A(G119), .B(new_n190), .C1(new_n191), .C2(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT71), .B1(new_n194), .B2(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(KEYINPUT72), .A3(G110), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT73), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(KEYINPUT73), .A2(G125), .A3(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(KEYINPUT16), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT74), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n216), .A3(G146), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT24), .B(G110), .Z(new_n218));
  XNOR2_X1  g032(.A(G119), .B(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n202), .A2(new_n215), .A3(new_n217), .A4(new_n220), .ZN(new_n221));
  OAI22_X1  g035(.A1(new_n197), .A2(G110), .B1(new_n219), .B2(new_n218), .ZN(new_n222));
  XNOR2_X1  g036(.A(G125), .B(G140), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n213), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n212), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT75), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n221), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n221), .B2(new_n225), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n234), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT25), .B1(new_n234), .B2(new_n188), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n189), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n189), .A2(G902), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT76), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(G472), .A2(G902), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT64), .A2(G143), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(G146), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT65), .B1(new_n247), .B2(G146), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n248), .A2(new_n254), .A3(G146), .A4(new_n249), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n245), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n245), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT64), .A2(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT64), .A2(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n213), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n247), .A2(G146), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT67), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n245), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n259), .A2(new_n260), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n251), .B1(new_n266), .B2(G146), .ZN(new_n267));
  INV_X1    g081(.A(new_n255), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n270));
  INV_X1    g084(.A(new_n263), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT11), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G134), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT66), .B1(new_n276), .B2(G134), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n273), .A3(G137), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n277), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n279), .A4(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n264), .A2(new_n272), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n194), .A2(G116), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G119), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT2), .B(G113), .Z(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n273), .A2(G137), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n276), .A2(G134), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n253), .B2(new_n255), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n261), .A2(new_n262), .B1(G128), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n286), .B(new_n298), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n295), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n226), .A3(G210), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n305), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n288), .A2(KEYINPUT30), .A3(new_n304), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n259), .A2(new_n260), .A3(new_n213), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n255), .B1(new_n314), .B2(new_n251), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n263), .B1(new_n315), .B2(new_n265), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n287), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n304), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n313), .A2(new_n294), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n306), .B1(new_n305), .B2(new_n311), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n244), .B(KEYINPUT31), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n305), .A2(new_n311), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT68), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n312), .A3(new_n321), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n244), .B1(new_n328), .B2(KEYINPUT31), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n318), .A2(new_n294), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n305), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n305), .B2(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT70), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n305), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n311), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n327), .A2(new_n341), .A3(new_n312), .A4(new_n321), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n243), .B1(new_n330), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT31), .B1(new_n322), .B2(new_n323), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n324), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n322), .A2(new_n323), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n341), .A2(new_n350), .B1(new_n338), .B2(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n243), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(new_n345), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n321), .A2(new_n305), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n339), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n355), .B(new_n357), .C1(new_n338), .C2(new_n339), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n288), .A2(new_n304), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n294), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n334), .B1(new_n360), .B2(new_n305), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n305), .A2(new_n334), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n339), .A2(new_n355), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n352), .A2(new_n354), .B1(new_n367), .B2(G472), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n242), .B1(new_n346), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G214), .B1(G237), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  INV_X1    g186(.A(new_n300), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n315), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n303), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n209), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G125), .B1(new_n256), .B2(new_n263), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT82), .B(G224), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G953), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n376), .B2(new_n377), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G122), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  AOI21_X1  g200(.A(G101), .B1(new_n385), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G104), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n386), .A2(new_n387), .A3(new_n390), .A4(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n385), .A2(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n398), .B2(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n396), .A3(G101), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n294), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n389), .A2(G104), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n397), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n393), .A2(new_n394), .B1(G101), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G113), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n290), .A2(G119), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT5), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n292), .A2(new_n293), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(KEYINPUT6), .B(new_n384), .C1(new_n402), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n412), .A3(new_n384), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n412), .A4(new_n384), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n384), .B1(new_n402), .B2(new_n412), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n383), .B(new_n413), .C1(new_n418), .C2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n416), .A2(new_n417), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n384), .B(KEYINPUT8), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n404), .A2(G101), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n395), .A2(new_n411), .A3(KEYINPUT83), .A4(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n405), .B2(new_n411), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT83), .B1(new_n405), .B2(new_n411), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n379), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n376), .A2(new_n377), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT84), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n376), .A2(new_n377), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n430), .B2(new_n379), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n429), .A2(new_n434), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n188), .B1(new_n423), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n372), .B1(new_n422), .B2(new_n439), .ZN(new_n440));
  AND4_X1   g254(.A1(new_n429), .A2(new_n435), .A3(new_n437), .A4(new_n434), .ZN(new_n441));
  AOI21_X1  g255(.A(G902), .B1(new_n441), .B2(new_n418), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n418), .A2(new_n421), .ZN(new_n443));
  INV_X1    g257(.A(new_n383), .ZN(new_n444));
  INV_X1    g258(.A(new_n413), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n446), .A3(KEYINPUT85), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n440), .A2(new_n447), .A3(KEYINPUT86), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n442), .A2(new_n446), .A3(new_n448), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n371), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G469), .ZN(new_n457));
  INV_X1    g271(.A(new_n401), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n395), .B2(new_n399), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n264), .A3(new_n272), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n395), .A2(new_n425), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT64), .B(G143), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n299), .B1(new_n462), .B2(new_n213), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n253), .B(new_n255), .C1(new_n463), .C2(new_n190), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n301), .B1(new_n464), .B2(KEYINPUT78), .ZN(new_n465));
  AOI21_X1  g279(.A(G146), .B1(new_n248), .B2(new_n249), .ZN(new_n466));
  OAI21_X1  g280(.A(G128), .B1(new_n466), .B2(new_n299), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n253), .A4(new_n255), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n461), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n460), .B1(new_n470), .B2(KEYINPUT10), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT10), .B1(new_n301), .B2(new_n303), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(new_n461), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n374), .A2(new_n375), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n405), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n287), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n190), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT78), .B1(new_n315), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n469), .A3(new_n374), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n405), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT10), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n474), .A2(new_n476), .ZN(new_n485));
  INV_X1    g299(.A(new_n287), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n460), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G140), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n226), .A2(G227), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n478), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n484), .A2(new_n485), .A3(new_n460), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n405), .A2(new_n303), .A3(new_n301), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n405), .B2(new_n481), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n496), .B2(new_n486), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n461), .A2(new_n375), .A3(new_n374), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n482), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(KEYINPUT12), .A3(new_n287), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n493), .A2(new_n486), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n492), .B1(new_n501), .B2(new_n491), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n457), .B1(new_n502), .B2(new_n188), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT12), .B1(new_n499), .B2(new_n287), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n494), .B(new_n486), .C1(new_n482), .C2(new_n498), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n487), .A2(new_n491), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n491), .B1(new_n478), .B2(new_n487), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n457), .B(new_n188), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT80), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n264), .A2(new_n272), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n483), .A2(new_n482), .B1(new_n513), .B2(new_n459), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n486), .B1(new_n514), .B2(new_n485), .ZN(new_n515));
  INV_X1    g329(.A(new_n487), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n490), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n497), .A2(new_n500), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n487), .A3(new_n491), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT80), .A3(new_n457), .A4(new_n188), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n503), .B1(new_n512), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT9), .B(G234), .ZN(new_n523));
  OAI21_X1  g337(.A(G221), .B1(new_n523), .B2(G902), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(G128), .A3(new_n266), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n266), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n190), .A2(G143), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(G134), .B(new_n527), .C1(new_n530), .C2(new_n526), .ZN(new_n531));
  INV_X1    g345(.A(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G116), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n290), .A2(G122), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n389), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n533), .A2(new_n534), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT90), .B1(new_n532), .B2(G116), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G107), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n528), .A2(new_n273), .A3(new_n529), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n531), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n535), .B(new_n536), .C1(KEYINPUT14), .C2(new_n389), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT14), .B1(new_n538), .B2(new_n539), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n546), .A3(G107), .ZN(new_n547));
  INV_X1    g361(.A(new_n543), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n273), .B1(new_n528), .B2(new_n529), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n545), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n523), .A2(new_n187), .A3(G953), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n544), .A2(new_n550), .A3(new_n554), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n544), .A2(new_n550), .ZN(new_n556));
  INV_X1    g370(.A(new_n551), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n188), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G952), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  INV_X1    g379(.A(G234), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n307), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n188), .B(new_n226), .C1(G234), .C2(G237), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n559), .B(new_n188), .C1(KEYINPUT15), .C2(new_n561), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n563), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G214), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n575), .A2(G237), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT87), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n266), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n247), .A2(new_n307), .A3(new_n226), .A4(G214), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n266), .B2(KEYINPUT87), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n285), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n307), .A2(new_n226), .A3(G214), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n462), .B2(KEYINPUT87), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n576), .B(new_n247), .C1(new_n246), .C2(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(G131), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT88), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND4_X1   g403(.A1(KEYINPUT17), .A2(new_n584), .A3(G131), .A4(new_n585), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n215), .B2(new_n217), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(KEYINPUT88), .A3(new_n582), .A4(new_n586), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G113), .B(G122), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(new_n385), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n205), .A2(new_n206), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G146), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n224), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n578), .A2(new_n580), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n285), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n598), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n586), .A2(new_n600), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n595), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n595), .B1(new_n593), .B2(new_n605), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n188), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G475), .ZN(new_n610));
  NOR2_X1   g424(.A1(G475), .A2(G902), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n595), .ZN(new_n613));
  MUX2_X1   g427(.A(new_n223), .B(new_n596), .S(KEYINPUT19), .Z(new_n614));
  OAI21_X1  g428(.A(new_n212), .B1(new_n614), .B2(G146), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n586), .B2(new_n581), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n613), .B1(new_n616), .B2(new_n604), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n612), .B1(new_n606), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n606), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT89), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT20), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n620), .A2(new_n621), .A3(new_n618), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n574), .B(new_n610), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n522), .A2(new_n525), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n369), .A2(new_n456), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  NOR3_X1   g441(.A1(new_n522), .A2(new_n242), .A3(new_n525), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n352), .B2(new_n188), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n353), .B1(new_n349), .B2(new_n351), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n449), .B1(new_n422), .B2(new_n439), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n371), .B1(new_n634), .B2(new_n455), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n572), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n610), .B1(new_n623), .B2(new_n622), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n556), .B2(new_n557), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n559), .A2(new_n638), .B1(new_n552), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(G478), .A3(new_n188), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n560), .A2(new_n561), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n633), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT94), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  AND2_X1   g464(.A1(new_n563), .A2(new_n573), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n618), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(KEYINPUT20), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(KEYINPUT20), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT96), .B1(new_n618), .B2(new_n656), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n610), .B(new_n652), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n636), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n633), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NAND2_X1  g481(.A1(new_n221), .A2(new_n225), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT97), .Z(new_n669));
  INV_X1    g483(.A(new_n230), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT36), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n668), .B(KEYINPUT97), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n671), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n675), .A3(new_n239), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n237), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n456), .A2(new_n625), .A3(new_n632), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  OAI21_X1  g494(.A(new_n354), .B1(new_n330), .B2(new_n343), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n367), .A2(G472), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n681), .B(new_n682), .C1(new_n631), .C2(KEYINPUT32), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n512), .A2(new_n521), .ZN(new_n684));
  INV_X1    g498(.A(new_n503), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n525), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n569), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n567), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n663), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n635), .A2(new_n677), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NAND2_X1  g509(.A1(new_n454), .A2(new_n455), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n360), .A2(new_n305), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n339), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT98), .ZN(new_n700));
  AOI21_X1  g514(.A(G902), .B1(new_n700), .B2(new_n328), .ZN(new_n701));
  OAI221_X1 g515(.A(new_n681), .B1(new_n629), .B2(new_n701), .C1(new_n631), .C2(KEYINPUT32), .ZN(new_n702));
  INV_X1    g516(.A(new_n677), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n651), .A2(new_n371), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n637), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT99), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n697), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n690), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n686), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT40), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n266), .ZN(G45));
  NOR2_X1   g528(.A1(new_n644), .A2(new_n691), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n683), .A2(new_n686), .A3(new_n693), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  NAND2_X1  g531(.A1(new_n520), .A2(new_n188), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n525), .B1(new_n718), .B2(G469), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n684), .A2(new_n241), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n683), .A3(new_n645), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT101), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G15));
  NAND3_X1  g538(.A1(new_n720), .A2(new_n664), .A3(new_n683), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND2_X1  g540(.A1(new_n620), .A2(new_n621), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n653), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n620), .A2(new_n621), .A3(new_n618), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n728), .A2(new_n729), .B1(G475), .B2(new_n609), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n574), .A3(new_n677), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n681), .A2(new_n682), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT32), .B1(new_n352), .B2(new_n243), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n684), .A2(new_n719), .A3(new_n635), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n684), .A2(new_n635), .A3(new_n719), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n194), .ZN(G21));
  NAND2_X1  g555(.A1(new_n698), .A2(KEYINPUT28), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n362), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT103), .B1(new_n361), .B2(new_n363), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n744), .A2(new_n745), .A3(new_n339), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n347), .A2(new_n342), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n243), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n630), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n684), .A2(new_n719), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n634), .A2(new_n455), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n704), .A2(new_n637), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n571), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n751), .A3(new_n754), .A4(new_n241), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  INV_X1    g570(.A(new_n715), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n739), .B2(new_n737), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n188), .B1(new_n330), .B2(new_n343), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(G472), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n677), .A4(new_n748), .ZN(new_n762));
  AOI21_X1  g576(.A(G902), .B1(new_n349), .B2(new_n351), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n677), .B(new_n748), .C1(new_n763), .C2(new_n629), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT104), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n455), .A2(new_n370), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n452), .B2(new_n453), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n686), .A2(new_n772), .A3(new_n715), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n683), .A2(new_n241), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n769), .B(new_n770), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n369), .A2(new_n686), .A3(new_n715), .A4(new_n772), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n769), .B1(new_n777), .B2(new_n770), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n773), .A2(new_n774), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT106), .B1(new_n779), .B2(KEYINPUT42), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n773), .A2(new_n774), .A3(new_n781), .A4(new_n770), .ZN(new_n782));
  OAI22_X1  g596(.A1(new_n776), .A2(new_n778), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  NAND4_X1  g598(.A1(new_n369), .A2(new_n686), .A3(new_n692), .A4(new_n772), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  INV_X1    g600(.A(new_n771), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n454), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n730), .A2(new_n643), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT108), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT109), .B1(new_n789), .B2(new_n790), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n730), .A2(new_n796), .A3(KEYINPUT43), .A4(new_n643), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n792), .A2(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n677), .B1(new_n630), .B2(new_n631), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n788), .B1(new_n800), .B2(KEYINPUT44), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(KEYINPUT44), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n457), .B1(new_n502), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT45), .B(new_n492), .C1(new_n501), .C2(new_n491), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n457), .A2(new_n188), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n684), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n809), .A2(new_n810), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n525), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT107), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(new_n710), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n815), .B2(new_n710), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n801), .B(new_n802), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  XNOR2_X1  g634(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n811), .A2(new_n684), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n524), .B1(new_n823), .B2(new_n813), .ZN(new_n824));
  INV_X1    g638(.A(new_n821), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n757), .A2(new_n788), .A3(new_n683), .A4(new_n241), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  NAND2_X1  g644(.A1(new_n792), .A2(new_n794), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n795), .A2(new_n797), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n751), .A2(new_n568), .A3(new_n772), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n369), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT48), .Z(new_n836));
  NOR2_X1   g650(.A1(new_n702), .A2(new_n242), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n750), .A2(new_n241), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n833), .A2(new_n568), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n842));
  INV_X1    g656(.A(new_n737), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI221_X1 g658(.A(new_n565), .B1(new_n838), .B2(new_n644), .C1(new_n841), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n836), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n696), .B(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n371), .A3(new_n751), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n849), .B2(new_n841), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT50), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  OAI211_X1 g666(.A(KEYINPUT116), .B(new_n852), .C1(new_n849), .C2(new_n841), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n833), .A2(new_n766), .A3(new_n834), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n730), .A2(new_n642), .A3(new_n641), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n838), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n718), .A2(G469), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n684), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n822), .B(new_n826), .C1(new_n524), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n841), .A2(new_n788), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n854), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n854), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n846), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(KEYINPUT117), .B(new_n846), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n686), .A2(new_n715), .A3(new_n772), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n766), .A2(KEYINPUT114), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT114), .B1(new_n766), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n563), .A2(new_n573), .A3(new_n690), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n237), .B2(new_n676), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n876), .B(new_n610), .C1(new_n661), .C2(new_n662), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n788), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT113), .B1(new_n687), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n683), .A2(new_n686), .ZN(new_n880));
  INV_X1    g694(.A(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n772), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n785), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n720), .B(new_n683), .C1(new_n664), .C2(new_n645), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n755), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n889), .B2(new_n740), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n731), .B1(new_n346), .B2(new_n368), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n842), .B2(new_n843), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(KEYINPUT111), .A3(new_n755), .A4(new_n888), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n644), .A2(new_n571), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n456), .A2(new_n628), .A3(new_n632), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n896), .A2(new_n626), .A3(KEYINPUT112), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT112), .B1(new_n896), .B2(new_n626), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n730), .A2(new_n652), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n571), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n456), .A2(new_n628), .A3(new_n900), .A4(new_n632), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n678), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n886), .A2(new_n894), .A3(new_n783), .A4(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(KEYINPUT53), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n753), .A2(new_n677), .A3(new_n691), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n702), .A2(new_n906), .A3(new_n686), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n716), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n767), .A3(new_n694), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT52), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(KEYINPUT115), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n767), .A3(KEYINPUT52), .A4(new_n694), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n905), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n912), .A2(new_n914), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT53), .B1(new_n904), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(KEYINPUT54), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n904), .B2(new_n917), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n922));
  OAI221_X1 g736(.A(new_n785), .B1(new_n879), .B2(new_n884), .C1(new_n872), .C2(new_n873), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT105), .B1(new_n779), .B2(KEYINPUT42), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n781), .B1(new_n777), .B2(new_n770), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n779), .A2(KEYINPUT106), .A3(KEYINPUT42), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n775), .A2(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n755), .A4(new_n888), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n929), .A2(new_n897), .A3(new_n898), .A4(new_n902), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n928), .A2(new_n911), .A3(new_n915), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n921), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  OAI22_X1  g747(.A1(new_n870), .A2(new_n933), .B1(G952), .B2(G953), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n859), .B(KEYINPUT49), .Z(new_n935));
  NOR3_X1   g749(.A1(new_n789), .A2(new_n371), .A3(new_n525), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n848), .A2(new_n935), .A3(new_n837), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(G75));
  NAND2_X1  g752(.A1(new_n564), .A2(G953), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT120), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n188), .B1(new_n921), .B2(new_n931), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT56), .B1(new_n941), .B2(G210), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n443), .A2(new_n445), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n383), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n446), .ZN(new_n945));
  XOR2_X1   g759(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n940), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n941), .B2(G210), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(KEYINPUT119), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(KEYINPUT119), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(G51));
  INV_X1    g768(.A(new_n940), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n807), .B(KEYINPUT57), .ZN(new_n956));
  INV_X1    g770(.A(new_n932), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n922), .B1(new_n921), .B2(new_n931), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n520), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n941), .A2(new_n805), .A3(new_n804), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(G54));
  NAND2_X1  g776(.A1(new_n921), .A2(new_n931), .ZN(new_n963));
  AND2_X1   g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(G902), .A3(new_n619), .A4(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT121), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n619), .B1(new_n941), .B2(new_n964), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n955), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n966), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT59), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n640), .B(new_n973), .C1(new_n957), .C2(new_n958), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n940), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n640), .B1(new_n933), .B2(new_n973), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G63));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  XNOR2_X1  g792(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n187), .A2(new_n188), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n921), .B2(new_n931), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n673), .A3(new_n675), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n940), .B1(new_n983), .B2(new_n234), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n983), .A2(new_n234), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n940), .A4(new_n984), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(G66));
  OAI21_X1  g804(.A(G953), .B1(new_n378), .B2(new_n570), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n894), .A2(new_n903), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(G953), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n943), .B1(G898), .B2(new_n226), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT123), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n994), .B(new_n996), .ZN(G69));
  AND3_X1   g811(.A1(new_n819), .A2(new_n785), .A3(new_n829), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n774), .A2(new_n753), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n817), .B2(new_n818), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n767), .A2(new_n694), .A3(new_n716), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n998), .A2(new_n1003), .A3(new_n226), .A4(new_n783), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n313), .A2(new_n320), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(new_n614), .Z(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(G900), .B2(G953), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n226), .B1(G227), .B2(G900), .ZN(new_n1009));
  AOI22_X1  g823(.A1(new_n1004), .A2(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1002), .B(new_n1011), .C1(new_n712), .C2(new_n708), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT62), .B1(new_n713), .B2(new_n1001), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n899), .A2(new_n644), .ZN(new_n1014));
  NOR4_X1   g828(.A1(new_n774), .A2(new_n711), .A3(new_n788), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n827), .B2(new_n828), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n819), .A2(new_n1012), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n226), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n1006), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1010), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1009), .A2(new_n1008), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G72));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1017), .B2(new_n992), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT125), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n339), .B1(new_n321), .B2(new_n305), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n916), .A2(new_n918), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n350), .B1(KEYINPUT127), .B2(new_n357), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(KEYINPUT127), .B2(new_n357), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n1024), .ZN(new_n1033));
  OAI22_X1  g847(.A1(new_n1028), .A2(new_n1029), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n321), .A2(new_n339), .A3(new_n305), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n998), .A2(new_n1003), .A3(new_n783), .A4(new_n993), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n1036), .B2(new_n1024), .ZN(new_n1037));
  OR3_X1    g851(.A1(new_n1037), .A2(KEYINPUT126), .A3(new_n955), .ZN(new_n1038));
  OAI21_X1  g852(.A(KEYINPUT126), .B1(new_n1037), .B2(new_n955), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1034), .B1(new_n1038), .B2(new_n1039), .ZN(G57));
endmodule


