//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT82), .B1(new_n193), .B2(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT69), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT69), .A2(G128), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .A4(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G119), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G119), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n202), .A2(new_n207), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT69), .B(G128), .Z(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n213), .B2(G119), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT24), .B(G110), .Z(new_n215));
  OAI22_X1  g029(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n211), .A2(new_n212), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n194), .B(new_n199), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n207), .A3(new_n210), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n214), .A2(new_n215), .B1(new_n219), .B2(G110), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n197), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n194), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n220), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n218), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT22), .B(G137), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n228), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n218), .B(new_n233), .C1(new_n225), .C2(new_n226), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G217), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(G234), .B2(new_n237), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n235), .A2(G902), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n235), .B2(G902), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n237), .A4(new_n234), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n239), .B1(new_n243), .B2(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G472), .A2(G902), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G119), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n247), .A2(KEYINPUT71), .A3(G119), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT71), .B1(new_n247), .B2(G119), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G113), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT2), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G113), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n257), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G137), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n262), .A2(G134), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI211_X1 g084(.A(KEYINPUT67), .B(KEYINPUT11), .C1(new_n262), .C2(G134), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n265), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n269), .B1(new_n264), .B2(G137), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n268), .A2(new_n267), .A3(new_n269), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n197), .B2(G143), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(KEYINPUT66), .A3(G146), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n282), .B(new_n284), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT0), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n203), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n197), .A2(G143), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n284), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n282), .A2(KEYINPUT64), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT0), .A3(G128), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n289), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n294), .A2(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n197), .A2(G143), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n283), .A2(G146), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n300), .A2(new_n301), .B1(new_n290), .B2(new_n203), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n302), .A3(KEYINPUT65), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n288), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n200), .A2(new_n201), .B1(new_n300), .B2(KEYINPUT1), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n284), .A2(new_n292), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT70), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n301), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(G143), .B2(new_n197), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n308), .B(new_n309), .C1(new_n213), .C2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n283), .A2(KEYINPUT66), .A3(G146), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT66), .B1(new_n283), .B2(G146), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n300), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n307), .A2(new_n312), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  XNOR2_X1  g132(.A(G134), .B(G137), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(new_n279), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n268), .A2(new_n265), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT68), .A3(G131), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n278), .A2(new_n279), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n281), .A2(new_n304), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n261), .B1(new_n324), .B2(KEYINPUT30), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT30), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n281), .A2(new_n304), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n317), .A2(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT30), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT72), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n325), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G237), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G237), .ZN(new_n336));
  AOI21_X1  g150(.A(G953), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G210), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT27), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G101), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n261), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n328), .A2(new_n329), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT74), .B(KEYINPUT31), .C1(new_n332), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n328), .A2(new_n329), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n261), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .A4(new_n342), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n341), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT75), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT75), .B1(new_n351), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n345), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n342), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  AND4_X1   g172(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT30), .A4(new_n329), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n326), .B1(new_n324), .B2(KEYINPUT30), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT31), .ZN(new_n362));
  INV_X1    g176(.A(new_n344), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n362), .B1(new_n361), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(KEYINPUT74), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n246), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT76), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n246), .C1(new_n356), .C2(new_n366), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n350), .B1(new_n324), .B2(new_n342), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT28), .B1(new_n324), .B2(new_n342), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n352), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n353), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n331), .A2(new_n327), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n344), .B1(new_n380), .B2(new_n358), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n381), .B2(new_n362), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n378), .A2(new_n382), .A3(new_n364), .A4(new_n345), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT32), .A3(new_n246), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n324), .A2(new_n342), .ZN(new_n385));
  INV_X1    g199(.A(new_n343), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(KEYINPUT77), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n343), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n346), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n374), .B(KEYINPUT78), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n392));
  NOR4_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n352), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n341), .B1(new_n361), .B2(new_n343), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n351), .B2(new_n352), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n237), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G472), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n384), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n245), .B1(new_n372), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G221), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n237), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G140), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n229), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT3), .B1(new_n408), .B2(G107), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n410));
  INV_X1    g224(.A(G107), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G104), .ZN(new_n412));
  INV_X1    g226(.A(G101), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(G107), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n409), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n408), .A2(G107), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n411), .A2(G104), .ZN(new_n417));
  OAI21_X1  g231(.A(G101), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n307), .A2(new_n312), .A3(new_n316), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n311), .A2(new_n203), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n316), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n281), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(KEYINPUT12), .A3(new_n281), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n419), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n432), .A2(new_n425), .B1(new_n317), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n281), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n409), .A2(new_n412), .A3(new_n414), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(G101), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(G101), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT4), .A3(new_n415), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n304), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n407), .B1(new_n431), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n407), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n435), .B1(new_n434), .B2(new_n441), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT83), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n426), .A2(KEYINPUT12), .A3(new_n281), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT12), .B1(new_n426), .B2(new_n281), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n317), .A2(new_n433), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n425), .A2(new_n432), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n281), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n406), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n281), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n442), .A3(new_n407), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n447), .A2(new_n459), .A3(G469), .ZN(new_n460));
  INV_X1    g274(.A(G469), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n237), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n406), .B1(new_n454), .B2(new_n445), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n442), .B(new_n407), .C1(new_n448), .C2(new_n449), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n465), .B2(new_n461), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n403), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G214), .B1(G237), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(G224), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n421), .A2(KEYINPUT0), .A3(G128), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n293), .A2(new_n289), .A3(new_n297), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT65), .B1(new_n299), .B2(new_n302), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n307), .A2(new_n312), .A3(new_n191), .A4(new_n316), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT86), .B1(new_n475), .B2(G125), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n304), .B2(new_n191), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT86), .ZN(new_n482));
  INV_X1    g296(.A(new_n479), .ZN(new_n483));
  INV_X1    g297(.A(new_n470), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n249), .B(KEYINPUT5), .C1(new_n250), .C2(new_n251), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT5), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n253), .B1(new_n248), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n489), .B1(new_n488), .B2(new_n491), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n260), .A2(new_n415), .A3(new_n418), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n261), .A2(new_n438), .A3(new_n440), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n487), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(new_n491), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT84), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n499), .A2(new_n260), .A3(new_n424), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n261), .A2(new_n438), .A3(new_n440), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G122), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n497), .A2(new_n510), .A3(new_n503), .A4(new_n505), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n486), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n484), .A2(KEYINPUT7), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n478), .B2(new_n479), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n482), .A2(new_n483), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n504), .B(KEYINPUT8), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n492), .A2(new_n493), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n424), .B1(new_n518), .B2(new_n260), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n494), .B1(new_n488), .B2(new_n491), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n514), .A2(new_n507), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n237), .ZN(new_n523));
  OAI21_X1  g337(.A(G210), .B1(G237), .B2(G902), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n512), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n478), .A2(new_n479), .A3(new_n513), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n515), .B1(new_n482), .B2(new_n483), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n521), .A2(new_n507), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n486), .A2(new_n509), .A3(new_n511), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n524), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n468), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G952), .ZN(new_n535));
  AOI211_X1 g349(.A(G953), .B(new_n535), .C1(G234), .C2(G237), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n237), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n283), .A2(G128), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n540), .B(KEYINPUT13), .Z(new_n541));
  NAND3_X1  g355(.A1(new_n200), .A2(G143), .A3(new_n201), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G134), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G122), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G116), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n247), .A2(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(G107), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(new_n264), .A3(new_n540), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n542), .A2(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G134), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n546), .A2(KEYINPUT14), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G107), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n548), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n555), .A2(G107), .A3(new_n546), .A4(new_n547), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(KEYINPUT90), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT90), .B1(new_n554), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n551), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n401), .A2(new_n236), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n551), .B(new_n564), .C1(new_n561), .C2(new_n562), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n237), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n572), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n569), .A3(new_n237), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n335), .A2(G237), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n578));
  OAI211_X1 g392(.A(G214), .B(new_n229), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n283), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n337), .A2(G143), .A3(G214), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n279), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n224), .B1(new_n582), .B2(KEYINPUT17), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n283), .ZN(new_n584));
  AOI21_X1  g398(.A(G143), .B1(new_n337), .B2(G214), .ZN(new_n585));
  OAI21_X1  g399(.A(G131), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n580), .A2(new_n279), .A3(new_n581), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G113), .B(G122), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n408), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT18), .B(G131), .C1(new_n584), .C2(new_n585), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n193), .A2(KEYINPUT87), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT87), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n190), .A2(new_n192), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(G146), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n199), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(KEYINPUT18), .A2(G131), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n580), .A2(new_n581), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n593), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n590), .A2(new_n592), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n598), .A2(new_n600), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n589), .A2(new_n583), .B1(new_n604), .B2(new_n593), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT89), .B1(new_n605), .B2(new_n592), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n590), .A2(new_n601), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n608));
  INV_X1    g422(.A(new_n592), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n603), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G475), .B1(new_n611), .B2(G902), .ZN(new_n612));
  NOR2_X1   g426(.A1(G475), .A2(G902), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n594), .A2(KEYINPUT19), .A3(new_n596), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n193), .A2(KEYINPUT19), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n197), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n588), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n194), .B(new_n617), .C1(new_n618), .C2(new_n582), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n592), .B1(new_n619), .B2(new_n601), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(KEYINPUT88), .B1(new_n605), .B2(new_n592), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT88), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n586), .A2(new_n588), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n617), .A2(new_n194), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n623), .A2(new_n624), .B1(new_n604), .B2(new_n593), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n622), .B1(new_n625), .B2(new_n592), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT20), .B(new_n614), .C1(new_n621), .C2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n619), .A2(new_n601), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT88), .A3(new_n609), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n602), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n631), .B2(new_n613), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n612), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NOR4_X1   g447(.A1(new_n534), .A2(new_n539), .A3(new_n576), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n399), .A2(new_n467), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n460), .A2(new_n466), .ZN(new_n637));
  INV_X1    g451(.A(new_n403), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n637), .A2(new_n244), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n237), .B1(new_n356), .B2(new_n366), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n639), .A2(new_n368), .A3(new_n641), .A4(new_n371), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT92), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n371), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n370), .B1(new_n383), .B2(new_n246), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n647), .A2(KEYINPUT92), .A3(new_n641), .A4(new_n639), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n468), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT93), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n526), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n525), .B1(new_n512), .B2(new_n523), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n531), .A2(new_n532), .A3(new_n524), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(KEYINPUT93), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT94), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n567), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n568), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n566), .B(new_n567), .C1(new_n658), .C2(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n571), .A2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT95), .B(G478), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n568), .B2(new_n237), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n539), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n633), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n656), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n649), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  NAND2_X1  g489(.A1(new_n630), .A2(new_n602), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n620), .A2(KEYINPUT88), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n613), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT20), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n631), .A2(new_n628), .A3(new_n613), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n576), .A3(new_n612), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n656), .A2(new_n539), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n649), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT35), .B(G107), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  INV_X1    g500(.A(new_n238), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n241), .B2(new_n242), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n227), .B1(KEYINPUT36), .B2(new_n231), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n218), .B(new_n691), .C1(new_n225), .C2(new_n226), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n237), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT96), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n467), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n634), .A2(new_n647), .A3(new_n641), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  AOI21_X1  g515(.A(new_n697), .B1(new_n372), .B2(new_n398), .ZN(new_n702));
  INV_X1    g516(.A(new_n656), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT97), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n537), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n536), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n704), .B1(new_n682), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n611), .A2(G902), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n711), .A2(G475), .B1(new_n679), .B2(new_n680), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(KEYINPUT97), .A3(new_n576), .A4(new_n708), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n702), .A2(new_n703), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XNOR2_X1  g531(.A(new_n708), .B(KEYINPUT39), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n467), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(KEYINPUT40), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n526), .A2(new_n533), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT38), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT38), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n633), .A2(new_n576), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n693), .B(KEYINPUT96), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n688), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n468), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n720), .A2(new_n724), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n341), .B1(new_n387), .B2(new_n389), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n237), .B1(new_n730), .B2(new_n381), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G472), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n372), .A2(new_n384), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n719), .A2(KEYINPUT40), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  AOI21_X1  g550(.A(new_n667), .B1(new_n662), .B2(new_n663), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n681), .B2(new_n612), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT98), .B1(new_n738), .B2(new_n708), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n633), .A2(new_n669), .A3(KEYINPUT98), .A4(new_n708), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n702), .A2(new_n703), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G146), .ZN(G48));
  NAND2_X1  g558(.A1(new_n372), .A2(new_n398), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n463), .A2(new_n464), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n237), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n465), .A2(new_n461), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n748), .A2(new_n749), .A3(new_n638), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n745), .A2(new_n672), .A3(new_n244), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT41), .B(G113), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G15));
  NAND4_X1  g567(.A1(new_n745), .A2(new_n683), .A3(new_n244), .A4(new_n750), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G116), .ZN(G18));
  NAND3_X1  g569(.A1(new_n652), .A2(new_n655), .A3(new_n750), .ZN(new_n756));
  INV_X1    g570(.A(new_n576), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n696), .A2(new_n712), .A3(new_n670), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n745), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  INV_X1    g575(.A(G472), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n383), .B2(new_n237), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n748), .A2(new_n749), .A3(new_n638), .A4(new_n670), .ZN(new_n764));
  INV_X1    g578(.A(new_n246), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n332), .A2(KEYINPUT31), .A3(new_n344), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n365), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n352), .B1(new_n390), .B2(new_n391), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n763), .A2(new_n245), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n656), .A2(new_n725), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G122), .ZN(G24));
  INV_X1    g587(.A(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n633), .A2(new_n669), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(new_n709), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n769), .B1(new_n640), .B2(G472), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n696), .A3(new_n777), .A4(new_n740), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT99), .B1(new_n778), .B2(new_n756), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n763), .A2(new_n727), .A3(new_n769), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT99), .ZN(new_n781));
  INV_X1    g595(.A(new_n756), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n742), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  NAND2_X1  g599(.A1(new_n367), .A2(new_n369), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n384), .A3(new_n397), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n244), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT101), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT101), .A3(new_n244), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n776), .A2(new_n740), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n653), .A2(new_n468), .A3(new_n654), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT100), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n653), .A2(new_n654), .A3(new_n797), .A4(new_n468), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n443), .A2(new_n446), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(G469), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n403), .B1(new_n466), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n796), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n793), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n802), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n745), .A2(new_n742), .A3(new_n804), .A4(new_n244), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n792), .A2(new_n803), .B1(new_n805), .B2(new_n794), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n279), .ZN(G33));
  INV_X1    g621(.A(KEYINPUT102), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n714), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n710), .A2(KEYINPUT102), .A3(new_n713), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n399), .A2(new_n809), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G134), .ZN(G36));
  NAND2_X1  g626(.A1(new_n447), .A2(new_n459), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n461), .B1(new_n799), .B2(KEYINPUT45), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n462), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n749), .B1(new_n817), .B2(KEYINPUT46), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n638), .B(new_n718), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT103), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n796), .A2(new_n798), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n712), .A2(new_n669), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT43), .B1(new_n824), .B2(KEYINPUT104), .ZN(new_n825));
  OAI211_X1 g639(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n633), .C2(new_n737), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n647), .A2(new_n641), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n696), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT44), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(KEYINPUT44), .A3(new_n829), .A4(new_n696), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n821), .A2(new_n823), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G137), .ZN(G39));
  OAI21_X1  g649(.A(new_n638), .B1(new_n818), .B2(new_n819), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT47), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n745), .A2(new_n793), .A3(new_n244), .A4(new_n822), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  NOR2_X1   g657(.A1(G952), .A2(G953), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT117), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n750), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n707), .B1(new_n846), .B2(KEYINPUT113), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n828), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n763), .A2(new_n245), .A3(new_n707), .A4(new_n769), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n828), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n750), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n468), .B(new_n854), .C1(new_n723), .C2(new_n722), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n853), .A2(KEYINPUT50), .A3(new_n855), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n780), .A2(new_n850), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n852), .A2(KEYINPUT112), .A3(new_n822), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT112), .B1(new_n852), .B2(new_n822), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n748), .A2(new_n749), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n638), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n861), .B(new_n862), .C1(new_n840), .C2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n733), .A2(new_n245), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n712), .A2(new_n737), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n847), .A2(new_n848), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n867), .A2(KEYINPUT115), .A3(new_n875), .A4(KEYINPUT51), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n860), .A2(new_n866), .A3(new_n874), .A4(new_n873), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n792), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n882));
  OR3_X1    g696(.A1(new_n849), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n847), .A2(new_n848), .A3(new_n738), .A4(new_n868), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n849), .B2(new_n881), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n535), .B(G953), .C1(new_n853), .C2(new_n782), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n876), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n702), .B(new_n703), .C1(new_n715), .C2(new_n742), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n727), .A2(new_n708), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT109), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n733), .A3(new_n771), .A4(new_n801), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n784), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n784), .A2(new_n890), .A3(new_n897), .A4(new_n893), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n745), .A2(new_n759), .B1(new_n770), .B2(new_n771), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n754), .A3(new_n751), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n805), .A2(new_n794), .ZN(new_n902));
  INV_X1    g716(.A(new_n791), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT101), .B1(new_n787), .B2(new_n244), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n803), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT108), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n778), .B2(new_n802), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n742), .A2(new_n804), .A3(new_n780), .A4(KEYINPUT108), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n633), .A2(new_n576), .A3(new_n709), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n702), .A2(new_n823), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n910), .A2(new_n811), .A3(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT106), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n671), .B2(new_n534), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n738), .A2(new_n918), .A3(KEYINPUT106), .A4(new_n670), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n644), .A2(new_n920), .A3(new_n648), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n635), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT107), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n635), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n534), .A2(new_n682), .A3(new_n539), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n644), .A2(new_n648), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n699), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n923), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n899), .A2(new_n914), .A3(new_n915), .A4(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(KEYINPUT107), .B2(new_n922), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n906), .A2(new_n933), .A3(new_n925), .A4(new_n913), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n894), .A2(KEYINPUT52), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n898), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT53), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n937), .A3(KEYINPUT54), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT111), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n806), .A2(new_n939), .A3(new_n901), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n905), .A2(new_n902), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n900), .A2(new_n754), .A3(new_n751), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT111), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n910), .A2(KEYINPUT53), .A3(new_n811), .A4(new_n912), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n930), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n899), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n915), .B1(new_n934), .B2(new_n936), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT54), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n938), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n845), .B1(new_n889), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n244), .A2(new_n638), .A3(new_n468), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n953), .B(new_n824), .C1(KEYINPUT49), .C2(new_n864), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT105), .Z(new_n955));
  OAI21_X1  g769(.A(new_n724), .B1(KEYINPUT49), .B2(new_n864), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(new_n733), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n955), .B2(new_n957), .ZN(G75));
  NAND2_X1  g772(.A1(new_n947), .A2(new_n948), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(G210), .A3(G902), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n509), .A2(new_n511), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n486), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT55), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n960), .B2(new_n961), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n229), .A2(G952), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(G51));
  XNOR2_X1  g782(.A(new_n462), .B(KEYINPUT57), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n746), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n237), .B1(new_n947), .B2(new_n948), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n815), .A3(new_n816), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n967), .B1(new_n973), .B2(new_n975), .ZN(G54));
  INV_X1    g790(.A(new_n967), .ZN(new_n977));
  NAND2_X1  g791(.A1(KEYINPUT58), .A2(G475), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n237), .B(new_n978), .C1(new_n947), .C2(new_n948), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n979), .B2(new_n631), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n974), .A2(KEYINPUT58), .A3(G475), .A4(new_n631), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT118), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT118), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n983), .A3(new_n631), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(G60));
  NAND2_X1  g799(.A1(G478), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT59), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n662), .B1(new_n951), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n662), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n959), .A2(KEYINPUT54), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n950), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n989), .A2(new_n992), .A3(new_n967), .ZN(G63));
  XNOR2_X1  g807(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(G217), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT119), .Z(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT60), .Z(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n947), .B2(new_n948), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n235), .B(KEYINPUT120), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n977), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n690), .A2(new_n692), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n959), .A2(new_n1004), .A3(new_n998), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n995), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n959), .A2(new_n998), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1001), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1008), .A2(new_n977), .A3(new_n1009), .A4(new_n994), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1006), .A2(new_n1010), .ZN(G66));
  NOR2_X1   g825(.A1(new_n930), .A2(new_n901), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(G953), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT122), .ZN(new_n1014));
  OAI21_X1  g828(.A(G953), .B1(new_n538), .B2(new_n469), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n962), .B1(G898), .B2(new_n229), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1017), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1014), .A2(new_n1019), .A3(new_n1015), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1018), .A2(new_n1020), .ZN(G69));
  AND2_X1   g835(.A1(new_n784), .A2(new_n890), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n821), .A2(new_n771), .A3(new_n792), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n834), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n842), .A2(new_n941), .A3(new_n811), .ZN(new_n1025));
  OR3_X1    g839(.A1(new_n1024), .A2(G953), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n380), .B1(KEYINPUT30), .B2(new_n324), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n615), .A2(new_n616), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1026), .B(new_n1029), .C1(new_n705), .C2(new_n229), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n719), .B1(new_n775), .B2(new_n682), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n399), .A2(new_n823), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n834), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(KEYINPUT124), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT124), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n834), .A2(new_n1035), .A3(new_n1032), .ZN(new_n1036));
  AOI22_X1  g850(.A1(new_n1034), .A2(new_n1036), .B1(new_n840), .B2(new_n841), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1022), .A2(new_n735), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(G953), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1029), .B(KEYINPUT123), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1030), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n229), .B1(G227), .B2(G900), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1044), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1030), .B(new_n1046), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(G72));
  NAND2_X1  g862(.A1(new_n361), .A2(new_n343), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1049), .B(KEYINPUT126), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1050), .A2(new_n341), .ZN(new_n1051));
  NOR4_X1   g865(.A1(new_n1024), .A2(new_n1025), .A3(new_n930), .A4(new_n901), .ZN(new_n1052));
  NAND2_X1  g866(.A1(G472), .A2(G902), .ZN(new_n1053));
  XOR2_X1   g867(.A(new_n1053), .B(KEYINPUT63), .Z(new_n1054));
  INV_X1    g868(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1051), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1054), .B1(new_n394), .B2(new_n381), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1057), .B(KEYINPUT127), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n932), .A2(new_n937), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1056), .A2(new_n977), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1050), .A2(new_n341), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1062));
  NAND4_X1  g876(.A1(new_n1062), .A2(new_n842), .A3(new_n1040), .A4(new_n1012), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1063), .A2(new_n1054), .ZN(new_n1064));
  INV_X1    g878(.A(KEYINPUT125), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1063), .A2(KEYINPUT125), .A3(new_n1054), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1060), .B1(new_n1066), .B2(new_n1067), .ZN(G57));
endmodule


