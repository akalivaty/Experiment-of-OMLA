//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n465), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(new_n464), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n483));
  OAI211_X1 g058(.A(G138), .B(new_n466), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n470), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n470), .A2(KEYINPUT68), .A3(new_n487), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n476), .B2(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(KEYINPUT69), .A3(G651), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n501), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n499), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n509), .A2(new_n499), .A3(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n517), .A2(new_n518), .B1(G651), .B2(new_n524), .ZN(G166));
  NAND2_X1  g100(.A1(new_n508), .A2(G51), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n514), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n511), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n508), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n514), .A2(G90), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n503), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  AOI22_X1  g115(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT71), .B1(new_n541), .B2(new_n503), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n522), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(new_n546), .A3(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT72), .B(G43), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n506), .A2(G543), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n506), .A2(G81), .A3(new_n511), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND4_X1  g135(.A1(new_n510), .A2(G53), .A3(G543), .A4(new_n512), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT73), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n506), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n506), .A2(new_n567), .A3(new_n511), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(G91), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n561), .A2(KEYINPUT73), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n503), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n565), .A2(new_n569), .A3(new_n571), .A4(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n524), .A2(G651), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n509), .A2(new_n499), .A3(new_n515), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n516), .ZN(G303));
  AND4_X1   g153(.A1(new_n567), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n567), .B1(new_n506), .B2(new_n511), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G87), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n511), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n508), .A2(G49), .B1(G651), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n522), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n507), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n566), .A2(G86), .A3(new_n568), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(G47), .A2(new_n508), .B1(new_n514), .B2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n522), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n503), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(new_n599), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n596), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT76), .B(G66), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n511), .A2(new_n606), .B1(G79), .B2(G543), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n507), .A2(new_n605), .B1(new_n607), .B2(new_n503), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n566), .A2(G92), .A3(new_n568), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .A4(new_n568), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G868), .ZN(G284));
  XOR2_X1   g189(.A(G284), .B(KEYINPUT77), .Z(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT78), .ZN(new_n617));
  AND4_X1   g192(.A1(new_n565), .A2(new_n569), .A3(new_n571), .A4(new_n574), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(G868), .B2(new_n618), .ZN(G280));
  XOR2_X1   g194(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n613), .B1(new_n621), .B2(G860), .ZN(G148));
  NOR2_X1   g197(.A1(new_n553), .A2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n613), .A2(new_n621), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(new_n625));
  AOI21_X1  g200(.A(new_n623), .B1(new_n625), .B2(G868), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n470), .A2(new_n467), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G111), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n632), .A2(KEYINPUT81), .B1(new_n633), .B2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(KEYINPUT81), .B2(new_n632), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n476), .A2(G123), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n465), .A2(G135), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n631), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G14), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  AOI21_X1  g241(.A(KEYINPUT18), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n674), .B2(new_n680), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT84), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(KEYINPUT84), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n683), .A2(KEYINPUT84), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n689), .A3(new_n685), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT85), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(new_n693), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n687), .A2(new_n696), .A3(new_n690), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(new_n694), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(G160), .A2(G29), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  AND2_X1   g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT92), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G2084), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT94), .ZN(new_n711));
  NOR2_X1   g286(.A1(G29), .A2(G35), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G162), .B2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2090), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n703), .A2(G33), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n465), .A2(KEYINPUT89), .A3(G139), .ZN(new_n724));
  AOI21_X1  g299(.A(KEYINPUT89), .B1(new_n465), .B2(G139), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n722), .B1(new_n466), .B2(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n719), .B1(new_n728), .B2(new_n703), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT91), .B(G2072), .Z(new_n730));
  XOR2_X1   g305(.A(new_n729), .B(new_n730), .Z(new_n731));
  AOI211_X1 g306(.A(new_n718), .B(new_n731), .C1(new_n716), .C2(new_n715), .ZN(new_n732));
  NOR2_X1   g307(.A1(G4), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n613), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT87), .B(G1348), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G16), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n554), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(G19), .ZN(new_n740));
  INV_X1    g315(.A(G1341), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G11), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(G28), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n703), .B1(new_n744), .B2(G28), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n743), .B1(new_n745), .B2(new_n746), .C1(new_n638), .C2(new_n703), .ZN(new_n747));
  INV_X1    g322(.A(new_n708), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G2084), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n703), .A2(G32), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n753), .A2(new_n754), .B1(G105), .B2(new_n467), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n465), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n476), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n750), .B1(new_n759), .B2(new_n703), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(G164), .A2(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G27), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n742), .A2(new_n749), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n703), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT88), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n465), .A2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n476), .A2(G128), .ZN(new_n773));
  OR2_X1    g348(.A1(G104), .A2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(G29), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2067), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n738), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n738), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  NOR2_X1   g356(.A1(G5), .A2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT93), .Z(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G301), .B2(new_n738), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n768), .A2(new_n778), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n740), .A2(new_n741), .B1(G1966), .B2(new_n780), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n784), .A2(new_n785), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n767), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n738), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n618), .B2(new_n738), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n737), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G6), .B(G305), .S(G16), .Z(new_n800));
  XOR2_X1   g375(.A(KEYINPUT32), .B(G1981), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n738), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n738), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(G1971), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G1971), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n738), .A2(G23), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n585), .B2(new_n738), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT33), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1976), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G24), .B(G290), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT86), .B(G1986), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n476), .A2(G119), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n465), .A2(G131), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n466), .A2(G107), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(G29), .Z(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n813), .A2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT36), .B1(new_n832), .B2(new_n815), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n799), .B1(new_n831), .B2(new_n833), .ZN(G311));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n798), .ZN(G150));
  NAND2_X1  g411(.A1(new_n613), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  INV_X1    g414(.A(G80), .ZN(new_n840));
  INV_X1    g415(.A(G543), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n522), .A2(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT97), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n844));
  OAI221_X1 g419(.A(new_n844), .B1(new_n840), .B2(new_n841), .C1(new_n522), .C2(new_n839), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(G651), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n506), .A2(G55), .A3(G543), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n506), .A2(G93), .A3(new_n511), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n553), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n548), .A2(new_n846), .A3(new_n552), .A4(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n838), .B(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n856), .A2(new_n857), .A3(G860), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n850), .A2(G860), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(G160), .B(KEYINPUT98), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n465), .A2(G142), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n476), .A2(G130), .ZN(new_n865));
  OR2_X1    g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n497), .B(new_n776), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n759), .ZN(new_n870));
  NOR2_X1   g445(.A1(G164), .A2(new_n776), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n492), .A2(new_n496), .A3(new_n776), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n758), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n873), .A3(new_n726), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n727), .B1(new_n870), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n629), .B(new_n825), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n873), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n728), .ZN(new_n880));
  INV_X1    g455(.A(new_n868), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n874), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n878), .B1(new_n877), .B2(new_n882), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n863), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n638), .B(new_n480), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n877), .A2(new_n882), .ZN(new_n889));
  INV_X1    g464(.A(new_n878), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n891), .A2(new_n884), .A3(new_n883), .A4(new_n862), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n888), .B1(new_n887), .B2(new_n892), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n895), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(G395));
  INV_X1    g477(.A(G868), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT102), .B1(new_n850), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G166), .A2(G288), .ZN(new_n905));
  NAND2_X1  g480(.A1(G303), .A2(new_n585), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G305), .B(G290), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n908), .A3(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n912), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n611), .A2(new_n612), .ZN(new_n916));
  INV_X1    g491(.A(new_n608), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(G299), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n573), .B1(new_n581), .B2(G91), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(KEYINPUT100), .A3(new_n565), .A4(new_n571), .ZN(new_n922));
  NAND2_X1  g497(.A1(G299), .A2(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n613), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n625), .A2(new_n854), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n625), .A2(new_n854), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n625), .A2(new_n854), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n625), .A2(new_n854), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT41), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n922), .A2(new_n613), .A3(new_n923), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n613), .A2(new_n618), .A3(KEYINPUT100), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n915), .A2(new_n929), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G868), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n915), .B1(new_n937), .B2(new_n929), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n904), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n915), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n929), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(KEYINPUT102), .A3(G868), .A4(new_n938), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(G295));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n941), .A2(new_n947), .A3(new_n945), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n941), .B2(new_n945), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n951));
  INV_X1    g526(.A(new_n852), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n548), .A2(new_n552), .B1(new_n846), .B2(new_n849), .ZN(new_n953));
  OAI21_X1  g528(.A(G171), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n851), .A2(G301), .A3(new_n852), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G168), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n851), .A2(G301), .A3(new_n852), .ZN(new_n957));
  AOI21_X1  g532(.A(G301), .B1(new_n851), .B2(new_n852), .ZN(new_n958));
  OAI21_X1  g533(.A(G286), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n936), .A2(new_n932), .A3(new_n956), .A4(new_n959), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n957), .A2(new_n958), .A3(G286), .ZN(new_n961));
  AOI21_X1  g536(.A(G168), .B1(new_n954), .B2(new_n955), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n926), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n912), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(KEYINPUT104), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n961), .A2(new_n962), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n932), .A4(new_n936), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n963), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n912), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT105), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n966), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n951), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n976), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n971), .B2(new_n972), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n965), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n965), .B1(new_n912), .B2(new_n964), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n979), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n991), .ZN(G397));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n492), .B2(new_n496), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n469), .A2(new_n473), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n582), .A2(G1976), .A3(new_n584), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT52), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n585), .B2(G1976), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n593), .A2(new_n1004), .A3(new_n594), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n514), .A2(G86), .ZN(new_n1006));
  OAI21_X1  g581(.A(G1981), .B1(new_n1006), .B2(new_n592), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(new_n1007), .A3(KEYINPUT49), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n997), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT110), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1010), .A2(new_n1014), .A3(new_n1011), .A4(new_n997), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1003), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n497), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT109), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n471), .A2(new_n472), .ZN(new_n1027));
  OAI211_X1 g602(.A(G40), .B(new_n468), .C1(new_n1027), .C2(new_n466), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1971), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n996), .B1(new_n994), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1030), .A2(new_n1031), .B1(new_n1035), .B2(new_n716), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1020), .B1(new_n1036), .B2(new_n993), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1019), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1017), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n716), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(G8), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1016), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1030), .B2(G2078), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT111), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1028), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1045), .A2(G2078), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n994), .A2(new_n1050), .A3(KEYINPUT45), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT119), .B(G1961), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(G171), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(G171), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT120), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1044), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1061));
  INV_X1    g636(.A(G1966), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1061), .A2(new_n1062), .B1(new_n1035), .B2(new_n709), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n993), .B1(new_n1063), .B2(G168), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1035), .A2(new_n709), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G286), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT51), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  AOI211_X1 g646(.A(KEYINPUT51), .B(new_n993), .C1(new_n1063), .C2(G168), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT62), .B1(new_n1076), .B2(new_n1072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1060), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1036), .A2(new_n993), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1016), .A2(new_n1039), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1005), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G288), .A2(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n997), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1080), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1067), .A2(G8), .A3(G168), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1044), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1079), .B1(new_n1090), .B2(new_n1039), .ZN(new_n1091));
  NOR4_X1   g666(.A1(new_n1063), .A2(new_n1087), .A3(new_n993), .A4(G286), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1020), .B(KEYINPUT112), .C1(new_n1036), .C2(new_n993), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1016), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1086), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1078), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n618), .B(KEYINPUT57), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n795), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .A4(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n994), .A2(new_n996), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G2067), .ZN(new_n1104));
  XOR2_X1   g679(.A(new_n1104), .B(KEYINPUT113), .Z(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(G1348), .B2(new_n1035), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n613), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(new_n1098), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G299), .B(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT114), .B(G1996), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .A4(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(new_n741), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1103), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1118), .B2(new_n554), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1112), .A3(new_n554), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT59), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  AOI211_X1 g701(.A(KEYINPUT116), .B(new_n553), .C1(new_n1114), .C2(new_n1117), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1110), .A2(new_n1101), .A3(KEYINPUT61), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1122), .A2(new_n1125), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT117), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1129), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT61), .B1(new_n1110), .B2(new_n1101), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1128), .A4(new_n1122), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1106), .A2(KEYINPUT60), .A3(new_n918), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1106), .B(new_n613), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(KEYINPUT60), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1111), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n765), .A2(KEYINPUT122), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1049), .B2(KEYINPUT122), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1048), .A2(KEYINPUT121), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT121), .B(new_n996), .C1(new_n994), .C2(KEYINPUT45), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1142), .A2(new_n1143), .A3(G301), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT123), .B1(new_n1152), .B2(G171), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1059), .A2(new_n1151), .A3(new_n1153), .A4(new_n1057), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1044), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1157));
  AOI21_X1  g732(.A(G301), .B1(new_n1152), .B2(KEYINPUT124), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(KEYINPUT124), .B2(new_n1152), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1055), .A2(G171), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1159), .A2(KEYINPUT125), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT125), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1156), .B(new_n1157), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1096), .B1(new_n1141), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n776), .B(G2067), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT107), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n825), .B(new_n828), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT108), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n758), .B(G1996), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(G290), .B(G1986), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n994), .A2(KEYINPUT45), .A3(new_n1028), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1176), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1179), .A2(G1986), .A3(G290), .ZN(new_n1181));
  XOR2_X1   g756(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1182));
  XNOR2_X1  g757(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1176), .B1(new_n1169), .B2(new_n758), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT46), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1179), .B2(G1996), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n1179), .A2(new_n1186), .A3(G1996), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT47), .Z(new_n1190));
  OR4_X1    g765(.A1(new_n828), .A2(new_n1169), .A3(new_n825), .A4(new_n1172), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(G2067), .B2(new_n776), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n1184), .B(new_n1190), .C1(new_n1176), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1178), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g769(.A1(new_n896), .A2(new_n898), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n1197));
  NOR2_X1   g771(.A1(G227), .A2(new_n459), .ZN(new_n1198));
  INV_X1    g772(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1197), .B1(G401), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g774(.A(new_n660), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1201), .A2(new_n658), .ZN(new_n1202));
  OAI211_X1 g776(.A(KEYINPUT127), .B(new_n1198), .C1(new_n1202), .C2(new_n655), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n1200), .A2(new_n700), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g778(.A1(new_n1196), .A2(new_n990), .A3(new_n1204), .ZN(G308));
  NAND3_X1  g779(.A1(new_n1196), .A2(new_n990), .A3(new_n1204), .ZN(G225));
endmodule


