

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n621), .A2(n688), .ZN(n670) );
  NOR2_X1 U552 ( .A1(n670), .A2(n1018), .ZN(n622) );
  XNOR2_X1 U553 ( .A(n627), .B(n670), .ZN(n650) );
  INV_X1 U554 ( .A(G2104), .ZN(n546) );
  XOR2_X1 U555 ( .A(KEYINPUT1), .B(n535), .Z(n800) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n687) );
  AND2_X1 U557 ( .A1(n544), .A2(n519), .ZN(G160) );
  NAND2_X1 U558 ( .A1(n527), .A2(n526), .ZN(n525) );
  INV_X1 U559 ( .A(n649), .ZN(n526) );
  XNOR2_X1 U560 ( .A(n648), .B(KEYINPUT29), .ZN(n649) );
  NAND2_X1 U561 ( .A1(n546), .A2(n531), .ZN(n530) );
  INV_X1 U562 ( .A(G2105), .ZN(n531) );
  NOR2_X1 U563 ( .A1(n650), .A2(n1012), .ZN(n637) );
  AND2_X1 U564 ( .A1(n525), .A2(n517), .ZN(n524) );
  XNOR2_X1 U565 ( .A(n687), .B(KEYINPUT89), .ZN(n621) );
  NOR2_X1 U566 ( .A1(G651), .A2(n588), .ZN(n804) );
  AND2_X1 U567 ( .A1(n545), .A2(n518), .ZN(n519) );
  XNOR2_X1 U568 ( .A(n647), .B(KEYINPUT28), .ZN(n516) );
  OR2_X1 U569 ( .A1(G301), .A2(n657), .ZN(n517) );
  AND2_X1 U570 ( .A1(n548), .A2(n547), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n662) );
  NOR2_X1 U572 ( .A1(n528), .A2(n649), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n524), .A2(n522), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n528), .A2(n523), .ZN(n522) );
  AND2_X1 U575 ( .A1(n516), .A2(n649), .ZN(n523) );
  INV_X1 U576 ( .A(n516), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n643), .B(n529), .ZN(n528) );
  INV_X1 U578 ( .A(KEYINPUT95), .ZN(n529) );
  XNOR2_X2 U579 ( .A(n530), .B(KEYINPUT17), .ZN(n888) );
  INV_X1 U580 ( .A(KEYINPUT94), .ZN(n639) );
  INV_X1 U581 ( .A(KEYINPUT96), .ZN(n648) );
  NOR2_X2 U582 ( .A1(G2105), .A2(n546), .ZN(n890) );
  XOR2_X1 U583 ( .A(KEYINPUT69), .B(n541), .Z(G299) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n588) );
  NAND2_X1 U585 ( .A1(n804), .A2(G53), .ZN(n540) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n798) );
  NAND2_X1 U587 ( .A1(G91), .A2(n798), .ZN(n533) );
  INV_X1 U588 ( .A(G651), .ZN(n534) );
  NOR2_X1 U589 ( .A1(n588), .A2(n534), .ZN(n803) );
  NAND2_X1 U590 ( .A1(G78), .A2(n803), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n538) );
  NOR2_X1 U592 ( .A1(G543), .A2(n534), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n800), .A2(G65), .ZN(n536) );
  XOR2_X1 U594 ( .A(KEYINPUT68), .B(n536), .Z(n537) );
  NOR2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U597 ( .A1(G101), .A2(n890), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n542), .Z(n545) );
  NAND2_X1 U599 ( .A1(G137), .A2(n888), .ZN(n543) );
  XOR2_X1 U600 ( .A(n543), .B(KEYINPUT65), .Z(n544) );
  AND2_X1 U601 ( .A1(n546), .A2(G2105), .ZN(n894) );
  NAND2_X1 U602 ( .A1(G125), .A2(n894), .ZN(n548) );
  AND2_X1 U603 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U604 ( .A1(G113), .A2(n897), .ZN(n547) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U606 ( .A(G120), .ZN(G236) );
  NAND2_X1 U607 ( .A1(G64), .A2(n800), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G52), .A2(n804), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n798), .A2(G90), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT67), .B(n551), .Z(n553) );
  NAND2_X1 U612 ( .A1(n803), .A2(G77), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U615 ( .A1(n556), .A2(n555), .ZN(G171) );
  NAND2_X1 U616 ( .A1(G126), .A2(n894), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G138), .A2(n888), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G114), .A2(n897), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G102), .A2(n890), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT85), .B(n563), .Z(G164) );
  NAND2_X1 U624 ( .A1(n798), .A2(G89), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G76), .A2(n803), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G63), .A2(n800), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G51), .A2(n804), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U636 ( .A(G171), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G75), .A2(n803), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G62), .A2(n800), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G88), .A2(n798), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT79), .B(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n804), .A2(G50), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(G303) );
  INV_X1 U645 ( .A(G303), .ZN(G166) );
  NAND2_X1 U646 ( .A1(G85), .A2(n798), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G60), .A2(n800), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G72), .A2(n803), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G47), .A2(n804), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT66), .B(n587), .Z(G290) );
  NAND2_X1 U654 ( .A1(G87), .A2(n588), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G74), .A2(G651), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U657 ( .A1(n800), .A2(n591), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G49), .A2(n804), .ZN(n592) );
  XOR2_X1 U659 ( .A(KEYINPUT77), .B(n592), .Z(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(G288) );
  NAND2_X1 U661 ( .A1(G48), .A2(n804), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n595), .B(KEYINPUT78), .ZN(n602) );
  NAND2_X1 U663 ( .A1(G86), .A2(n798), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G61), .A2(n800), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n803), .A2(G73), .ZN(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT2), .B(n598), .Z(n599) );
  NOR2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(G305) );
  NAND2_X1 U670 ( .A1(G79), .A2(n803), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G54), .A2(n804), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U673 ( .A(KEYINPUT72), .B(n605), .ZN(n609) );
  NAND2_X1 U674 ( .A1(G92), .A2(n798), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G66), .A2(n800), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  XNOR2_X1 U678 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n611), .B(n610), .ZN(n796) );
  NAND2_X1 U680 ( .A1(G56), .A2(n800), .ZN(n612) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n612), .Z(n618) );
  NAND2_X1 U682 ( .A1(n798), .A2(G81), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT12), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G68), .A2(n803), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT13), .B(n616), .Z(n617) );
  NOR2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n804), .A2(G43), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n999) );
  NOR2_X1 U690 ( .A1(G164), .A2(G1384), .ZN(n688) );
  INV_X1 U691 ( .A(G1996), .ZN(n1018) );
  XOR2_X1 U692 ( .A(n622), .B(KEYINPUT26), .Z(n624) );
  NAND2_X1 U693 ( .A1(n670), .A2(G1341), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U695 ( .A1(n999), .A2(n625), .ZN(n626) );
  OR2_X1 U696 ( .A1(n796), .A2(n626), .ZN(n634) );
  NAND2_X1 U697 ( .A1(n796), .A2(n626), .ZN(n632) );
  INV_X1 U698 ( .A(KEYINPUT91), .ZN(n627) );
  INV_X1 U699 ( .A(n650), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G2067), .A2(n628), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G1348), .A2(n670), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n642) );
  XOR2_X1 U705 ( .A(G1956), .B(KEYINPUT93), .Z(n934) );
  NAND2_X1 U706 ( .A1(n650), .A2(n934), .ZN(n644) );
  INV_X1 U707 ( .A(G299), .ZN(n635) );
  AND2_X1 U708 ( .A1(n644), .A2(n635), .ZN(n638) );
  INV_X1 U709 ( .A(G2072), .ZN(n1012) );
  XNOR2_X1 U710 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(n645) );
  AND2_X1 U712 ( .A1(n638), .A2(n645), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U716 ( .A1(G299), .A2(n646), .ZN(n647) );
  XOR2_X1 U717 ( .A(G2078), .B(KEYINPUT25), .Z(n1013) );
  NOR2_X1 U718 ( .A1(n1013), .A2(n650), .ZN(n653) );
  INV_X1 U719 ( .A(n670), .ZN(n651) );
  NOR2_X1 U720 ( .A1(n651), .A2(G1961), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U722 ( .A1(G8), .A2(n670), .ZN(n745) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n745), .ZN(n664) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n670), .ZN(n666) );
  NOR2_X1 U725 ( .A1(n664), .A2(n666), .ZN(n654) );
  NAND2_X1 U726 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U728 ( .A1(G168), .A2(n656), .ZN(n659) );
  AND2_X1 U729 ( .A1(G301), .A2(n657), .ZN(n658) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(KEYINPUT31), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT97), .ZN(n669) );
  INV_X1 U734 ( .A(n669), .ZN(n665) );
  NOR2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U736 ( .A1(G8), .A2(n666), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n730) );
  AND2_X1 U738 ( .A1(n669), .A2(G286), .ZN(n678) );
  INV_X1 U739 ( .A(G8), .ZN(n676) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(KEYINPUT98), .ZN(n673) );
  NOR2_X1 U742 ( .A1(n745), .A2(G1971), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n674), .A2(G303), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n680) );
  XOR2_X1 U747 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(n732) );
  NAND2_X1 U749 ( .A1(n730), .A2(n732), .ZN(n683) );
  NAND2_X1 U750 ( .A1(G166), .A2(G8), .ZN(n681) );
  OR2_X1 U751 ( .A1(G2090), .A2(n681), .ZN(n682) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n685) );
  INV_X1 U753 ( .A(KEYINPUT103), .ZN(n684) );
  XNOR2_X1 U754 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n686), .A2(n745), .ZN(n728) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U757 ( .A(KEYINPUT86), .B(n689), .Z(n761) );
  NAND2_X1 U758 ( .A1(G128), .A2(n894), .ZN(n691) );
  NAND2_X1 U759 ( .A1(G116), .A2(n897), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT35), .ZN(n697) );
  NAND2_X1 U762 ( .A1(G140), .A2(n888), .ZN(n694) );
  NAND2_X1 U763 ( .A1(G104), .A2(n890), .ZN(n693) );
  NAND2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U765 ( .A(KEYINPUT34), .B(n695), .Z(n696) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n698), .B(KEYINPUT36), .ZN(n882) );
  XOR2_X1 U768 ( .A(G2067), .B(KEYINPUT37), .Z(n699) );
  NOR2_X1 U769 ( .A1(n882), .A2(n699), .ZN(n955) );
  NAND2_X1 U770 ( .A1(n882), .A2(n699), .ZN(n760) );
  INV_X1 U771 ( .A(n760), .ZN(n956) );
  NAND2_X1 U772 ( .A1(G105), .A2(n890), .ZN(n700) );
  XNOR2_X1 U773 ( .A(n700), .B(KEYINPUT38), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G129), .A2(n894), .ZN(n702) );
  NAND2_X1 U775 ( .A1(G117), .A2(n897), .ZN(n701) );
  NAND2_X1 U776 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U777 ( .A1(G141), .A2(n888), .ZN(n703) );
  XNOR2_X1 U778 ( .A(KEYINPUT87), .B(n703), .ZN(n704) );
  NOR2_X1 U779 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U780 ( .A1(n707), .A2(n706), .ZN(n881) );
  NOR2_X1 U781 ( .A1(G1996), .A2(n881), .ZN(n966) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n881), .ZN(n715) );
  NAND2_X1 U783 ( .A1(G119), .A2(n894), .ZN(n709) );
  NAND2_X1 U784 ( .A1(G131), .A2(n888), .ZN(n708) );
  NAND2_X1 U785 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U786 ( .A1(G107), .A2(n897), .ZN(n711) );
  NAND2_X1 U787 ( .A1(G95), .A2(n890), .ZN(n710) );
  NAND2_X1 U788 ( .A1(n711), .A2(n710), .ZN(n712) );
  OR2_X1 U789 ( .A1(n713), .A2(n712), .ZN(n902) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n902), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U792 ( .A(KEYINPUT88), .B(n716), .Z(n959) );
  NOR2_X1 U793 ( .A1(n761), .A2(n959), .ZN(n759) );
  NOR2_X1 U794 ( .A1(G1986), .A2(G290), .ZN(n718) );
  NOR2_X1 U795 ( .A1(G1991), .A2(n902), .ZN(n717) );
  XNOR2_X1 U796 ( .A(KEYINPUT104), .B(n717), .ZN(n962) );
  NOR2_X1 U797 ( .A1(n718), .A2(n962), .ZN(n719) );
  XOR2_X1 U798 ( .A(KEYINPUT105), .B(n719), .Z(n720) );
  NOR2_X1 U799 ( .A1(n759), .A2(n720), .ZN(n721) );
  NOR2_X1 U800 ( .A1(n966), .A2(n721), .ZN(n722) );
  XOR2_X1 U801 ( .A(KEYINPUT39), .B(n722), .Z(n723) );
  NOR2_X1 U802 ( .A1(n956), .A2(n723), .ZN(n724) );
  NOR2_X1 U803 ( .A1(n955), .A2(n724), .ZN(n725) );
  NOR2_X1 U804 ( .A1(n761), .A2(n725), .ZN(n726) );
  XNOR2_X1 U805 ( .A(n726), .B(KEYINPUT106), .ZN(n767) );
  INV_X1 U806 ( .A(n767), .ZN(n727) );
  AND2_X1 U807 ( .A1(n728), .A2(n727), .ZN(n758) );
  NAND2_X1 U808 ( .A1(G288), .A2(G1976), .ZN(n729) );
  XNOR2_X1 U809 ( .A(n729), .B(KEYINPUT101), .ZN(n1004) );
  NOR2_X1 U810 ( .A1(n1004), .A2(n745), .ZN(n733) );
  AND2_X1 U811 ( .A1(n730), .A2(n733), .ZN(n731) );
  NAND2_X1 U812 ( .A1(n732), .A2(n731), .ZN(n738) );
  INV_X1 U813 ( .A(n733), .ZN(n736) );
  NOR2_X1 U814 ( .A1(G1971), .A2(G303), .ZN(n735) );
  NOR2_X1 U815 ( .A1(G288), .A2(G1976), .ZN(n734) );
  XNOR2_X1 U816 ( .A(n734), .B(KEYINPUT100), .ZN(n746) );
  NOR2_X1 U817 ( .A1(n735), .A2(n746), .ZN(n991) );
  OR2_X1 U818 ( .A1(n736), .A2(n991), .ZN(n737) );
  AND2_X1 U819 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U820 ( .A(n739), .B(KEYINPUT64), .ZN(n744) );
  INV_X1 U821 ( .A(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n740) );
  XOR2_X1 U823 ( .A(n740), .B(KEYINPUT90), .Z(n741) );
  XNOR2_X1 U824 ( .A(KEYINPUT24), .B(n741), .ZN(n742) );
  OR2_X1 U825 ( .A1(n745), .A2(n742), .ZN(n754) );
  AND2_X1 U826 ( .A1(n749), .A2(n754), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n744), .A2(n743), .ZN(n756) );
  INV_X1 U828 ( .A(n745), .ZN(n747) );
  NAND2_X1 U829 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U830 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U831 ( .A(n750), .B(KEYINPUT102), .Z(n752) );
  XNOR2_X1 U832 ( .A(G1981), .B(G305), .ZN(n986) );
  INV_X1 U833 ( .A(n986), .ZN(n751) );
  NAND2_X1 U834 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U835 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U836 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U837 ( .A1(n758), .A2(n757), .ZN(n769) );
  INV_X1 U838 ( .A(n759), .ZN(n765) );
  XOR2_X1 U839 ( .A(G1986), .B(G290), .Z(n1003) );
  NAND2_X1 U840 ( .A1(n760), .A2(n1003), .ZN(n763) );
  INV_X1 U841 ( .A(n761), .ZN(n762) );
  NAND2_X1 U842 ( .A1(n763), .A2(n762), .ZN(n764) );
  AND2_X1 U843 ( .A1(n765), .A2(n764), .ZN(n766) );
  OR2_X1 U844 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U845 ( .A1(n769), .A2(n768), .ZN(n771) );
  INV_X1 U846 ( .A(KEYINPUT40), .ZN(n770) );
  XNOR2_X1 U847 ( .A(n771), .B(n770), .ZN(G329) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U849 ( .A(n772), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n838) );
  NAND2_X1 U851 ( .A1(n838), .A2(G567), .ZN(n773) );
  XNOR2_X1 U852 ( .A(n773), .B(KEYINPUT11), .ZN(n774) );
  XNOR2_X1 U853 ( .A(KEYINPUT71), .B(n774), .ZN(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n780) );
  OR2_X1 U855 ( .A1(n999), .A2(n780), .ZN(G153) );
  INV_X1 U856 ( .A(n796), .ZN(n996) );
  NOR2_X1 U857 ( .A1(G868), .A2(n996), .ZN(n776) );
  INV_X1 U858 ( .A(G868), .ZN(n818) );
  NOR2_X1 U859 ( .A1(n818), .A2(G301), .ZN(n775) );
  NOR2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U861 ( .A(KEYINPUT74), .B(n777), .ZN(G284) );
  NAND2_X1 U862 ( .A1(G286), .A2(G868), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G299), .A2(n818), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U865 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n781), .A2(n796), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U868 ( .A1(G868), .A2(n999), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G868), .A2(n796), .ZN(n783) );
  NOR2_X1 U870 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U872 ( .A(KEYINPUT75), .B(n786), .Z(G282) );
  NAND2_X1 U873 ( .A1(n894), .A2(G123), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT18), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G111), .A2(n897), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G135), .A2(n888), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G99), .A2(n890), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n958) );
  XNOR2_X1 U881 ( .A(n958), .B(G2096), .ZN(n795) );
  INV_X1 U882 ( .A(G2100), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(G156) );
  NAND2_X1 U884 ( .A1(G559), .A2(n796), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n999), .B(n797), .ZN(n815) );
  NOR2_X1 U886 ( .A1(n815), .A2(G860), .ZN(n809) );
  NAND2_X1 U887 ( .A1(n798), .A2(G93), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT76), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G67), .A2(n800), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G80), .A2(n803), .ZN(n806) );
  NAND2_X1 U892 ( .A1(G55), .A2(n804), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n817) );
  XNOR2_X1 U895 ( .A(n809), .B(n817), .ZN(G145) );
  XNOR2_X1 U896 ( .A(G166), .B(KEYINPUT19), .ZN(n814) );
  XNOR2_X1 U897 ( .A(n817), .B(G288), .ZN(n812) );
  XOR2_X1 U898 ( .A(G290), .B(G299), .Z(n810) );
  XNOR2_X1 U899 ( .A(G305), .B(n810), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n814), .B(n813), .ZN(n906) );
  XOR2_X1 U902 ( .A(n815), .B(n906), .Z(n816) );
  NAND2_X1 U903 ( .A1(n816), .A2(G868), .ZN(n820) );
  NAND2_X1 U904 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U906 ( .A(KEYINPUT80), .B(n821), .Z(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U911 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XOR2_X1 U912 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U914 ( .A1(G661), .A2(G483), .ZN(n836) );
  NOR2_X1 U915 ( .A1(G237), .A2(G236), .ZN(n826) );
  NAND2_X1 U916 ( .A1(G69), .A2(n826), .ZN(n827) );
  XNOR2_X1 U917 ( .A(KEYINPUT83), .B(n827), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n828), .A2(G108), .ZN(n927) );
  NAND2_X1 U919 ( .A1(n927), .A2(G567), .ZN(n835) );
  XOR2_X1 U920 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n830) );
  NAND2_X1 U921 ( .A1(G132), .A2(G82), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n830), .B(n829), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n831), .A2(G218), .ZN(n832) );
  NAND2_X1 U924 ( .A1(G96), .A2(n832), .ZN(n926) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n926), .ZN(n833) );
  XNOR2_X1 U926 ( .A(KEYINPUT82), .B(n833), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(n844) );
  NOR2_X1 U928 ( .A1(n836), .A2(n844), .ZN(n837) );
  XNOR2_X1 U929 ( .A(n837), .B(KEYINPUT84), .ZN(n842) );
  NAND2_X1 U930 ( .A1(G36), .A2(n842), .ZN(G176) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n838), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  XNOR2_X1 U933 ( .A(KEYINPUT107), .B(n839), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n840), .A2(G661), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(KEYINPUT108), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(G188) );
  XNOR2_X1 U938 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  INV_X1 U939 ( .A(n844), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1986), .B(G1976), .Z(n854) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1956), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U952 ( .A(n855), .B(G2474), .Z(n857) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1981), .Z(n859) );
  XNOR2_X1 U956 ( .A(G1961), .B(G1971), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U959 ( .A1(n894), .A2(G124), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U961 ( .A1(G136), .A2(n888), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U963 ( .A(KEYINPUT110), .B(n865), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G112), .A2(n897), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G100), .A2(n890), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n879) );
  NAND2_X1 U969 ( .A1(G139), .A2(n888), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G103), .A2(n890), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U972 ( .A1(n894), .A2(G127), .ZN(n872) );
  XOR2_X1 U973 ( .A(KEYINPUT113), .B(n872), .Z(n874) );
  NAND2_X1 U974 ( .A1(n897), .A2(G115), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n969) );
  XNOR2_X1 U978 ( .A(n969), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n887) );
  XOR2_X1 U980 ( .A(G162), .B(n958), .Z(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n883) );
  XOR2_X1 U982 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U983 ( .A(G164), .B(G160), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n904) );
  NAND2_X1 U986 ( .A1(n888), .A2(G142), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(KEYINPUT112), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G106), .A2(n890), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n893), .B(KEYINPUT45), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G130), .A2(n894), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G118), .A2(n897), .ZN(n898) );
  XNOR2_X1 U994 ( .A(KEYINPUT111), .B(n898), .ZN(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n906), .B(KEYINPUT115), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(n999), .B(G286), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1002 ( .A(n996), .B(G171), .Z(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n911), .ZN(G397) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2430), .Z(n913) );
  XNOR2_X1 U1006 ( .A(G2438), .B(G2443), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n919) );
  XOR2_X1 U1008 ( .A(G2435), .B(G2454), .Z(n915) );
  XNOR2_X1 U1009 ( .A(G1341), .B(G1348), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1011 ( .A(G2446), .B(G2427), .Z(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1013 ( .A(n919), .B(n918), .Z(n920) );
  NAND2_X1 U1014 ( .A1(G14), .A2(n920), .ZN(n928) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n928), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(G225) );
  XOR2_X1 U1021 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1023 ( .A(G132), .ZN(G219) );
  INV_X1 U1024 ( .A(G108), .ZN(G238) );
  INV_X1 U1025 ( .A(G96), .ZN(G221) );
  INV_X1 U1026 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(G325) );
  INV_X1 U1028 ( .A(G325), .ZN(G261) );
  INV_X1 U1029 ( .A(n928), .ZN(G401) );
  XNOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(n929), .B(G4), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(G6), .B(G1981), .ZN(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(G20), .B(n934), .ZN(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT60), .B(n937), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G21), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(G5), .B(G1961), .ZN(n938) );
  NOR2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1971), .B(G22), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(G23), .B(G1976), .ZN(n942) );
  NOR2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1046 ( .A(G1986), .B(KEYINPUT126), .Z(n944) );
  XNOR2_X1 U1047 ( .A(G24), .B(n944), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(n947), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1051 ( .A(KEYINPUT61), .B(n950), .Z(n952) );
  XOR2_X1 U1052 ( .A(G16), .B(KEYINPUT125), .Z(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(KEYINPUT127), .B(n953), .ZN(n954) );
  NAND2_X1 U1055 ( .A1(n954), .A2(G11), .ZN(n984) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G2084), .B(G160), .Z(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n977) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1064 ( .A(KEYINPUT117), .B(n967), .Z(n968) );
  XOR2_X1 U1065 ( .A(KEYINPUT51), .B(n968), .Z(n975) );
  XOR2_X1 U1066 ( .A(G164), .B(G2078), .Z(n972) );
  XOR2_X1 U1067 ( .A(n969), .B(KEYINPUT118), .Z(n970) );
  XNOR2_X1 U1068 ( .A(G2072), .B(n970), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(KEYINPUT50), .B(n973), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT52), .ZN(n980) );
  INV_X1 U1074 ( .A(KEYINPUT55), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(G29), .A2(n981), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT119), .B(n982), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n1011) );
  XNOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XOR2_X1 U1080 ( .A(G1966), .B(G168), .Z(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(n987), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(n988), .B(KEYINPUT57), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G1956), .B(KEYINPUT124), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(n989), .B(G299), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(G1971), .A2(G303), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n996), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G301), .B(G1961), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n999), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1036) );
  XOR2_X1 U1100 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n1027) );
  XNOR2_X1 U1101 ( .A(G1991), .B(G25), .ZN(n1024) );
  XNOR2_X1 U1102 ( .A(G33), .B(n1012), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1013), .B(G27), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G2067), .B(G26), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(G32), .B(n1018), .Z(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT120), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(KEYINPUT121), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(G28), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(n1027), .B(n1026), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(G2090), .B(G35), .Z(n1030) );
  XOR2_X1 U1115 ( .A(KEYINPUT54), .B(G34), .Z(n1028) );
  XNOR2_X1 U1116 ( .A(n1028), .B(G2084), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1119 ( .A(KEYINPUT55), .B(n1033), .Z(n1034) );
  NOR2_X1 U1120 ( .A1(G29), .A2(n1034), .ZN(n1035) );
  NOR2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1122 ( .A(n1037), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

