//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT10), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(KEYINPUT68), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n189), .A2(KEYINPUT69), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n192), .A2(new_n194), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n188), .B1(new_n199), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT3), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n212), .B2(G104), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(KEYINPUT81), .A3(G107), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n210), .A2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n212), .A2(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n219), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n212), .A2(KEYINPUT3), .A3(G104), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(new_n212), .B2(G104), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n217), .A2(new_n218), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n219), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT0), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(new_n189), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n206), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(KEYINPUT0), .B2(G128), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n189), .A3(KEYINPUT64), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n237), .A2(new_n238), .B1(new_n192), .B2(new_n194), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n235), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n241), .B(G101), .C1(new_n229), .C2(new_n230), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n232), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n226), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n219), .A2(new_n223), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n204), .A2(G128), .B1(new_n192), .B2(new_n194), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n197), .B2(new_n198), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n188), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT82), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(new_n188), .C1(new_n245), .C2(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT67), .A3(G131), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT66), .B(G131), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n261), .A2(new_n256), .A3(new_n255), .A4(new_n258), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT67), .B1(new_n259), .B2(G131), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n244), .A2(new_n252), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(G227), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(KEYINPUT84), .A3(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n245), .A2(new_n247), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n245), .A2(new_n199), .A3(new_n207), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n265), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT12), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT84), .B1(new_n266), .B2(new_n271), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n187), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n244), .B2(new_n252), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n266), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n271), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT84), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT85), .A3(new_n276), .A4(new_n272), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n271), .B1(new_n276), .B2(new_n266), .ZN(new_n292));
  INV_X1    g106(.A(new_n284), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n281), .ZN(new_n294));
  OAI21_X1  g108(.A(G469), .B1(new_n294), .B2(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G237), .A2(G953), .ZN(new_n297));
  AND2_X1   g111(.A1(KEYINPUT93), .A2(G143), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT93), .A2(G143), .ZN(new_n299));
  OAI211_X1 g113(.A(G214), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G237), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n268), .A3(G214), .ZN(new_n302));
  NAND2_X1  g116(.A1(KEYINPUT93), .A2(G143), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n261), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT95), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT17), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n310), .A3(new_n306), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n300), .A2(new_n304), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n261), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n308), .A2(new_n309), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n317), .A2(G140), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(KEYINPUT16), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n191), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n316), .B(G146), .C1(KEYINPUT16), .C2(new_n318), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n310), .B1(new_n305), .B2(new_n306), .ZN(new_n323));
  AOI211_X1 g137(.A(KEYINPUT95), .B(new_n261), .C1(new_n300), .C2(new_n304), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT17), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n314), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT18), .A2(G131), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT94), .B1(new_n312), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT94), .ZN(new_n329));
  INV_X1    g143(.A(new_n327), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n305), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n312), .A2(new_n327), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n315), .B(new_n191), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G113), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n210), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n326), .A2(new_n338), .A3(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n290), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(G475), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G475), .A2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT19), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n315), .B(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n321), .B1(new_n349), .B2(G146), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n323), .A2(new_n324), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(new_n313), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n334), .B1(new_n330), .B2(new_n305), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n331), .B2(new_n328), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n339), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g169(.A(KEYINPUT20), .B(new_n347), .C1(new_n341), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n341), .A2(KEYINPUT96), .A3(new_n355), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT96), .B1(new_n341), .B2(new_n355), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n358), .A2(new_n359), .A3(new_n347), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(G116), .B(G122), .Z(new_n363));
  INV_X1    g177(.A(G122), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G116), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n212), .B1(new_n365), .B2(KEYINPUT14), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n363), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT69), .B(G128), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G143), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n193), .A2(G128), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n254), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n370), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G134), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n367), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n363), .B(G107), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT13), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n370), .B(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n203), .A2(new_n193), .ZN(new_n378));
  OAI21_X1  g192(.A(G134), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n379), .A3(new_n371), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n375), .A2(new_n379), .A3(KEYINPUT97), .A4(new_n371), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n374), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  INV_X1    g199(.A(G217), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n385), .A2(new_n386), .A3(G953), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n387), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n389), .B(new_n374), .C1(new_n382), .C2(new_n383), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n290), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G478), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n391), .B(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n345), .A2(new_n362), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n296), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n268), .A2(G952), .ZN(new_n400));
  INV_X1    g214(.A(G234), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n301), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n290), .B(new_n268), .C1(G234), .C2(G237), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT21), .B(G898), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G214), .B1(G237), .B2(G902), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n408), .B(KEYINPUT86), .Z(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n199), .A2(new_n207), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n317), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n240), .A2(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT90), .B(G224), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n415), .A2(new_n268), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n414), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G116), .B(G119), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT71), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT2), .ZN(new_n426));
  INV_X1    g240(.A(G113), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT70), .B1(KEYINPUT2), .B2(G113), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT2), .A2(G113), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n424), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g247(.A(KEYINPUT72), .B(new_n431), .C1(new_n428), .C2(new_n429), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n423), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n429), .ZN(new_n436));
  NOR3_X1   g250(.A1(KEYINPUT70), .A2(KEYINPUT2), .A3(G113), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT72), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n431), .B1(new_n428), .B2(new_n429), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n424), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n422), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n242), .A4(new_n232), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n446));
  INV_X1    g260(.A(G119), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(G116), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n427), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n446), .A2(new_n450), .B1(new_n440), .B2(new_n421), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n224), .B2(new_n225), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n232), .A2(new_n242), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n444), .B1(new_n454), .B2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n420), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT89), .B1(new_n456), .B2(KEYINPUT6), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n435), .A2(new_n442), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n232), .A2(new_n242), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT87), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n452), .A3(new_n445), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n420), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n461), .B2(new_n420), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n460), .A2(new_n419), .A3(new_n452), .A4(new_n445), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND4_X1   g283(.A1(new_n466), .A2(new_n456), .A3(KEYINPUT6), .A4(new_n468), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n418), .B(new_n465), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G210), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n414), .B1(new_n473), .B2(new_n416), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n412), .A2(KEYINPUT7), .A3(new_n417), .A4(new_n413), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n440), .A2(new_n421), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n446), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n450), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n446), .A2(new_n477), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n219), .A3(new_n223), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n419), .B(KEYINPUT8), .Z(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n451), .B2(new_n245), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n474), .A2(new_n475), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n485), .B2(new_n468), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n471), .A2(new_n472), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n472), .B1(new_n471), .B2(new_n488), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n407), .B(new_n410), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n240), .B1(new_n263), .B2(new_n264), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n257), .A2(G134), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n256), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G131), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n262), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n411), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n492), .B1(new_n499), .B2(new_n458), .ZN(new_n500));
  AND4_X1   g314(.A1(new_n492), .A2(new_n458), .A3(new_n498), .A4(new_n493), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n499), .A2(new_n458), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G101), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n297), .A2(G210), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT74), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n507), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n504), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n238), .A2(new_n237), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n234), .B1(new_n516), .B2(new_n206), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n206), .A2(new_n234), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n235), .B(KEYINPUT65), .C1(new_n239), .C2(new_n234), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n498), .B1(new_n521), .B2(new_n265), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n493), .A2(new_n498), .A3(KEYINPUT30), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n443), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n499), .A2(new_n458), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n512), .B1(new_n528), .B2(new_n510), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n443), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n500), .B2(new_n501), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n511), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n514), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n527), .A3(new_n510), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n511), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n526), .A2(new_n538), .A3(new_n527), .A4(new_n510), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n534), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n315), .A2(new_n191), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n321), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n368), .A2(G119), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n189), .A2(G119), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n548), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT75), .B(new_n550), .C1(new_n368), .C2(G119), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT24), .B(G110), .Z(new_n554));
  NOR3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT76), .B1(new_n447), .B2(G128), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT76), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n189), .A3(G119), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT23), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n556), .B(new_n558), .C1(new_n550), .C2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT23), .A4(G119), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G110), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n547), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(KEYINPUT77), .A3(new_n561), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(KEYINPUT78), .A3(new_n568), .A4(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n320), .A2(new_n321), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n554), .B1(new_n552), .B2(new_n553), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G110), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n562), .B2(new_n566), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT78), .B1(new_n574), .B2(new_n568), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n564), .B(new_n565), .C1(new_n572), .C2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT79), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT22), .B(G137), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n549), .A2(new_n551), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n549), .A2(new_n548), .A3(new_n551), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n586), .A2(new_n554), .B1(new_n320), .B2(new_n321), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n574), .A2(new_n568), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n590), .A3(new_n569), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n565), .B1(new_n591), .B2(new_n564), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n564), .B1(new_n572), .B2(new_n575), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n580), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n290), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT25), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n594), .A2(KEYINPUT80), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n576), .A3(new_n581), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n595), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT25), .A3(new_n290), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n386), .B1(G234), .B2(new_n290), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(G902), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n604), .A2(new_n605), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n545), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n399), .A2(new_n491), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n215), .ZN(G3));
  NAND2_X1  g424(.A1(new_n540), .A2(new_n290), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n540), .A2(new_n542), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT25), .B1(new_n602), .B2(new_n290), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n598), .B(G902), .C1(new_n601), .C2(new_n595), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n605), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n602), .A2(new_n606), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n398), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n291), .B2(new_n295), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n345), .A2(new_n362), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n392), .A2(new_n290), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n391), .B2(G478), .ZN(new_n629));
  OR3_X1    g443(.A1(new_n388), .A2(new_n390), .A3(KEYINPUT33), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT33), .B1(new_n388), .B2(new_n390), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n629), .B1(new_n633), .B2(G478), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n625), .B1(new_n491), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n471), .A2(new_n488), .ZN(new_n638));
  INV_X1    g452(.A(new_n472), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n471), .A2(new_n472), .A3(new_n488), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n409), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(KEYINPUT98), .A3(new_n407), .A4(new_n635), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n624), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  XNOR2_X1  g460(.A(new_n360), .B(KEYINPUT20), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n344), .A3(new_n395), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n491), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n624), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(new_n491), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n621), .B(new_n396), .C1(new_n291), .C2(new_n295), .ZN(new_n655));
  INV_X1    g469(.A(new_n605), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n599), .B2(new_n603), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n594), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n606), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT99), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n617), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n614), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n654), .A2(new_n655), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT100), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT37), .B(G110), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  INV_X1    g483(.A(new_n544), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n662), .A2(new_n664), .B1(new_n672), .B2(new_n534), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n404), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n402), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n648), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n677), .A3(new_n642), .A4(new_n622), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT101), .B(G128), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G30));
  XNOR2_X1  g494(.A(new_n676), .B(KEYINPUT39), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n622), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT40), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n489), .A2(new_n490), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n662), .A2(new_n664), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n528), .A2(new_n511), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n527), .A2(new_n511), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n290), .B1(new_n691), .B2(new_n503), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n672), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n395), .B1(new_n345), .B2(new_n362), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n410), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n683), .A2(new_n687), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT103), .B(G143), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G45));
  NAND3_X1  g513(.A1(new_n626), .A2(new_n634), .A3(new_n676), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n673), .A2(new_n642), .A3(new_n622), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(new_n288), .A2(new_n290), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n398), .A3(new_n291), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n608), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n637), .A2(new_n643), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n637), .A2(new_n643), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND2_X1  g528(.A1(new_n707), .A2(new_n650), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT105), .B(G116), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G18));
  AND3_X1   g531(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n621), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n396), .A2(new_n406), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n673), .A2(new_n642), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT106), .B(G119), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G21));
  OAI211_X1 g538(.A(new_n695), .B(new_n410), .C1(new_n489), .C2(new_n490), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n536), .B(new_n539), .C1(new_n510), .C2(new_n504), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n542), .B(KEYINPUT107), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n612), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n619), .A3(new_n406), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n726), .A2(new_n720), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  AOI21_X1  g547(.A(new_n730), .B1(new_n662), .B2(new_n664), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n720), .A3(new_n642), .A4(new_n701), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(new_n608), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n293), .A2(KEYINPUT108), .A3(new_n281), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n284), .B2(new_n280), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n292), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(G902), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n291), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n291), .A2(KEYINPUT109), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n621), .A2(new_n409), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n489), .A2(new_n490), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n738), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n291), .A2(KEYINPUT109), .A3(new_n743), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT109), .B1(new_n291), .B2(new_n743), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n751), .B(new_n738), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n737), .B(new_n701), .C1(new_n752), .C2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n608), .B1(new_n761), .B2(new_n755), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  OAI211_X1 g579(.A(new_n737), .B(new_n677), .C1(new_n752), .C2(new_n756), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  OAI21_X1  g581(.A(G469), .B1(new_n294), .B2(KEYINPUT45), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(KEYINPUT111), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(G469), .A2(G902), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n718), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n773), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n777), .A2(new_n398), .A3(new_n681), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n640), .A2(new_n641), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n409), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n634), .A2(new_n345), .A3(new_n362), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT43), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n614), .A3(new_n688), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n781), .B1(new_n785), .B2(KEYINPUT44), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n778), .B(new_n786), .C1(KEYINPUT44), .C2(new_n785), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  NOR4_X1   g602(.A1(new_n781), .A2(new_n545), .A3(new_n607), .A4(new_n700), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n777), .A2(KEYINPUT47), .A3(new_n398), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT47), .B1(new_n777), .B2(new_n398), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n705), .A2(new_n291), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT49), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n694), .A3(new_n782), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n619), .A2(new_n750), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(KEYINPUT49), .B2(new_n794), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(KEYINPUT112), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n687), .A2(new_n796), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n647), .A2(new_n344), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n395), .A2(new_n676), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n684), .A2(new_n410), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n622), .A3(new_n673), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n734), .A2(new_n701), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n752), .B2(new_n756), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n766), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n759), .B2(new_n763), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n626), .A2(new_n395), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n654), .A2(new_n622), .A3(new_n620), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n715), .A2(new_n814), .A3(new_n722), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n666), .A2(new_n732), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n779), .A2(new_n407), .A3(new_n410), .A4(new_n635), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n623), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n819), .B2(new_n609), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n654), .A2(new_n622), .A3(new_n635), .A4(new_n620), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n654), .A2(new_n655), .A3(new_n737), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n817), .A2(new_n712), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n676), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n398), .B1(new_n827), .B2(KEYINPUT115), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n657), .A2(new_n661), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n748), .A2(new_n726), .A3(new_n694), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n678), .A3(new_n702), .A4(new_n735), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(new_n832), .B2(KEYINPUT116), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n812), .A2(new_n826), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n839));
  INV_X1    g653(.A(new_n811), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n678), .A2(new_n702), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n735), .A4(new_n831), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n832), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n826), .A2(new_n764), .A3(new_n840), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n837), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n838), .B2(KEYINPUT117), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n839), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n837), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n835), .A4(new_n826), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n794), .A2(new_n779), .A3(new_n402), .A4(new_n750), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(new_n783), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n737), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT48), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n855), .A2(new_n672), .A3(new_n607), .A4(new_n693), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n859), .A2(new_n636), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n730), .A2(new_n619), .A3(new_n402), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n783), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n642), .A3(new_n720), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n858), .A2(new_n400), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n409), .A2(new_n862), .A3(new_n687), .A4(new_n720), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT50), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(KEYINPUT50), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n856), .A2(new_n734), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n859), .A2(new_n626), .A3(new_n634), .ZN(new_n870));
  AND4_X1   g684(.A1(KEYINPUT51), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n862), .A2(new_n780), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT118), .ZN(new_n873));
  INV_X1    g687(.A(new_n790), .ZN(new_n874));
  INV_X1    g688(.A(new_n791), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n794), .A2(new_n398), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n864), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n877), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n875), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(new_n873), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n879), .B1(new_n885), .B2(KEYINPUT51), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n850), .A2(new_n854), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n801), .B1(new_n887), .B2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n268), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n290), .B1(new_n851), .B2(new_n852), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n418), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n891), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n893), .B2(new_n896), .ZN(G51));
  XNOR2_X1  g712(.A(new_n853), .B(KEYINPUT54), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n773), .B(KEYINPUT57), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n288), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n892), .A2(new_n770), .A3(new_n771), .A4(new_n769), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n890), .B1(new_n902), .B2(new_n903), .ZN(G54));
  NOR2_X1   g718(.A1(new_n358), .A2(new_n359), .ZN(new_n905));
  NAND2_X1  g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT120), .Z(new_n907));
  AND3_X1   g721(.A1(new_n892), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n892), .B2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n890), .ZN(G60));
  XOR2_X1   g724(.A(new_n627), .B(KEYINPUT59), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n899), .A2(new_n632), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n891), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n850), .B2(new_n854), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n633), .ZN(G63));
  NAND2_X1  g729(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n891), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n918));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT121), .Z(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n853), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n921), .ZN(new_n923));
  AOI211_X1 g737(.A(KEYINPUT122), .B(new_n923), .C1(new_n851), .C2(new_n852), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n602), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n659), .B1(new_n922), .B2(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n916), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n853), .A2(new_n921), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n853), .A2(new_n918), .A3(new_n921), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n926), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n917), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n916), .A2(new_n933), .A3(new_n928), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n929), .A2(new_n935), .ZN(G66));
  INV_X1    g750(.A(new_n405), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n268), .B1(new_n937), .B2(new_n415), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT124), .Z(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n826), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n894), .B1(G898), .B2(new_n268), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  NAND2_X1  g756(.A1(new_n524), .A2(new_n525), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n349), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n787), .A2(new_n792), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n841), .A2(new_n735), .ZN(new_n946));
  OR3_X1    g760(.A1(new_n946), .A2(new_n697), .A3(KEYINPUT62), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n946), .B2(new_n697), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n780), .B(new_n737), .C1(new_n635), .C2(new_n813), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(new_n682), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n945), .A2(new_n947), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n944), .B1(new_n951), .B2(new_n268), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n725), .A2(new_n608), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n946), .B1(new_n778), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n787), .A2(new_n792), .A3(new_n955), .A4(new_n766), .ZN(new_n956));
  INV_X1    g770(.A(new_n764), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n955), .A2(new_n766), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n945), .A2(new_n959), .A3(KEYINPUT126), .A4(new_n764), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n960), .A3(new_n268), .ZN(new_n961));
  INV_X1    g775(.A(new_n944), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT125), .B1(new_n961), .B2(new_n963), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n268), .B1(G227), .B2(G900), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  AOI221_X4 g782(.A(new_n952), .B1(KEYINPUT125), .B2(new_n968), .C1(new_n961), .C2(new_n963), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  NAND3_X1  g784(.A1(new_n958), .A2(new_n960), .A3(new_n826), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n511), .A3(new_n528), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n528), .B(new_n510), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n849), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n826), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n951), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n890), .B1(new_n980), .B2(new_n690), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n976), .A2(new_n978), .A3(new_n981), .ZN(G57));
endmodule


