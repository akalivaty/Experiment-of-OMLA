//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n591, new_n593, new_n594, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1084, new_n1085, new_n1086, new_n1087;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n462), .A2(KEYINPUT64), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(KEYINPUT64), .ZN(new_n469));
  NOR3_X1   g044(.A1(new_n468), .A2(new_n469), .A3(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT3), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(new_n461), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n467), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT65), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n474), .A2(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n472), .A2(G2105), .A3(new_n461), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(G124), .B2(new_n484), .ZN(G162));
  XOR2_X1   g060(.A(KEYINPUT66), .B(G114), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n473), .A2(G138), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT64), .B(G2104), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n461), .B(new_n493), .C1(new_n494), .C2(new_n460), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n472), .A2(KEYINPUT67), .A3(new_n461), .A4(new_n493), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n464), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n493), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n492), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT68), .B(G89), .Z(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT69), .Z(new_n523));
  INV_X1    g098(.A(new_n515), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(G51), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n510), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n513), .A2(new_n531), .B1(new_n515), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n507), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n513), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G81), .B1(G43), .B2(new_n524), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT72), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  XOR2_X1   g127(.A(new_n513), .B(KEYINPUT75), .Z(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT73), .Z(new_n558));
  NOR3_X1   g133(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT74), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n554), .B1(new_n510), .B2(new_n555), .C1(new_n558), .C2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n553), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n524), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT76), .Z(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n524), .A2(G48), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT77), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n510), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(G86), .B2(new_n553), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n541), .A2(G85), .B1(G47), .B2(new_n524), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n510), .B2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G301), .A2(G868), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n553), .A2(G92), .ZN(new_n579));
  XOR2_X1   g154(.A(new_n579), .B(KEYINPUT10), .Z(new_n580));
  NAND2_X1  g155(.A1(G79), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G66), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n507), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(G54), .A2(new_n524), .B1(new_n583), .B2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n578), .B1(new_n586), .B2(G868), .ZN(G284));
  OAI21_X1  g162(.A(new_n578), .B1(new_n586), .B2(G868), .ZN(G321));
  MUX2_X1   g163(.A(G299), .B(G286), .S(G868), .Z(G297));
  XOR2_X1   g164(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n586), .B1(new_n591), .B2(G860), .ZN(G148));
  NAND2_X1  g167(.A1(new_n586), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G868), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g170(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n596));
  XNOR2_X1  g171(.A(G323), .B(new_n596), .ZN(G282));
  OR2_X1    g172(.A1(G99), .A2(G2105), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n598), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n599));
  INV_X1    g174(.A(G135), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n474), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(G123), .B2(new_n484), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(G2096), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n470), .A2(new_n461), .A3(new_n463), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT13), .B(G2100), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT81), .Z(G156));
  XNOR2_X1  g185(.A(G2427), .B(G2438), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(G2430), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT15), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2435), .Z(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT14), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(G2451), .B(G2454), .Z(new_n618));
  XNOR2_X1  g193(.A(G2443), .B(G2446), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n617), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G1341), .B(G1348), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n621), .B(new_n622), .Z(new_n623));
  AND2_X1   g198(.A1(new_n623), .A2(G14), .ZN(G401));
  XOR2_X1   g199(.A(G2072), .B(G2078), .Z(new_n625));
  XOR2_X1   g200(.A(G2067), .B(G2678), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2084), .B(G2090), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n629), .B2(KEYINPUT18), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2100), .Z(new_n632));
  AND2_X1   g207(.A1(new_n629), .A2(KEYINPUT17), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n627), .A2(new_n628), .ZN(new_n634));
  AOI21_X1  g209(.A(KEYINPUT18), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(G227));
  XNOR2_X1  g211(.A(G1971), .B(G1976), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT19), .ZN(new_n638));
  XOR2_X1   g213(.A(G1956), .B(G2474), .Z(new_n639));
  XOR2_X1   g214(.A(G1961), .B(G1966), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT20), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n639), .A2(new_n640), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n645), .A2(new_n638), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT83), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n638), .A3(new_n641), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1991), .B(G1996), .ZN(new_n652));
  INV_X1    g227(.A(G1981), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G1986), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n651), .B(new_n655), .Z(G229));
  INV_X1    g231(.A(G16), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G21), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(G168), .B2(new_n657), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT93), .ZN(new_n660));
  INV_X1    g235(.A(G1966), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT24), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n663), .A2(G34), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(G34), .ZN(new_n665));
  AOI21_X1  g240(.A(G29), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n476), .B2(G29), .ZN(new_n667));
  INV_X1    g242(.A(G2084), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G29), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT30), .B(G28), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(G27), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(G164), .B2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(G2078), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(G29), .A2(G33), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G139), .ZN(new_n681));
  INV_X1    g256(.A(G127), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n464), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G115), .B2(G2104), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n680), .B1(new_n681), .B2(new_n474), .C1(new_n684), .C2(new_n473), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT90), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n677), .B1(new_n686), .B2(G29), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(G2072), .Z(new_n688));
  NAND4_X1  g263(.A1(new_n662), .A2(new_n672), .A3(new_n676), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n602), .A2(G29), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT94), .Z(new_n691));
  INV_X1    g266(.A(G11), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n660), .B2(new_n661), .ZN(new_n695));
  NOR4_X1   g270(.A1(new_n689), .A2(new_n691), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n670), .A2(G32), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n470), .A2(G105), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n484), .A2(G129), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  INV_X1    g277(.A(new_n474), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G141), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n699), .A2(new_n700), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT92), .Z(new_n706));
  OAI21_X1  g281(.A(new_n697), .B1(new_n706), .B2(new_n670), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT27), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1996), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n657), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n657), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n696), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT95), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n657), .A2(G6), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n573), .B2(new_n657), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G23), .B(G288), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT33), .B(G1976), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n657), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n657), .ZN(new_n724));
  MUX2_X1   g299(.A(new_n723), .B(new_n724), .S(KEYINPUT87), .Z(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1971), .Z(new_n726));
  NAND3_X1  g301(.A1(new_n719), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT34), .Z(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G24), .ZN(new_n729));
  XNOR2_X1  g304(.A(G290), .B(KEYINPUT86), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1986), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n703), .A2(G131), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT84), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n484), .A2(G119), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n473), .A2(G107), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT85), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n739), .B(new_n741), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n728), .A2(new_n732), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n670), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n670), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2090), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  NAND2_X1  g325(.A1(G299), .A2(G16), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n657), .A2(KEYINPUT23), .A3(G20), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT23), .ZN(new_n753));
  INV_X1    g328(.A(G20), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G16), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n751), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1956), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n670), .A2(G26), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n474), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G128), .B2(new_n484), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(new_n670), .ZN(new_n764));
  MUX2_X1   g339(.A(new_n758), .B(new_n764), .S(KEYINPUT28), .Z(new_n765));
  AOI22_X1  g340(.A1(new_n748), .A2(G2090), .B1(new_n765), .B2(G2067), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n750), .A2(new_n757), .A3(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n715), .A2(new_n745), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n765), .A2(G2067), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n657), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n586), .B2(new_n657), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n545), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1341), .Z(new_n776));
  NAND4_X1  g351(.A1(new_n768), .A2(new_n769), .A3(new_n773), .A4(new_n776), .ZN(G150));
  INV_X1    g352(.A(G150), .ZN(G311));
  AOI22_X1  g353(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n510), .ZN(new_n780));
  INV_X1    g355(.A(G93), .ZN(new_n781));
  INV_X1    g356(.A(G55), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n513), .A2(new_n781), .B1(new_n515), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G860), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT37), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n585), .A2(new_n591), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n785), .B1(new_n542), .B2(new_n540), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n545), .A2(new_n785), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n790), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n787), .B1(new_n795), .B2(G860), .ZN(G145));
  XNOR2_X1  g371(.A(new_n602), .B(new_n476), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G162), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n484), .A2(G130), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n703), .A2(G142), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n473), .A2(G118), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n738), .B(new_n804), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(new_n606), .ZN(new_n807));
  MUX2_X1   g382(.A(new_n705), .B(new_n706), .S(new_n686), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n763), .B(KEYINPUT99), .ZN(new_n809));
  INV_X1    g384(.A(new_n492), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n499), .A2(KEYINPUT98), .A3(new_n501), .ZN(new_n811));
  AOI21_X1  g386(.A(KEYINPUT98), .B1(new_n499), .B2(new_n501), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n809), .B(new_n813), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n808), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n807), .A2(KEYINPUT102), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n807), .B(new_n815), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n798), .B(new_n816), .C1(new_n817), .C2(KEYINPUT102), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n798), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT103), .B(G37), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g397(.A(new_n585), .B(G299), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(KEYINPUT41), .B2(new_n823), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n593), .B(new_n794), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n823), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n573), .B(G303), .ZN(new_n830));
  XNOR2_X1  g405(.A(G288), .B(G290), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT42), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n829), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G868), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G868), .B2(new_n784), .ZN(G295));
  OAI21_X1  g411(.A(new_n835), .B1(G868), .B2(new_n784), .ZN(G331));
  INV_X1    g412(.A(KEYINPUT109), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n839));
  XNOR2_X1  g414(.A(G286), .B(G171), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n794), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT105), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n794), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n823), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT106), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n841), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n823), .A2(new_n824), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(KEYINPUT108), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n823), .A2(KEYINPUT41), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n832), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n844), .A2(new_n826), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n848), .A2(new_n823), .ZN(new_n856));
  INV_X1    g431(.A(new_n832), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n820), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n856), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(KEYINPUT107), .A3(new_n832), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n832), .A2(KEYINPUT107), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n855), .A2(new_n856), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n860), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n839), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n859), .A2(KEYINPUT43), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(KEYINPUT43), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT44), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n838), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n869), .A2(new_n873), .A3(KEYINPUT109), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(G397));
  INV_X1    g452(.A(G1384), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n813), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(G160), .A2(G40), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n884), .A2(new_n885), .A3(G1996), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n763), .B(G2067), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n883), .B1(new_n705), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n884), .B2(G1996), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT47), .Z(new_n892));
  NOR2_X1   g467(.A1(G290), .A2(G1986), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT111), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n883), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT48), .Z(new_n896));
  INV_X1    g471(.A(new_n706), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n887), .B1(new_n897), .B2(G1996), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G1996), .B2(new_n705), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n738), .A2(new_n741), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n738), .A2(new_n741), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n896), .B1(new_n883), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(KEYINPUT126), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n901), .A2(KEYINPUT126), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G2067), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n763), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n884), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n892), .A2(new_n904), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n912));
  INV_X1    g487(.A(new_n882), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n813), .A2(new_n878), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G8), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G1976), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(G288), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT114), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n917), .B(new_n922), .C1(new_n918), .C2(G288), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n921), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n573), .A2(new_n653), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n541), .A2(G86), .ZN(new_n926));
  OAI21_X1  g501(.A(G1981), .B1(new_n572), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT49), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n929), .A2(new_n917), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n499), .A2(new_n501), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT98), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n499), .A2(KEYINPUT98), .A3(new_n501), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G1384), .B1(new_n936), .B2(new_n810), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n882), .B1(new_n937), .B2(KEYINPUT45), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n932), .B2(new_n810), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n880), .ZN(new_n941));
  AOI21_X1  g516(.A(G1971), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G2090), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n813), .A2(new_n944), .A3(new_n878), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n913), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n939), .B2(new_n944), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT112), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n942), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(new_n916), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n954));
  NAND3_X1  g529(.A1(G303), .A2(G8), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n956));
  OAI22_X1  g531(.A1(G166), .A2(new_n916), .B1(KEYINPUT113), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n940), .A2(KEYINPUT50), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n882), .B(new_n961), .C1(KEYINPUT50), .C2(new_n879), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n942), .B1(new_n943), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n963), .B2(new_n916), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n931), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n913), .C1(new_n937), .C2(KEYINPUT45), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n940), .A2(new_n880), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n913), .A2(KEYINPUT45), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n914), .A2(KEYINPUT117), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n661), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n946), .A2(G2084), .A3(new_n950), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n916), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G168), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n912), .B1(new_n965), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n931), .A2(KEYINPUT115), .ZN(new_n978));
  INV_X1    g553(.A(new_n960), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT63), .B1(new_n953), .B2(new_n959), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n924), .B2(new_n930), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n977), .B1(new_n976), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n978), .A2(new_n979), .A3(new_n983), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n930), .A2(G1976), .A3(G288), .ZN(new_n987));
  INV_X1    g562(.A(new_n925), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n917), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n986), .A2(KEYINPUT116), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT116), .B1(new_n986), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(G168), .A2(new_n916), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n975), .A2(KEYINPUT51), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT121), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n973), .C1(new_n661), .C2(new_n971), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT121), .B1(new_n972), .B2(new_n974), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT122), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(G8), .C1(new_n996), .C2(new_n997), .ZN(new_n1001));
  INV_X1    g576(.A(new_n993), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n994), .B1(new_n1003), .B2(KEYINPUT51), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n972), .A2(new_n974), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n995), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n972), .A2(KEYINPUT121), .A3(new_n974), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n938), .A2(new_n941), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(G2078), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT119), .B1(new_n946), .B2(new_n950), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n948), .A2(new_n949), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n913), .A4(new_n945), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1016), .A3(new_n712), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n675), .A2(KEYINPUT53), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1012), .B(new_n1017), .C1(new_n971), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G171), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT62), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1008), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n916), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n993), .B1(new_n1025), .B2(new_n1000), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1026), .B2(new_n999), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1022), .B(new_n1023), .C1(new_n1027), .C2(new_n994), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1009), .A2(new_n1021), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1023), .B1(new_n1027), .B2(new_n994), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT56), .B(G2072), .Z(new_n1031));
  OAI22_X1  g606(.A1(new_n962), .A2(G1956), .B1(new_n1011), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G299), .B(KEYINPUT57), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1033), .ZN(new_n1035));
  OAI221_X1 g610(.A(new_n1035), .B1(new_n1011), .B2(new_n1031), .C1(new_n962), .C2(G1956), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1034), .A2(new_n1036), .A3(KEYINPUT61), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT61), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1013), .A2(new_n1016), .A3(new_n772), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n915), .A2(new_n908), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT60), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT120), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1040), .A2(new_n1045), .A3(KEYINPUT60), .A4(new_n1041), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n586), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT58), .B(G1341), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1011), .A2(G1996), .B1(new_n915), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n545), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT59), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1044), .A2(new_n586), .A3(new_n1048), .A4(new_n1046), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1039), .A2(new_n1050), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1036), .A2(new_n586), .A3(new_n1042), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1034), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1017), .A2(KEYINPUT123), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n938), .A2(KEYINPUT53), .A3(new_n675), .A4(new_n881), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1013), .A2(new_n1016), .A3(new_n1061), .A4(new_n712), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1059), .A2(new_n1012), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G171), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(KEYINPUT54), .C1(G171), .C2(new_n1019), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1020), .B1(new_n1063), .B2(G171), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1030), .A2(new_n1058), .A3(new_n1065), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1029), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n965), .B(KEYINPUT125), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n992), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n903), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n894), .B1(G1986), .B2(G290), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n884), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n911), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT127), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT127), .B(new_n911), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g657(.A(new_n821), .ZN(new_n1084));
  NOR3_X1   g658(.A1(new_n1084), .A2(G401), .A3(G227), .ZN(new_n1085));
  INV_X1    g659(.A(G229), .ZN(new_n1086));
  NAND2_X1  g660(.A1(new_n871), .A2(new_n872), .ZN(new_n1087));
  NAND4_X1  g661(.A1(new_n1085), .A2(G319), .A3(new_n1086), .A4(new_n1087), .ZN(G225));
  INV_X1    g662(.A(G225), .ZN(G308));
endmodule


