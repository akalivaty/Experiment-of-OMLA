

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XNOR2_X1 U323 ( .A(n480), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U324 ( .A(n455), .B(n454), .ZN(n504) );
  XOR2_X1 U325 ( .A(n368), .B(n367), .Z(n519) );
  XNOR2_X1 U326 ( .A(n340), .B(G43GAT), .ZN(n341) );
  XNOR2_X1 U327 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  INV_X1 U328 ( .A(KEYINPUT11), .ZN(n303) );
  XNOR2_X1 U329 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U331 ( .A(n304), .B(n303), .ZN(n305) );
  NOR2_X1 U332 ( .A1(n414), .A2(n413), .ZN(n489) );
  XNOR2_X1 U333 ( .A(n306), .B(n305), .ZN(n311) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n481) );
  XOR2_X1 U335 ( .A(n452), .B(n451), .Z(n562) );
  XNOR2_X1 U336 ( .A(n369), .B(n347), .ZN(n532) );
  XNOR2_X1 U337 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U338 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U339 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n459), .B(n458), .ZN(G1330GAT) );
  INV_X1 U341 ( .A(KEYINPUT77), .ZN(n312) );
  INV_X1 U342 ( .A(G85GAT), .ZN(n291) );
  NAND2_X1 U343 ( .A1(G92GAT), .A2(n291), .ZN(n294) );
  INV_X1 U344 ( .A(G92GAT), .ZN(n292) );
  NAND2_X1 U345 ( .A1(n292), .A2(G85GAT), .ZN(n293) );
  NAND2_X1 U346 ( .A1(n294), .A2(n293), .ZN(n296) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n432) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(n432), .ZN(n302) );
  XNOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n297), .B(G218GAT), .ZN(n374) );
  XNOR2_X1 U352 ( .A(KEYINPUT9), .B(KEYINPUT76), .ZN(n299) );
  AND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U355 ( .A(n374), .B(n300), .Z(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G162GAT), .Z(n386) );
  XNOR2_X1 U358 ( .A(n386), .B(KEYINPUT10), .ZN(n304) );
  XOR2_X1 U359 ( .A(KEYINPUT67), .B(KEYINPUT7), .Z(n308) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(KEYINPUT8), .B(n309), .Z(n448) );
  INV_X1 U363 ( .A(n448), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n560) );
  XNOR2_X1 U365 ( .A(n312), .B(n560), .ZN(n485) );
  XNOR2_X1 U366 ( .A(KEYINPUT36), .B(n485), .ZN(n586) );
  XOR2_X1 U367 ( .A(G211GAT), .B(G78GAT), .Z(n314) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G22GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U370 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n316) );
  XNOR2_X1 U371 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n328) );
  XOR2_X1 U374 ( .A(G8GAT), .B(G183GAT), .Z(n377) );
  XOR2_X1 U375 ( .A(G57GAT), .B(KEYINPUT13), .Z(n418) );
  XOR2_X1 U376 ( .A(n377), .B(n418), .Z(n320) );
  XNOR2_X1 U377 ( .A(G71GAT), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U379 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n322) );
  NAND2_X1 U380 ( .A1(G231GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U382 ( .A(n324), .B(n323), .Z(n326) );
  XOR2_X1 U383 ( .A(G15GAT), .B(G127GAT), .Z(n334) );
  XNOR2_X1 U384 ( .A(n334), .B(KEYINPUT15), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n569) );
  XOR2_X1 U387 ( .A(KEYINPUT84), .B(KEYINPUT18), .Z(n330) );
  XNOR2_X1 U388 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(n331), .ZN(n369) );
  XOR2_X1 U391 ( .A(G183GAT), .B(KEYINPUT83), .Z(n333) );
  XNOR2_X1 U392 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n346) );
  XOR2_X1 U394 ( .A(G99GAT), .B(G190GAT), .Z(n336) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XNOR2_X1 U396 ( .A(n429), .B(n334), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U398 ( .A(n337), .B(KEYINPUT86), .Z(n344) );
  XOR2_X1 U399 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n339) );
  XNOR2_X1 U400 ( .A(G113GAT), .B(G134GAT), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n364) );
  XOR2_X1 U402 ( .A(G176GAT), .B(n364), .Z(n342) );
  NAND2_X1 U403 ( .A1(G227GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U405 ( .A(n346), .B(n345), .Z(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n349) );
  XNOR2_X1 U407 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n368) );
  XOR2_X1 U409 ( .A(G148GAT), .B(G127GAT), .Z(n351) );
  XNOR2_X1 U410 ( .A(G29GAT), .B(G120GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U412 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n353) );
  XNOR2_X1 U413 ( .A(G1GAT), .B(G141GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n362) );
  XOR2_X1 U416 ( .A(G155GAT), .B(KEYINPUT2), .Z(n357) );
  XNOR2_X1 U417 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n398) );
  XOR2_X1 U419 ( .A(G85GAT), .B(G162GAT), .Z(n359) );
  NAND2_X1 U420 ( .A1(G225GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n398), .B(n360), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U424 ( .A(n363), .B(G57GAT), .Z(n366) );
  XNOR2_X1 U425 ( .A(n364), .B(KEYINPUT1), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n367) );
  INV_X1 U427 ( .A(n369), .ZN(n373) );
  XOR2_X1 U428 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n371) );
  XNOR2_X1 U429 ( .A(G204GAT), .B(G92GAT), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n384) );
  XOR2_X1 U432 ( .A(n374), .B(KEYINPUT94), .Z(n376) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U435 ( .A(n378), .B(n377), .Z(n382) );
  XOR2_X1 U436 ( .A(G211GAT), .B(KEYINPUT21), .Z(n380) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n385) );
  XOR2_X1 U439 ( .A(G176GAT), .B(G64GAT), .Z(n419) );
  XNOR2_X1 U440 ( .A(n385), .B(n419), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n472) );
  INV_X1 U443 ( .A(n472), .ZN(n521) );
  XNOR2_X1 U444 ( .A(n521), .B(KEYINPUT27), .ZN(n408) );
  NAND2_X1 U445 ( .A1(n519), .A2(n408), .ZN(n530) );
  NOR2_X1 U446 ( .A1(n532), .A2(n530), .ZN(n401) );
  XOR2_X1 U447 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U448 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U450 ( .A(n389), .B(G106GAT), .Z(n391) );
  XOR2_X1 U451 ( .A(G141GAT), .B(G22GAT), .Z(n441) );
  XNOR2_X1 U452 ( .A(n441), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n393) );
  XNOR2_X1 U455 ( .A(KEYINPUT89), .B(KEYINPUT22), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U457 ( .A(n395), .B(n394), .Z(n400) );
  XOR2_X1 U458 ( .A(G78GAT), .B(G148GAT), .Z(n397) );
  XNOR2_X1 U459 ( .A(KEYINPUT70), .B(G204GAT), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n433) );
  XNOR2_X1 U461 ( .A(n398), .B(n433), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n477) );
  XNOR2_X1 U463 ( .A(n477), .B(KEYINPUT28), .ZN(n497) );
  NAND2_X1 U464 ( .A1(n401), .A2(n497), .ZN(n402) );
  XOR2_X1 U465 ( .A(KEYINPUT96), .B(n402), .Z(n414) );
  AND2_X1 U466 ( .A1(n521), .A2(n532), .ZN(n403) );
  XNOR2_X1 U467 ( .A(KEYINPUT99), .B(n403), .ZN(n404) );
  NAND2_X1 U468 ( .A1(n404), .A2(n477), .ZN(n405) );
  XNOR2_X1 U469 ( .A(KEYINPUT25), .B(n405), .ZN(n411) );
  XNOR2_X1 U470 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n407) );
  NOR2_X1 U471 ( .A1(n532), .A2(n477), .ZN(n406) );
  XOR2_X1 U472 ( .A(n407), .B(n406), .Z(n573) );
  AND2_X1 U473 ( .A1(n573), .A2(n408), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n409), .B(KEYINPUT98), .ZN(n410) );
  NOR2_X1 U475 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U476 ( .A1(n519), .A2(n412), .ZN(n413) );
  NOR2_X1 U477 ( .A1(n569), .A2(n489), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n415), .B(KEYINPUT101), .ZN(n416) );
  NOR2_X1 U479 ( .A1(n586), .A2(n416), .ZN(n417) );
  XNOR2_X1 U480 ( .A(KEYINPUT37), .B(n417), .ZN(n518) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n421) );
  AND2_X1 U482 ( .A1(G230GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U484 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n423) );
  XNOR2_X1 U485 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n431) );
  XOR2_X1 U488 ( .A(KEYINPUT69), .B(KEYINPUT33), .Z(n427) );
  XNOR2_X1 U489 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U493 ( .A(n433), .B(n432), .Z(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n579) );
  XOR2_X1 U495 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n437) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(G8GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n452) );
  XOR2_X1 U498 ( .A(G197GAT), .B(G15GAT), .Z(n439) );
  XNOR2_X1 U499 ( .A(G36GAT), .B(G50GAT), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U501 ( .A(n440), .B(G113GAT), .Z(n443) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n445) );
  NAND2_X1 U505 ( .A1(G229GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(n447), .B(n446), .Z(n450) );
  XNOR2_X1 U508 ( .A(n448), .B(KEYINPUT65), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U510 ( .A1(n579), .A2(n562), .ZN(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT75), .B(n453), .Z(n490) );
  NOR2_X1 U512 ( .A1(n518), .A2(n490), .ZN(n455) );
  XNOR2_X1 U513 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n454) );
  NAND2_X1 U514 ( .A1(n504), .A2(n532), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n457) );
  XNOR2_X1 U516 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(n579), .ZN(n564) );
  NAND2_X1 U520 ( .A1(n562), .A2(n564), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n569), .A2(n463), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n560), .A2(n464), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT47), .ZN(n470) );
  INV_X1 U525 ( .A(n569), .ZN(n582) );
  NOR2_X1 U526 ( .A1(n586), .A2(n582), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n466), .B(KEYINPUT45), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n467), .A2(n579), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n468), .A2(n562), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT48), .ZN(n531) );
  NOR2_X1 U532 ( .A1(n472), .A2(n531), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n519), .A2(n476), .ZN(n574) );
  NAND2_X1 U535 ( .A1(n477), .A2(n574), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT55), .B(n478), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n532), .ZN(n480) );
  INV_X1 U538 ( .A(n485), .ZN(n544) );
  NAND2_X1 U539 ( .A1(n570), .A2(n544), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n482) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n492) );
  XOR2_X1 U542 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n487) );
  NAND2_X1 U543 ( .A1(n569), .A2(n485), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(n488) );
  OR2_X1 U545 ( .A1(n489), .A2(n488), .ZN(n506) );
  NOR2_X1 U546 ( .A1(n490), .A2(n506), .ZN(n498) );
  NAND2_X1 U547 ( .A1(n519), .A2(n498), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n521), .A2(n498), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n495) );
  NAND2_X1 U552 ( .A1(n498), .A2(n532), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n496), .ZN(G1326GAT) );
  INV_X1 U555 ( .A(n497), .ZN(n535) );
  NAND2_X1 U556 ( .A1(n498), .A2(n535), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U558 ( .A1(n504), .A2(n519), .ZN(n502) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n521), .A2(n504), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n535), .A2(n504), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  INV_X1 U567 ( .A(n562), .ZN(n575) );
  NAND2_X1 U568 ( .A1(n575), .A2(n564), .ZN(n517) );
  NOR2_X1 U569 ( .A1(n517), .A2(n506), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n519), .A2(n512), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n521), .A2(n512), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n532), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n535), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT108), .Z(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n519), .A2(n526), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U586 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n532), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(KEYINPUT110), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n535), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT115), .Z(n538) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n532), .A2(n548), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT113), .B(n533), .Z(n534) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(KEYINPUT114), .B(n536), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n562), .A2(n545), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U604 ( .A1(n545), .A2(n564), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n545), .A2(n569), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n573), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n575), .A2(n559), .ZN(n549) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  INV_X1 U616 ( .A(n564), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n550), .A2(n559), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT52), .B(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n582), .A2(n559), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n570), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n566) );
  NAND2_X1 U633 ( .A1(n570), .A2(n564), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  XOR2_X1 U636 ( .A(G183GAT), .B(KEYINPUT125), .Z(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n585) );
  NOR2_X1 U640 ( .A1(n575), .A2(n585), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

