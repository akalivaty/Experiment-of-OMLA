//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n455), .A2(new_n449), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI211_X1 g051(.A(G137), .B(new_n466), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n477), .ZN(new_n479));
  INV_X1    g054(.A(G101), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n470), .B2(new_n471), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n467), .B1(new_n478), .B2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n464), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n464), .A2(new_n466), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n490), .B2(G136), .ZN(G162));
  NAND3_X1  g066(.A1(new_n464), .A2(G138), .A3(new_n466), .ZN(new_n492));
  OAI21_X1  g067(.A(G126), .B1(new_n475), .B2(new_n476), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n466), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n466), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT73), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G50), .A2(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT72), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n521), .B1(new_n516), .B2(new_n519), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n526), .A2(new_n527), .A3(G50), .A4(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n506), .A2(new_n508), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT74), .B(G88), .Z(new_n532));
  AOI22_X1  g107(.A1(new_n525), .A2(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n514), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n526), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT76), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(new_n538), .A3(G543), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n537), .A2(G51), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n542), .B1(new_n509), .B2(new_n543), .C1(new_n530), .C2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n540), .A2(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n509), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n531), .A2(G90), .B1(G651), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n537), .A2(new_n539), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n509), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  INV_X1    g135(.A(new_n551), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n560), .B1(new_n561), .B2(G43), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  AND2_X1   g142(.A1(G53), .A2(G543), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n520), .A2(new_n522), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n570), .B1(new_n526), .B2(new_n568), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n530), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n506), .A2(new_n508), .A3(G65), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n579), .A2(G78), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT79), .B1(new_n576), .B2(new_n581), .ZN(new_n584));
  NOR3_X1   g159(.A1(new_n583), .A2(new_n584), .A3(new_n515), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT80), .B1(new_n575), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n526), .A2(new_n529), .A3(G91), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n526), .A2(new_n570), .A3(new_n568), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n569), .A2(new_n571), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n576), .A2(new_n581), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n594), .A2(G651), .A3(new_n582), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n586), .A2(new_n596), .ZN(G299));
  INV_X1    g172(.A(G168), .ZN(G286));
  NAND2_X1  g173(.A1(new_n531), .A2(G87), .ZN(new_n599));
  INV_X1    g174(.A(new_n536), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G49), .ZN(new_n601));
  OAI211_X1 g176(.A(KEYINPUT81), .B(G651), .C1(new_n529), .C2(G74), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  AOI21_X1  g178(.A(G74), .B1(new_n506), .B2(new_n508), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n515), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n599), .A2(new_n601), .A3(new_n606), .ZN(G288));
  INV_X1    g182(.A(G48), .ZN(new_n608));
  INV_X1    g183(.A(G86), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n608), .A2(new_n536), .B1(new_n530), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n612));
  NAND2_X1  g187(.A1(G73), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G61), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n509), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n612), .B1(new_n615), .B2(G651), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n615), .A2(new_n612), .A3(G651), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(G305));
  NAND2_X1  g193(.A1(G72), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G60), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n509), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n531), .A2(G85), .B1(G651), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n537), .A2(G47), .A3(new_n539), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n530), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT10), .A4(G92), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n537), .A2(G54), .A3(new_n539), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(new_n515), .ZN(new_n633));
  AND3_X1   g208(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n625), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n625), .B1(new_n634), .B2(G868), .ZN(G321));
  NAND2_X1  g211(.A1(new_n589), .A2(new_n588), .ZN(new_n637));
  INV_X1    g212(.A(new_n587), .ZN(new_n638));
  AND4_X1   g213(.A1(new_n591), .A2(new_n595), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n591), .B1(new_n590), .B2(new_n595), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G868), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(G168), .A2(G868), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G297));
  XOR2_X1   g221(.A(new_n645), .B(KEYINPUT83), .Z(G280));
  INV_X1    g222(.A(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n634), .B1(new_n648), .B2(G860), .ZN(G148));
  NAND2_X1  g224(.A1(new_n634), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G868), .ZN(new_n651));
  INV_X1    g226(.A(G43), .ZN(new_n652));
  OAI221_X1 g227(.A(new_n558), .B1(new_n559), .B2(new_n530), .C1(new_n551), .C2(new_n652), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n651), .A2(KEYINPUT84), .B1(new_n642), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(KEYINPUT84), .B2(new_n651), .ZN(G323));
  XNOR2_X1  g230(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g231(.A(new_n484), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G123), .ZN(new_n658));
  NOR2_X1   g233(.A1(G99), .A2(G2105), .ZN(new_n659));
  OAI21_X1  g234(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n490), .A2(KEYINPUT85), .A3(G135), .ZN(new_n661));
  AOI21_X1  g236(.A(KEYINPUT85), .B1(new_n490), .B2(G135), .ZN(new_n662));
  OAI221_X1 g237(.A(new_n658), .B1(new_n659), .B2(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n472), .A2(new_n464), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT12), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT13), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n669), .ZN(G156));
  XNOR2_X1  g245(.A(G2427), .B(G2438), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2430), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(KEYINPUT14), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2451), .B(G2454), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT16), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n677), .A2(new_n679), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(new_n679), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1341), .B(G1348), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n690), .A3(new_n686), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  OAI211_X1 g269(.A(G14), .B(new_n689), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g271(.A(G2072), .B(G2078), .Z(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT17), .Z(new_n698));
  XOR2_X1   g273(.A(G2084), .B(G2090), .Z(new_n699));
  XNOR2_X1  g274(.A(G2067), .B(G2678), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(new_n697), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n700), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n697), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT18), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(new_n664), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G2100), .ZN(G227));
  XNOR2_X1  g285(.A(G1971), .B(G1976), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT19), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(G1956), .B(G2474), .Z(new_n714));
  XOR2_X1   g289(.A(G1961), .B(G1966), .Z(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n714), .A2(new_n715), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n721), .B(new_n720), .S(new_n713), .Z(new_n722));
  NOR2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1986), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(G1991), .B(G1996), .ZN(new_n727));
  INV_X1    g302(.A(G1981), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n726), .B(new_n729), .ZN(G229));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NOR2_X1   g306(.A1(G168), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n731), .B2(G21), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(G5), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G171), .B2(new_n731), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G1961), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G1961), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n733), .A2(new_n734), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n735), .A2(new_n738), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G34), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G160), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2078), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n663), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(G32), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT26), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n472), .A2(G105), .ZN(new_n757));
  INV_X1    g332(.A(G129), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n484), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G141), .B2(new_n490), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n752), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n752), .A2(G33), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  AOI22_X1  g342(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n466), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n490), .B2(G139), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(new_n752), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G2072), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n761), .A2(new_n763), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n753), .A2(new_n764), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(new_n749), .B2(G2078), .C1(new_n771), .C2(G2072), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n741), .A2(new_n751), .A3(new_n774), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n731), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n562), .B2(new_n731), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1341), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n752), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  INV_X1    g364(.A(G128), .ZN(new_n790));
  NOR2_X1   g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n484), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n490), .B2(G140), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(new_n752), .ZN(new_n795));
  INV_X1    g370(.A(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n731), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n634), .B2(new_n731), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT91), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n798), .A2(KEYINPUT91), .A3(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n752), .A2(G35), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G162), .B2(new_n752), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2090), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n731), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n641), .B2(new_n731), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1956), .Z(new_n812));
  AND4_X1   g387(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n784), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n784), .A2(KEYINPUT95), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n731), .A2(G22), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G166), .B2(new_n731), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(G1971), .ZN(new_n821));
  NOR2_X1   g396(.A1(G6), .A2(G16), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n617), .A2(new_n616), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n610), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n824), .B2(G16), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT32), .B(G1981), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n731), .A2(G23), .ZN(new_n828));
  INV_X1    g403(.A(G288), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n731), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT33), .B(G1976), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT90), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n820), .A2(G1971), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n821), .A2(new_n827), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n657), .A2(G119), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT89), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n490), .A2(G131), .ZN(new_n839));
  NOR2_X1   g414(.A1(G95), .A2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  MUX2_X1   g417(.A(G25), .B(new_n842), .S(G29), .Z(new_n843));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G1991), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G290), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G16), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G16), .B2(G24), .ZN(new_n849));
  INV_X1    g424(.A(G1986), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n846), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n836), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n818), .A2(new_n856), .ZN(G150));
  INV_X1    g432(.A(G150), .ZN(G311));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n509), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n515), .B1(new_n861), .B2(KEYINPUT96), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(KEYINPUT96), .B2(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n537), .A2(G55), .A3(new_n539), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n531), .A2(G93), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND4_X1  g443(.A1(new_n562), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n653), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n634), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT97), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n878));
  AOI21_X1  g453(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n868), .B1(new_n880), .B2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(new_n794), .B(new_n502), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n770), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n842), .B(new_n667), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n490), .A2(G142), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n657), .A2(G130), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n891), .A2(new_n466), .A3(G118), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n466), .B2(G118), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n889), .B(new_n890), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n760), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n888), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n663), .B(G160), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G162), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n888), .B(new_n897), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n901), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT40), .Z(G395));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n586), .A2(new_n596), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  AOI211_X1 g490(.A(new_n915), .B(new_n911), .C1(new_n586), .C2(new_n596), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT101), .B1(G299), .B2(new_n634), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n914), .B(KEYINPUT102), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n871), .B(new_n650), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(new_n824), .ZN(new_n929));
  NAND3_X1  g504(.A1(G305), .A2(new_n533), .A3(new_n514), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n847), .A2(G288), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n829), .A2(G290), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n929), .A2(new_n930), .A3(new_n932), .A4(new_n933), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n935), .A2(KEYINPUT103), .A3(new_n937), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT103), .B1(new_n935), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n941), .B2(new_n936), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n909), .B1(new_n928), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n927), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n924), .B2(new_n922), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n946), .B2(new_n942), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n928), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(KEYINPUT104), .A3(new_n942), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n944), .A2(new_n947), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(G868), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n866), .A2(new_n642), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(G295));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n952), .B2(new_n953), .ZN(new_n956));
  INV_X1    g531(.A(new_n953), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT106), .B(new_n957), .C1(new_n951), .C2(G868), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(G331));
  NAND2_X1  g534(.A1(G286), .A2(G171), .ZN(new_n960));
  NAND2_X1  g535(.A1(G168), .A2(G301), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n871), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n960), .A2(new_n869), .A3(new_n870), .A4(new_n961), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n913), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n910), .A2(new_n915), .ZN(new_n969));
  NAND3_X1  g544(.A1(G299), .A2(KEYINPUT101), .A3(new_n634), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n971), .B2(KEYINPUT102), .ZN(new_n972));
  INV_X1    g547(.A(new_n921), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n939), .A2(new_n940), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n965), .A2(new_n926), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n906), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n976), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n974), .A2(KEYINPUT107), .A3(new_n976), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n976), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n922), .B2(new_n966), .ZN(new_n987));
  AOI21_X1  g562(.A(G37), .B1(new_n987), .B2(new_n975), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT41), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n926), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n968), .B1(G299), .B2(new_n634), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n966), .B(new_n989), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n926), .B2(new_n990), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT108), .B(new_n976), .C1(new_n994), .C2(new_n965), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n995), .A3(new_n941), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n988), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n985), .B(KEYINPUT44), .C1(new_n984), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(new_n984), .A3(new_n996), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n983), .B2(new_n984), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT109), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n965), .B1(new_n920), .B2(new_n921), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n980), .B1(new_n1003), .B2(new_n986), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n982), .A3(new_n941), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n984), .B1(new_n1005), .B2(new_n988), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n984), .A2(new_n996), .A3(new_n906), .A4(new_n977), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT109), .B(new_n1001), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1002), .B2(new_n1009), .ZN(G397));
  OR2_X1    g585(.A1(new_n465), .A2(new_n466), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT69), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n474), .B1(new_n473), .B2(new_n477), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1011), .B(G40), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  NAND3_X1  g591(.A1(G160), .A2(new_n1016), .A3(G40), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT45), .B1(new_n502), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(G1996), .A3(new_n896), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT111), .Z(new_n1023));
  XNOR2_X1  g598(.A(new_n794), .B(new_n796), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT112), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G1996), .B2(new_n896), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1021), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n842), .B(new_n844), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G290), .B(G1986), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1021), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1033), .B(G1384), .C1(new_n497), .C2(new_n501), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1020), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2078), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1018), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(KEYINPUT125), .A3(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n502), .A2(new_n1019), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1015), .A2(new_n1017), .B1(new_n1043), .B2(KEYINPUT50), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n502), .A2(new_n1045), .A3(new_n1019), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1036), .A2(KEYINPUT53), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1014), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1035), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1041), .A2(new_n1042), .A3(new_n1049), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1039), .A2(new_n1040), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1035), .A2(new_n1018), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(new_n1050), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1055), .A2(G301), .A3(new_n1042), .A4(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1054), .A2(KEYINPUT54), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1041), .A2(new_n1042), .A3(new_n1049), .A4(new_n1057), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G171), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1055), .A2(G301), .A3(new_n1042), .A4(new_n1052), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT54), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1018), .A2(new_n746), .A3(new_n1064), .A4(new_n1046), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1044), .A2(KEYINPUT120), .A3(new_n746), .A4(new_n1046), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1056), .A2(new_n734), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G286), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1067), .A2(new_n1069), .A3(G168), .A4(new_n1068), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(KEYINPUT51), .A3(G8), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1059), .A2(new_n1063), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  AND4_X1   g655(.A1(new_n1080), .A2(new_n1018), .A3(new_n1064), .A4(new_n1046), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1971), .B1(new_n1035), .B2(new_n1018), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1971), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1056), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1044), .A2(new_n1080), .A3(new_n1046), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(KEYINPUT113), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G303), .A2(G8), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1088), .B(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1083), .A2(new_n1087), .A3(G8), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1079), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT115), .A3(new_n1091), .A4(new_n1087), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1043), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1095), .B1(new_n1018), .B2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n599), .A2(new_n601), .A3(new_n606), .A4(G1976), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT116), .ZN(new_n1103));
  INV_X1    g678(.A(G1976), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT52), .B1(G288), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1101), .A2(KEYINPUT117), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(G1981), .B1(new_n823), .B2(new_n610), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n611), .B(new_n728), .C1(new_n616), .C2(new_n617), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT49), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1114), .A2(new_n1101), .B1(new_n1115), .B2(KEYINPUT52), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1046), .B(KEYINPUT119), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1080), .A3(new_n1044), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1085), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1091), .B1(new_n1120), .B2(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1099), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1099), .A2(new_n1122), .A3(KEYINPUT126), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1956), .B1(new_n1118), .B2(new_n1044), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT56), .B(G2072), .Z(new_n1128));
  NOR2_X1   g703(.A1(new_n1056), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n590), .A2(new_n595), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT57), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1047), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1018), .A2(new_n796), .A3(new_n1100), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n911), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1134), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1018), .A2(new_n1100), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1996), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1035), .A2(new_n1144), .A3(new_n1018), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n653), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT123), .B1(new_n1146), .B2(KEYINPUT124), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1137), .A2(new_n911), .A3(new_n1138), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n1150), .B2(new_n1139), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1146), .A2(KEYINPUT123), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1149), .B(new_n1151), .C1(new_n1153), .C2(new_n1147), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1137), .A2(new_n1138), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT61), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n1158));
  NOR4_X1   g733(.A1(new_n1127), .A2(new_n1129), .A3(new_n1158), .A4(new_n1132), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1140), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1078), .A2(new_n1125), .A3(new_n1126), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1077), .A2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1072), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1165), .A2(new_n1071), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1061), .B1(new_n1166), .B2(KEYINPUT62), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1125), .A2(new_n1126), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1099), .A2(new_n1117), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1114), .A2(new_n1101), .ZN(new_n1170));
  NOR2_X1   g745(.A1(G288), .A2(G1976), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT118), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1112), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1101), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1162), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1070), .A2(G8), .A3(G168), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1099), .A2(new_n1176), .A3(new_n1122), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1099), .A2(KEYINPUT121), .A3(new_n1122), .A4(new_n1176), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1117), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1097), .A2(new_n1087), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1091), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1181), .B(KEYINPUT122), .C1(new_n1182), .C2(new_n1091), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1099), .A2(KEYINPUT63), .A3(new_n1176), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1179), .A2(new_n1180), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1032), .B1(new_n1175), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1028), .B1(new_n1025), .B2(new_n760), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT46), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1021), .A2(new_n1144), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1194), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT47), .Z(new_n1196));
  NAND3_X1  g771(.A1(new_n1021), .A2(new_n850), .A3(new_n847), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT48), .Z(new_n1198));
  NOR2_X1   g773(.A1(new_n1030), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n842), .A2(new_n845), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1027), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n794), .A2(new_n796), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1028), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1196), .A2(new_n1199), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1190), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g780(.A1(G227), .A2(new_n462), .ZN(new_n1207));
  NOR2_X1   g781(.A1(G229), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1208), .A2(new_n695), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n1208), .A2(new_n695), .A3(KEYINPUT127), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n907), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n1213), .A2(new_n1000), .ZN(G308));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1000), .ZN(G225));
endmodule


