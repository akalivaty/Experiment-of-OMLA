

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  INV_X1 U326 ( .A(n588), .ZN(n472) );
  XNOR2_X1 U327 ( .A(n379), .B(n378), .ZN(n389) );
  XNOR2_X1 U328 ( .A(n459), .B(KEYINPUT111), .ZN(n460) );
  INV_X1 U329 ( .A(n540), .ZN(n530) );
  INV_X1 U330 ( .A(n538), .ZN(n527) );
  NAND2_X1 U331 ( .A1(n557), .A2(n465), .ZN(n544) );
  XNOR2_X2 U332 ( .A(n403), .B(n402), .ZN(n485) );
  XOR2_X1 U333 ( .A(KEYINPUT37), .B(n460), .Z(n493) );
  XNOR2_X2 U334 ( .A(n494), .B(KEYINPUT38), .ZN(n523) );
  XNOR2_X1 U335 ( .A(n480), .B(KEYINPUT48), .ZN(n558) );
  XNOR2_X1 U336 ( .A(n348), .B(n347), .ZN(n349) );
  NAND2_X1 U337 ( .A1(n571), .A2(n570), .ZN(n294) );
  INV_X1 U338 ( .A(KEYINPUT74), .ZN(n302) );
  XNOR2_X1 U339 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U340 ( .A(n388), .B(n304), .ZN(n307) );
  INV_X1 U341 ( .A(KEYINPUT106), .ZN(n419) );
  XNOR2_X1 U342 ( .A(n407), .B(KEYINPUT104), .ZN(n408) );
  XNOR2_X1 U343 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U344 ( .A(n409), .B(n408), .ZN(n578) );
  XOR2_X1 U345 ( .A(n312), .B(n311), .Z(n585) );
  NOR2_X1 U346 ( .A1(n352), .A2(n572), .ZN(n576) );
  XNOR2_X1 U347 ( .A(n462), .B(n461), .ZN(n541) );
  XNOR2_X1 U348 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U349 ( .A(KEYINPUT44), .B(G106GAT), .ZN(n466) );
  XNOR2_X1 U350 ( .A(KEYINPUT118), .B(G99GAT), .ZN(n463) );
  XNOR2_X1 U351 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n464), .B(n463), .ZN(G1338GAT) );
  INV_X1 U353 ( .A(KEYINPUT116), .ZN(n462) );
  XOR2_X1 U354 ( .A(G92GAT), .B(G64GAT), .Z(n296) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U356 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U357 ( .A(KEYINPUT76), .B(n297), .Z(n383) );
  XOR2_X1 U358 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n299) );
  XNOR2_X1 U359 ( .A(KEYINPUT33), .B(KEYINPUT77), .ZN(n298) );
  XNOR2_X1 U360 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n383), .B(n300), .ZN(n312) );
  XNOR2_X1 U362 ( .A(G148GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n301), .B(G78GAT), .ZN(n388) );
  NAND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n303) );
  XOR2_X1 U365 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n306) );
  XNOR2_X1 U366 ( .A(G71GAT), .B(G57GAT), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n445) );
  XOR2_X1 U368 ( .A(n307), .B(n445), .Z(n310) );
  XOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .Z(n308) );
  XOR2_X1 U370 ( .A(KEYINPUT75), .B(n308), .Z(n421) );
  XNOR2_X1 U371 ( .A(G120GAT), .B(n421), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U373 ( .A(n585), .B(KEYINPUT41), .Z(n570) );
  XOR2_X1 U374 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U375 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n326) );
  XOR2_X1 U377 ( .A(G141GAT), .B(G1GAT), .Z(n316) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G50GAT), .ZN(n315) );
  XNOR2_X1 U379 ( .A(n316), .B(n315), .ZN(n324) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n318) );
  XNOR2_X1 U381 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U383 ( .A(G8GAT), .B(G197GAT), .Z(n320) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(G113GAT), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U386 ( .A(n322), .B(n321), .Z(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n332) );
  XOR2_X1 U389 ( .A(G29GAT), .B(G43GAT), .Z(n328) );
  XNOR2_X1 U390 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n422) );
  XOR2_X1 U392 ( .A(n422), .B(G22GAT), .Z(n330) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U395 ( .A(n332), .B(n331), .Z(n491) );
  AND2_X1 U396 ( .A1(n570), .A2(n491), .ZN(n526) );
  XOR2_X1 U397 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n334) );
  XNOR2_X1 U398 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U400 ( .A(G169GAT), .B(n335), .Z(n377) );
  XOR2_X1 U401 ( .A(G15GAT), .B(G127GAT), .Z(n453) );
  XOR2_X1 U402 ( .A(G190GAT), .B(G134GAT), .Z(n337) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(G99GAT), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U405 ( .A(n453), .B(n338), .Z(n340) );
  NAND2_X1 U406 ( .A1(G227GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n340), .B(n339), .ZN(n342) );
  INV_X1 U408 ( .A(KEYINPUT20), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n350) );
  XOR2_X1 U410 ( .A(G120GAT), .B(KEYINPUT86), .Z(n344) );
  XNOR2_X1 U411 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n359), .B(KEYINPUT89), .ZN(n348) );
  XOR2_X1 U414 ( .A(KEYINPUT87), .B(G71GAT), .Z(n346) );
  XNOR2_X1 U415 ( .A(G176GAT), .B(G183GAT), .ZN(n345) );
  XOR2_X1 U416 ( .A(n346), .B(n345), .Z(n347) );
  XOR2_X1 U417 ( .A(n377), .B(n351), .Z(n352) );
  XOR2_X1 U418 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n354) );
  XNOR2_X1 U419 ( .A(G1GAT), .B(G127GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U421 ( .A(G155GAT), .B(G162GAT), .Z(n356) );
  XNOR2_X1 U422 ( .A(G29GAT), .B(G85GAT), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n376) );
  XOR2_X1 U425 ( .A(G134GAT), .B(KEYINPUT79), .Z(n434) );
  XOR2_X1 U426 ( .A(n434), .B(n359), .Z(n361) );
  NAND2_X1 U427 ( .A1(G225GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U429 ( .A(n362), .B(G57GAT), .Z(n366) );
  XOR2_X1 U430 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n364) );
  XNOR2_X1 U431 ( .A(G141GAT), .B(KEYINPUT91), .ZN(n363) );
  XNOR2_X1 U432 ( .A(n364), .B(n363), .ZN(n399) );
  XNOR2_X1 U433 ( .A(n399), .B(G148GAT), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U435 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n368) );
  XNOR2_X1 U436 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n367) );
  XNOR2_X1 U437 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U438 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n370) );
  XNOR2_X1 U439 ( .A(KEYINPUT6), .B(KEYINPUT98), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U441 ( .A(n372), .B(n371), .Z(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U443 ( .A(n376), .B(n375), .Z(n538) );
  INV_X1 U444 ( .A(n377), .ZN(n387) );
  XOR2_X1 U445 ( .A(G211GAT), .B(KEYINPUT21), .Z(n379) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(G218GAT), .ZN(n378) );
  XOR2_X1 U447 ( .A(KEYINPUT101), .B(n389), .Z(n381) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U450 ( .A(G8GAT), .B(G183GAT), .Z(n441) );
  XOR2_X1 U451 ( .A(n382), .B(n441), .Z(n385) );
  XOR2_X1 U452 ( .A(G36GAT), .B(G190GAT), .Z(n424) );
  XNOR2_X1 U453 ( .A(n383), .B(n424), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U455 ( .A(n387), .B(n386), .Z(n540) );
  XNOR2_X1 U456 ( .A(KEYINPUT27), .B(n530), .ZN(n410) );
  NOR2_X1 U457 ( .A1(n527), .A2(n410), .ZN(n557) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n403) );
  XOR2_X1 U459 ( .A(KEYINPUT94), .B(KEYINPUT22), .Z(n391) );
  XNOR2_X1 U460 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U462 ( .A(G22GAT), .B(G155GAT), .Z(n442) );
  XOR2_X1 U463 ( .A(KEYINPUT90), .B(n442), .Z(n393) );
  XOR2_X1 U464 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U465 ( .A(G204GAT), .B(n423), .ZN(n392) );
  XNOR2_X1 U466 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U467 ( .A(n395), .B(n394), .ZN(n397) );
  AND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U469 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U470 ( .A(KEYINPUT24), .B(n398), .Z(n401) );
  XNOR2_X1 U471 ( .A(n399), .B(KEYINPUT23), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n485), .B(KEYINPUT67), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n404), .B(KEYINPUT28), .ZN(n465) );
  XOR2_X1 U475 ( .A(n544), .B(KEYINPUT102), .Z(n405) );
  NAND2_X1 U476 ( .A1(n352), .A2(n405), .ZN(n406) );
  XNOR2_X1 U477 ( .A(n406), .B(KEYINPUT103), .ZN(n418) );
  AND2_X1 U478 ( .A1(n485), .A2(n352), .ZN(n409) );
  INV_X1 U479 ( .A(KEYINPUT26), .ZN(n407) );
  NOR2_X1 U480 ( .A1(n578), .A2(n410), .ZN(n415) );
  NOR2_X1 U481 ( .A1(n352), .A2(n530), .ZN(n411) );
  NOR2_X1 U482 ( .A1(n485), .A2(n411), .ZN(n412) );
  XNOR2_X1 U483 ( .A(n412), .B(KEYINPUT25), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n413), .B(KEYINPUT105), .ZN(n414) );
  NOR2_X1 U485 ( .A1(n415), .A2(n414), .ZN(n416) );
  NOR2_X1 U486 ( .A1(n538), .A2(n416), .ZN(n417) );
  NOR2_X1 U487 ( .A1(n418), .A2(n417), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n503) );
  XOR2_X1 U489 ( .A(n422), .B(n421), .Z(n438) );
  XOR2_X1 U490 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U491 ( .A1(G232GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U493 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n428) );
  XNOR2_X1 U494 ( .A(G92GAT), .B(G106GAT), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U496 ( .A(n430), .B(n429), .Z(n436) );
  XOR2_X1 U497 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n432) );
  XNOR2_X1 U498 ( .A(G218GAT), .B(KEYINPUT66), .ZN(n431) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U502 ( .A(n438), .B(n437), .Z(n498) );
  INV_X1 U503 ( .A(n498), .ZN(n567) );
  XOR2_X1 U504 ( .A(KEYINPUT36), .B(n567), .Z(n593) );
  XOR2_X1 U505 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n440) );
  XNOR2_X1 U506 ( .A(G211GAT), .B(G78GAT), .ZN(n439) );
  XNOR2_X1 U507 ( .A(n440), .B(n439), .ZN(n457) );
  XOR2_X1 U508 ( .A(n442), .B(n441), .Z(n444) );
  XNOR2_X1 U509 ( .A(G1GAT), .B(G64GAT), .ZN(n443) );
  XNOR2_X1 U510 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U511 ( .A(KEYINPUT80), .B(n445), .Z(n447) );
  NAND2_X1 U512 ( .A1(G231GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U514 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U515 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n451) );
  XNOR2_X1 U516 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n450) );
  XNOR2_X1 U517 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U518 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U519 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U520 ( .A(n457), .B(n456), .Z(n588) );
  NOR2_X1 U521 ( .A1(n593), .A2(n588), .ZN(n458) );
  NAND2_X1 U522 ( .A1(n503), .A2(n458), .ZN(n459) );
  NAND2_X1 U523 ( .A1(n526), .A2(n493), .ZN(n461) );
  INV_X1 U524 ( .A(n352), .ZN(n571) );
  NAND2_X1 U525 ( .A1(n541), .A2(n571), .ZN(n464) );
  INV_X1 U526 ( .A(n465), .ZN(n513) );
  NAND2_X1 U527 ( .A1(n541), .A2(n513), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(G1339GAT) );
  INV_X1 U529 ( .A(KEYINPUT54), .ZN(n482) );
  INV_X1 U530 ( .A(n491), .ZN(n580) );
  NAND2_X1 U531 ( .A1(n580), .A2(n570), .ZN(n468) );
  XNOR2_X1 U532 ( .A(n468), .B(KEYINPUT46), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n469), .A2(n472), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n567), .A2(n470), .ZN(n471) );
  XNOR2_X1 U535 ( .A(KEYINPUT47), .B(n471), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n593), .A2(n472), .ZN(n473) );
  XNOR2_X1 U537 ( .A(KEYINPUT45), .B(n473), .ZN(n475) );
  INV_X1 U538 ( .A(n585), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U540 ( .A(KEYINPUT119), .B(n476), .ZN(n477) );
  NAND2_X1 U541 ( .A1(n477), .A2(n491), .ZN(n478) );
  NAND2_X1 U542 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U543 ( .A1(n558), .A2(n540), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U545 ( .A1(n483), .A2(n527), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(KEYINPUT64), .ZN(n579) );
  NOR2_X1 U547 ( .A1(n579), .A2(n485), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(KEYINPUT55), .ZN(n572) );
  NAND2_X1 U549 ( .A1(n576), .A2(n567), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n488) );
  INV_X1 U551 ( .A(G190GAT), .ZN(n487) );
  NOR2_X1 U552 ( .A1(n585), .A2(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT78), .ZN(n504) );
  NAND2_X1 U554 ( .A1(n493), .A2(n504), .ZN(n494) );
  NOR2_X1 U555 ( .A1(n523), .A2(n530), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(KEYINPUT112), .ZN(n497) );
  INV_X1 U557 ( .A(G36GAT), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n500) );
  NAND2_X1 U560 ( .A1(n588), .A2(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(n501), .B(KEYINPUT16), .Z(n502) );
  AND2_X1 U563 ( .A1(n503), .A2(n502), .ZN(n525) );
  NAND2_X1 U564 ( .A1(n525), .A2(n504), .ZN(n514) );
  NOR2_X1 U565 ( .A1(n527), .A2(n514), .ZN(n506) );
  XNOR2_X1 U566 ( .A(KEYINPUT107), .B(KEYINPUT34), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G1GAT), .B(n507), .ZN(G1324GAT) );
  NOR2_X1 U569 ( .A1(n530), .A2(n514), .ZN(n508) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(n508), .Z(n509) );
  XNOR2_X1 U571 ( .A(G8GAT), .B(n509), .ZN(G1325GAT) );
  NOR2_X1 U572 ( .A1(n352), .A2(n514), .ZN(n511) );
  XNOR2_X1 U573 ( .A(KEYINPUT109), .B(KEYINPUT35), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U575 ( .A(G15GAT), .B(n512), .Z(G1326GAT) );
  INV_X1 U576 ( .A(n513), .ZN(n534) );
  NOR2_X1 U577 ( .A1(n534), .A2(n514), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(n515), .Z(n516) );
  XNOR2_X1 U579 ( .A(G22GAT), .B(n516), .ZN(G1327GAT) );
  NOR2_X1 U580 ( .A1(n523), .A2(n527), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1328GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT40), .B(KEYINPUT114), .Z(n520) );
  XNOR2_X1 U584 ( .A(G43GAT), .B(KEYINPUT113), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n522) );
  NOR2_X1 U586 ( .A1(n352), .A2(n523), .ZN(n521) );
  XOR2_X1 U587 ( .A(n522), .B(n521), .Z(G1330GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n534), .ZN(n524) );
  XOR2_X1 U589 ( .A(G50GAT), .B(n524), .Z(G1331GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n527), .A2(n533), .ZN(n528) );
  XOR2_X1 U592 ( .A(G57GAT), .B(n528), .Z(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT42), .B(n529), .ZN(G1332GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n533), .ZN(n531) );
  XOR2_X1 U595 ( .A(G64GAT), .B(n531), .Z(G1333GAT) );
  NOR2_X1 U596 ( .A1(n352), .A2(n533), .ZN(n532) );
  XOR2_X1 U597 ( .A(G71GAT), .B(n532), .Z(G1334GAT) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT43), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(G78GAT), .B(n537), .Z(G1335GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n541), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G85GAT), .B(n539), .ZN(G1336GAT) );
  XOR2_X1 U604 ( .A(G92GAT), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(G1337GAT) );
  NOR2_X1 U607 ( .A1(n352), .A2(n544), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n545), .A2(n558), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(n546), .Z(n553) );
  NAND2_X1 U610 ( .A1(n553), .A2(n580), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U613 ( .A1(n553), .A2(n570), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(G120GAT), .B(n550), .Z(G1341GAT) );
  NAND2_X1 U616 ( .A1(n553), .A2(n588), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT50), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n567), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G134GAT), .B(n556), .ZN(G1343GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n578), .A2(n559), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n580), .A2(n566), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U628 ( .A1(n566), .A2(n570), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  XOR2_X1 U631 ( .A(G155GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n588), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n580), .A2(n576), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n574) );
  OR2_X1 U639 ( .A1(n294), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G176GAT), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U642 ( .A1(n576), .A2(n588), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .Z(n582) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n591), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U651 ( .A1(n591), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n591), .A2(n588), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(KEYINPUT126), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G211GAT), .B(n590), .ZN(G1354GAT) );
  INV_X1 U656 ( .A(n591), .ZN(n592) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

