//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT66), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NOR4_X1   g043(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT66), .A4(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n461), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT65), .B(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(KEYINPUT66), .B(new_n477), .C1(new_n488), .C2(new_n468), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n466), .A2(new_n490), .A3(KEYINPUT3), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n461), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n492), .B2(G124), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n489), .B2(new_n491), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n461), .A3(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n479), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n461), .C1(new_n467), .C2(new_n469), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n504), .A2(KEYINPUT67), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(KEYINPUT67), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n469), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n502), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n515), .B2(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n519), .B(G651), .C1(new_n512), .C2(new_n513), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n511), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n521), .A2(G50), .B1(G651), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n518), .B2(new_n520), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT70), .B(G88), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND2_X1  g107(.A1(new_n528), .A2(G89), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n536), .A2(KEYINPUT7), .A3(new_n537), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n521), .A2(G51), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n533), .A2(new_n542), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n524), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G52), .B1(G651), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n528), .A2(G90), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(new_n528), .A2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n521), .A2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G651), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(new_n515), .ZN(new_n566));
  NAND2_X1  g141(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n556), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n520), .B1(new_n568), .B2(new_n516), .ZN(new_n569));
  AND2_X1   g144(.A1(KEYINPUT72), .A2(G53), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(G543), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n524), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n528), .A2(G91), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n572), .A2(KEYINPUT73), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT73), .B1(new_n572), .B2(new_n576), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n556), .B1(new_n524), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n528), .B2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n521), .A2(G49), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  AND2_X1   g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n523), .B2(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n588), .B2(new_n556), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OR2_X1    g165(.A1(KEYINPUT5), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(KEYINPUT5), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g168(.A(KEYINPUT74), .B(G651), .C1(new_n593), .C2(new_n587), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n569), .A2(G86), .A3(new_n523), .ZN(new_n596));
  AND2_X1   g171(.A1(G48), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n569), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n524), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n521), .A2(G47), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n528), .A2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(new_n556), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n569), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G54), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n528), .A2(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G280));
  XOR2_X1   g196(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n559), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n623), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n625), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n492), .A2(G123), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT78), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(KEYINPUT79), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n634), .A2(KEYINPUT79), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n494), .A2(G135), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2096), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n479), .A2(new_n466), .A3(G2105), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2443), .B(G2446), .Z(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n658), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n666), .B2(KEYINPUT81), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(KEYINPUT81), .B2(new_n666), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n666), .B(KEYINPUT17), .Z(new_n673));
  INV_X1    g248(.A(new_n667), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n665), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT85), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1981), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(G171), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G5), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1341), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n559), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G16), .B2(G19), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n706), .A2(G1961), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n703), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n703), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n710), .B1(new_n707), .B2(new_n709), .C1(G1966), .C2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT29), .Z(new_n717));
  INV_X1    g292(.A(G2090), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n721));
  OAI22_X1  g296(.A1(G160), .A2(new_n714), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT95), .B(G2084), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n722), .A2(new_n724), .B1(G1966), .B2(new_n712), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n725), .B1(new_n722), .B2(new_n724), .C1(new_n706), .C2(G1961), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n713), .A2(new_n719), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n717), .A2(new_n718), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT99), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G11), .ZN(new_n730));
  INV_X1    g305(.A(G28), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n731), .B2(KEYINPUT30), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI22_X1  g308(.A1(new_n733), .A2(KEYINPUT98), .B1(KEYINPUT30), .B2(new_n731), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n730), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n714), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT94), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n494), .A2(G139), .ZN(new_n741));
  INV_X1    g316(.A(new_n479), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n742), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n741), .C1(new_n461), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(new_n442), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n736), .B(new_n746), .C1(G29), .C2(new_n639), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(new_n443), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n714), .A2(G32), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT26), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(KEYINPUT26), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(G105), .B2(new_n471), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n494), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n492), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(new_n714), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n616), .A2(new_n703), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G4), .B2(new_n703), .ZN(new_n766));
  INV_X1    g341(.A(G1348), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n747), .A2(new_n751), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n745), .A2(new_n442), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT96), .Z(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n443), .B2(new_n750), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n714), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n494), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n492), .A2(G128), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n461), .A2(G116), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n767), .B2(new_n766), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n769), .A2(new_n772), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G299), .A2(G16), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n703), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n727), .A2(new_n729), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n703), .A2(G22), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n703), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  MUX2_X1   g372(.A(G6), .B(G305), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT90), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT32), .B(G1981), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n796), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n703), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(G288), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n703), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n799), .B2(new_n801), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n803), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n714), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n494), .A2(G131), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n492), .A2(G119), .ZN(new_n817));
  OR2_X1    g392(.A1(G95), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n714), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n703), .A2(G24), .ZN(new_n825));
  INV_X1    g400(.A(G290), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n703), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT88), .B(G1986), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n813), .A2(new_n814), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT92), .B1(new_n812), .B2(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n811), .B1(new_n803), .B2(new_n809), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n834), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n791), .B1(new_n837), .B2(new_n839), .ZN(G311));
  INV_X1    g415(.A(new_n791), .ZN(new_n841));
  INV_X1    g416(.A(new_n839), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n838), .B1(new_n834), .B2(new_n835), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(G150));
  NAND2_X1  g419(.A1(new_n521), .A2(G55), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n569), .A2(G93), .A3(new_n523), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n556), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT100), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n851), .A3(new_n846), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n558), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n559), .A3(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT38), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n616), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n860), .A2(new_n861), .A3(G860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n849), .A2(G860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n780), .B(new_n760), .ZN(new_n866));
  XNOR2_X1  g441(.A(G164), .B(KEYINPUT101), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n494), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n492), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n461), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n644), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n820), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n870), .B(new_n879), .C1(new_n868), .C2(new_n869), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n871), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n871), .A2(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n483), .B(new_n496), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n639), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(new_n892), .A3(new_n881), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT40), .B1(new_n891), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(G395));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n849), .B2(new_n619), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n628), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n626), .B(KEYINPUT76), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n856), .ZN(new_n907));
  INV_X1    g482(.A(new_n856), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(new_n616), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n578), .A2(new_n579), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n572), .A2(new_n576), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT73), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n616), .B1(new_n915), .B2(new_n577), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n910), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n578), .B2(new_n579), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n577), .A3(new_n616), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n907), .A2(new_n909), .A3(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n919), .ZN(new_n924));
  INV_X1    g499(.A(new_n909), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n908), .B1(new_n903), .B2(new_n905), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n922), .A3(KEYINPUT105), .ZN(new_n928));
  XOR2_X1   g503(.A(G290), .B(G288), .Z(new_n929));
  XOR2_X1   g504(.A(G303), .B(G305), .Z(new_n930));
  XOR2_X1   g505(.A(new_n929), .B(new_n930), .Z(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT42), .Z(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G868), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n923), .B2(new_n928), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n901), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(new_n900), .A3(G868), .A4(new_n933), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(G295));
  AND2_X1   g514(.A1(new_n936), .A2(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  XNOR2_X1  g516(.A(G301), .B(G286), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n850), .A2(new_n559), .A3(new_n852), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n559), .B1(new_n850), .B2(new_n852), .ZN(new_n944));
  OR3_X1    g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n945), .A2(new_n924), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n856), .A2(new_n949), .A3(new_n942), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n945), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n947), .B1(new_n952), .B2(new_n921), .ZN(new_n953));
  INV_X1    g528(.A(new_n931), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n951), .A2(new_n924), .A3(new_n945), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n917), .A2(new_n920), .B1(new_n945), .B2(new_n946), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n931), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n951), .A2(new_n945), .B1(new_n917), .B2(new_n920), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n931), .B1(new_n962), .B2(new_n947), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n941), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n945), .A2(new_n924), .A3(new_n946), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n917), .A2(new_n920), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n856), .A2(new_n942), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n948), .B2(new_n950), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n954), .B(new_n966), .C1(new_n967), .C2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n963), .A2(new_n970), .A3(new_n961), .A4(new_n894), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n955), .A2(new_n973), .A3(new_n961), .A4(new_n963), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n941), .B1(new_n959), .B2(KEYINPUT43), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT109), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT109), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n965), .B1(new_n977), .B2(new_n978), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n502), .B2(new_n509), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n473), .A2(G40), .A3(new_n482), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT110), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n826), .ZN(new_n990));
  INV_X1    g565(.A(G2067), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n780), .B(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n760), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n821), .A2(new_n823), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n821), .A2(new_n823), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n985), .B1(new_n990), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT114), .B(G8), .Z(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G286), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n980), .C1(new_n502), .C2(new_n509), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n981), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n984), .A2(G2084), .ZN(new_n1009));
  INV_X1    g584(.A(G1966), .ZN(new_n1010));
  AND4_X1   g585(.A1(G40), .A2(new_n470), .A3(new_n482), .A4(new_n472), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n980), .C1(new_n502), .C2(new_n509), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n983), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1008), .A2(new_n1009), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1001), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1013), .A2(new_n1010), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1009), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1019));
  OAI211_X1 g594(.A(G286), .B(new_n1000), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(KEYINPUT51), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(new_n1001), .C1(new_n1014), .C2(new_n999), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT62), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n583), .A2(G1976), .A3(new_n584), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1000), .B(new_n1028), .C1(new_n981), .C2(new_n984), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n492), .A2(G126), .B1(new_n505), .B2(new_n506), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n498), .B1(new_n494), .B2(G138), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n500), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(new_n980), .A3(new_n1011), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1035), .A2(KEYINPUT115), .A3(new_n1000), .A4(new_n1028), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  OAI21_X1  g615(.A(G651), .B1(new_n593), .B2(new_n587), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n598), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT118), .B(G86), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n1043), .B(new_n524), .C1(new_n518), .C2(new_n520), .ZN(new_n1044));
  OAI21_X1  g619(.A(G1981), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n595), .A2(new_n1046), .A3(new_n596), .A4(new_n598), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1035), .A3(new_n1000), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1040), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n981), .A2(new_n984), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n999), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1056), .A2(new_n1058), .A3(KEYINPUT120), .A4(new_n1051), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1031), .A2(KEYINPUT116), .A3(new_n1036), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT117), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1064), .A2(new_n1029), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n1039), .A2(new_n1060), .A3(new_n1061), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G166), .A2(new_n1015), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(KEYINPUT113), .B2(KEYINPUT55), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n984), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1071), .A2(new_n718), .B1(new_n1013), .B2(new_n795), .ZN(new_n1072));
  OAI221_X1 g647(.A(new_n1068), .B1(new_n1067), .B2(new_n1069), .C1(new_n1072), .C2(new_n999), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1068), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1013), .A2(new_n795), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1013), .A2(new_n1077), .A3(new_n795), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(G2090), .B(new_n984), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1080));
  OAI211_X1 g655(.A(G8), .B(new_n1074), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1066), .A2(new_n1073), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1021), .A2(KEYINPUT62), .A3(new_n1023), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n983), .A2(new_n1012), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1011), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1013), .B2(G2078), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n984), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1085), .B(new_n1087), .C1(new_n1088), .C2(G1961), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1026), .A2(new_n1082), .A3(new_n1083), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1081), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1060), .A2(new_n1062), .A3(new_n805), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1047), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1056), .B(KEYINPUT121), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1092), .A2(new_n1066), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(new_n913), .B(KEYINPUT57), .Z(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n789), .B1(new_n1070), .B2(new_n984), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n983), .A2(new_n1011), .A3(new_n1012), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(KEYINPUT123), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1098), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n981), .B2(new_n984), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1034), .A2(KEYINPUT124), .A3(new_n980), .A4(new_n1011), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n991), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1088), .B2(G1348), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1105), .B1(new_n1112), .B2(new_n911), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(new_n1099), .A3(new_n1097), .A4(new_n1103), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n983), .A2(new_n993), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT58), .B(G1341), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1109), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n559), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(KEYINPUT59), .A3(new_n559), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT60), .B(new_n1110), .C1(new_n1088), .C2(G1348), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1122), .B(new_n1123), .C1(new_n616), .C2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1112), .A2(KEYINPUT60), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1124), .A2(new_n616), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1105), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT61), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1116), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1088), .A2(G1961), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1134), .A2(new_n1087), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G301), .B(KEYINPUT54), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n443), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1137));
  INV_X1    g712(.A(new_n473), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n481), .A2(KEYINPUT125), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n461), .B1(new_n481), .B2(KEYINPUT125), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1137), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1084), .B2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1135), .A2(new_n1142), .B1(new_n1089), .B2(new_n1136), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1082), .A2(new_n1133), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1091), .B(new_n1096), .C1(new_n1132), .C2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1015), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1066), .B1(new_n1147), .B2(new_n1074), .ZN(new_n1148));
  OAI211_X1 g723(.A(G168), .B(new_n1000), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1081), .A2(KEYINPUT63), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  AND4_X1   g727(.A1(new_n1066), .A2(new_n1073), .A3(new_n1081), .A4(new_n1150), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n1153), .B2(KEYINPUT122), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1066), .A2(new_n1073), .A3(new_n1081), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n1149), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1152), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n998), .B1(new_n1145), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n987), .A2(new_n985), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1162), .B(new_n1163), .C1(new_n985), .C2(new_n997), .ZN(new_n1164));
  INV_X1    g739(.A(new_n992), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n985), .B1(new_n1165), .B2(new_n760), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n985), .A2(new_n993), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1167), .A2(KEYINPUT46), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1167), .A2(KEYINPUT46), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1166), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT47), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n992), .A2(new_n994), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1172), .A2(new_n995), .B1(G2067), .B2(new_n780), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1164), .B(new_n1171), .C1(new_n985), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1159), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(G319), .ZN(new_n1177));
  NOR2_X1   g751(.A1(G227), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g752(.A(new_n1178), .B(KEYINPUT127), .ZN(new_n1179));
  NOR3_X1   g753(.A1(G229), .A2(G401), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n892), .B1(new_n886), .B2(new_n887), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n1181), .B2(new_n895), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n960), .A2(new_n964), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1183), .ZN(G308));
  INV_X1    g758(.A(G308), .ZN(G225));
endmodule


