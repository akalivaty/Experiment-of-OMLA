//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT0), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT0), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n191), .B(KEYINPUT64), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT0), .B(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(KEYINPUT0), .A3(G128), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n196), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n205), .A2(KEYINPUT3), .A3(G104), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT3), .B1(new_n205), .B2(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G101), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n210), .B(new_n204), .C1(new_n206), .C2(new_n207), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n213), .A3(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT10), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  AND4_X1   g031(.A1(new_n217), .A2(new_n188), .A3(new_n190), .A4(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n188), .A2(KEYINPUT77), .A3(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(G128), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n223), .B2(new_n191), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  XNOR2_X1  g039(.A(G104), .B(G107), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n210), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n205), .A2(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n204), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT76), .A3(G101), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n211), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n216), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n227), .A2(new_n230), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n217), .B1(G143), .B2(new_n187), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n191), .B1(new_n234), .B2(new_n194), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n198), .A2(new_n217), .A3(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n211), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n215), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G131), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n244), .A2(new_n246), .A3(new_n250), .A4(new_n247), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n215), .A2(new_n232), .A3(KEYINPUT80), .A4(new_n238), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n241), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n257), .A2(new_n258), .B1(G131), .B2(new_n248), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n215), .A2(new_n232), .A3(new_n259), .A4(new_n238), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT75), .ZN(new_n264));
  XNOR2_X1  g078(.A(G110), .B(G140), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n264), .B(new_n265), .Z(new_n266));
  NAND3_X1  g080(.A1(new_n260), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n261), .B1(new_n260), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n237), .B1(new_n233), .B2(new_n211), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n224), .A2(new_n231), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n254), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n237), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n231), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n224), .B2(new_n231), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n280), .A2(KEYINPUT78), .A3(new_n274), .A4(new_n254), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n260), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n266), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n270), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G469), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT81), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n260), .A2(new_n266), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT79), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n267), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n291), .A2(new_n256), .B1(new_n283), .B2(new_n282), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n288), .B(G469), .C1(new_n292), .C2(G902), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT82), .B(G469), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n289), .A2(KEYINPUT83), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n277), .A2(new_n281), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n260), .B2(new_n266), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n266), .B1(new_n256), .B2(new_n260), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n294), .B(new_n295), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n287), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT68), .B(G116), .ZN(new_n304));
  INV_X1    g118(.A(G122), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(G116), .B2(new_n305), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n205), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n189), .A2(G128), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n194), .A2(G143), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(KEYINPUT13), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT87), .B1(new_n310), .B2(KEYINPUT13), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n310), .A2(KEYINPUT87), .A3(KEYINPUT13), .ZN(new_n314));
  OAI21_X1  g128(.A(G134), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n310), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n243), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n308), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT14), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  OAI22_X1  g134(.A1(new_n306), .A2(new_n319), .B1(new_n320), .B2(G122), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n304), .A2(KEYINPUT14), .A3(new_n305), .ZN(new_n322));
  OAI21_X1  g136(.A(G107), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT88), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n307), .A2(new_n205), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(G107), .C1(new_n321), .C2(new_n322), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n316), .B(new_n243), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT9), .B(G234), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G217), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n331), .A2(new_n332), .A3(G953), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n318), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n318), .B2(new_n329), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n294), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G478), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT15), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI221_X1 g153(.A(new_n294), .B1(KEYINPUT15), .B2(new_n337), .C1(new_n334), .C2(new_n335), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G952), .ZN(new_n342));
  AOI211_X1 g156(.A(G953), .B(new_n342), .C1(G234), .C2(G237), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT21), .B(G898), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n294), .B(new_n262), .C1(G234), .C2(G237), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n262), .A3(G214), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n189), .ZN(new_n352));
  NOR2_X1   g166(.A1(G237), .A2(G953), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G131), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n250), .A3(new_n354), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT16), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT72), .A2(G125), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(new_n359), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n364), .B2(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  INV_X1    g180(.A(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G140), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT19), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n360), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n364), .B2(new_n369), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n358), .B(new_n366), .C1(G146), .C2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n360), .A3(new_n187), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n364), .B2(new_n187), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT18), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n250), .ZN(new_n376));
  OAI221_X1 g190(.A(new_n374), .B1(new_n355), .B2(new_n376), .C1(new_n356), .C2(new_n375), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G113), .B(G122), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n203), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n358), .A2(KEYINPUT17), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n187), .B(new_n362), .C1(new_n364), .C2(new_n361), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n355), .A2(KEYINPUT17), .A3(G131), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n366), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n380), .B(new_n377), .C1(new_n383), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(G475), .A2(G902), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n348), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT20), .B(new_n391), .C1(new_n382), .C2(new_n387), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n377), .B1(new_n383), .B2(new_n386), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n381), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n394), .B2(new_n387), .ZN(new_n395));
  INV_X1    g209(.A(G475), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n390), .A2(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n341), .A2(new_n347), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G221), .B1(new_n331), .B2(G902), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT74), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G210), .B1(G237), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n320), .A2(G119), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G119), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n304), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT2), .B(G113), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(new_n407), .C1(new_n408), .C2(new_n304), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n212), .A2(new_n414), .A3(new_n214), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(G113), .B(new_n417), .C1(new_n409), .C2(new_n416), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(new_n233), .A3(new_n211), .A4(new_n413), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G122), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n419), .A3(new_n421), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(G224), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n196), .A2(new_n200), .A3(new_n201), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n278), .A2(new_n367), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n428), .B1(new_n427), .B2(G125), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n262), .B(new_n426), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n432), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n426), .A2(new_n262), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n430), .A4(new_n429), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n420), .A2(new_n438), .A3(new_n422), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n425), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n429), .A2(new_n430), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n441), .A2(KEYINPUT7), .A3(new_n435), .A4(new_n434), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(KEYINPUT7), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n431), .B2(new_n432), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n421), .B(KEYINPUT8), .ZN(new_n445));
  INV_X1    g259(.A(new_n419), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n413), .A2(new_n418), .B1(new_n233), .B2(new_n211), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n444), .A3(new_n424), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n294), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n405), .B1(new_n440), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n425), .A2(new_n437), .A3(new_n439), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n294), .A3(new_n404), .A4(new_n449), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n403), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n303), .A2(new_n398), .A3(new_n401), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n251), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n245), .A2(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n247), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G131), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n237), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n458), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n254), .A2(new_n202), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n257), .A2(new_n258), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n235), .A2(new_n236), .B1(G131), .B2(new_n462), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT66), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n467), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT30), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n473), .A2(new_n414), .A3(new_n475), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n353), .A2(G210), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n210), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n482), .B(new_n483), .Z(new_n484));
  INV_X1    g298(.A(new_n414), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n466), .A2(new_n485), .A3(new_n476), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT31), .ZN(new_n488));
  INV_X1    g302(.A(new_n486), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT28), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n470), .A2(new_n414), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n486), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(new_n484), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT31), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n480), .A2(new_n496), .A3(new_n484), .A4(new_n486), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n488), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G472), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n294), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(KEYINPUT32), .A3(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n480), .A2(new_n486), .ZN(new_n506));
  INV_X1    g320(.A(new_n484), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT29), .B1(new_n494), .B2(new_n484), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n477), .A2(new_n414), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT71), .A3(new_n486), .ZN(new_n512));
  OR3_X1    g326(.A1(new_n477), .A2(KEYINPUT71), .A3(new_n414), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n490), .B1(new_n514), .B2(KEYINPUT28), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT29), .A3(new_n484), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n294), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G472), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n504), .A2(new_n505), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n451), .A2(new_n453), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n402), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n395), .A2(new_n396), .ZN(new_n522));
  INV_X1    g336(.A(new_n390), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n388), .A2(new_n348), .A3(new_n389), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n347), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n339), .A4(new_n340), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(KEYINPUT89), .A3(new_n401), .A4(new_n303), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n332), .B1(G234), .B2(new_n294), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n366), .A2(new_n384), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n194), .A2(G119), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n408), .A2(G128), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT24), .B(G110), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT23), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n535), .A2(new_n539), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n541), .A2(new_n542), .B1(G119), .B2(new_n194), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G110), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n533), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n543), .A2(G110), .B1(new_n536), .B2(new_n537), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n373), .A3(new_n366), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT22), .B(G137), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n532), .B1(new_n555), .B2(G902), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT25), .A4(new_n294), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n531), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n531), .A2(new_n294), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT73), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n554), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n457), .A2(new_n519), .A3(new_n529), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n451), .A2(KEYINPUT90), .A3(new_n453), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n402), .B1(new_n451), .B2(KEYINPUT90), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n450), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n404), .B1(new_n572), .B2(new_n452), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n403), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n451), .A2(KEYINPUT90), .A3(new_n453), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(KEYINPUT91), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n318), .A2(new_n329), .A3(new_n333), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(KEYINPUT92), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n334), .B2(new_n335), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n318), .A2(new_n329), .ZN(new_n582));
  INV_X1    g396(.A(new_n333), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(new_n579), .C1(KEYINPUT92), .C2(new_n578), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n337), .A2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n336), .A2(new_n337), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n525), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND4_X1   g404(.A1(new_n526), .A2(new_n571), .A3(new_n577), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n498), .A2(new_n294), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n592), .A2(G472), .B1(new_n498), .B2(new_n501), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n303), .A2(new_n565), .A3(new_n401), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT34), .B(G104), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  INV_X1    g411(.A(new_n341), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n397), .ZN(new_n599));
  AND4_X1   g413(.A1(new_n526), .A2(new_n571), .A3(new_n577), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n593), .A3(new_n594), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NOR2_X1   g418(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n548), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n562), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n559), .A2(KEYINPUT94), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n609));
  INV_X1    g423(.A(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n558), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n457), .A2(new_n529), .A3(new_n593), .A4(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT37), .B(G110), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G12));
  AND2_X1   g429(.A1(new_n303), .A2(new_n401), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n519), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n571), .A2(new_n577), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n611), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n343), .B1(new_n346), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n598), .A2(new_n397), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  XOR2_X1   g439(.A(new_n520), .B(KEYINPUT38), .Z(new_n626));
  NOR2_X1   g440(.A1(new_n598), .A2(new_n525), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n619), .A2(new_n402), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n622), .B(KEYINPUT39), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n616), .A2(new_n630), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n626), .B(new_n628), .C1(new_n631), .C2(KEYINPUT40), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n498), .A2(KEYINPUT32), .A3(new_n501), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT32), .B1(new_n498), .B2(new_n501), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n499), .A2(new_n294), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n499), .B1(new_n514), .B2(new_n507), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n637), .B2(new_n487), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT95), .Z(new_n639));
  AOI21_X1  g453(.A(KEYINPUT96), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n635), .A2(KEYINPUT96), .A3(new_n639), .ZN(new_n641));
  OAI221_X1 g455(.A(new_n632), .B1(KEYINPUT40), .B2(new_n631), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G143), .ZN(G45));
  INV_X1    g457(.A(new_n622), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n590), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n620), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G146), .ZN(G48));
  INV_X1    g462(.A(new_n300), .ZN(new_n649));
  INV_X1    g463(.A(new_n301), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n401), .B(new_n302), .C1(new_n651), .C2(new_n286), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT97), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n591), .A2(new_n653), .A3(new_n565), .A4(new_n519), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND4_X1  g470(.A1(new_n600), .A2(new_n653), .A3(new_n565), .A4(new_n519), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  NOR2_X1   g472(.A1(new_n618), .A2(new_n652), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n619), .A2(new_n527), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n519), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G119), .ZN(G21));
  AND4_X1   g476(.A1(new_n526), .A2(new_n571), .A3(new_n577), .A4(new_n627), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n592), .A2(G472), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n488), .B(new_n497), .C1(new_n515), .C2(new_n484), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n501), .B(KEYINPUT98), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n664), .A2(new_n565), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n663), .A2(new_n668), .A3(new_n653), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G122), .ZN(G24));
  NAND3_X1  g484(.A1(new_n664), .A2(new_n612), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT99), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n664), .A2(new_n612), .A3(new_n673), .A4(new_n667), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n645), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n659), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G125), .ZN(G27));
  AOI21_X1  g491(.A(new_n564), .B1(new_n635), .B2(new_n518), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n284), .A2(KEYINPUT101), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n282), .B2(new_n283), .ZN(new_n681));
  OAI211_X1 g495(.A(G469), .B(new_n270), .C1(new_n679), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(G469), .A2(G902), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT100), .Z(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n302), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n520), .A2(new_n403), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n685), .A2(new_n686), .A3(new_n401), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n678), .A2(KEYINPUT102), .A3(new_n646), .A4(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n519), .A2(new_n565), .A3(new_n646), .A4(new_n687), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT42), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n678), .A2(KEYINPUT42), .A3(new_n646), .A4(new_n687), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n688), .A2(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n691), .A2(new_n693), .A3(new_n688), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(G131), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G33));
  NAND4_X1  g512(.A1(new_n519), .A2(new_n565), .A3(new_n623), .A4(new_n687), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G134), .ZN(G36));
  INV_X1    g516(.A(new_n686), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n588), .A2(new_n589), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(KEYINPUT107), .B2(KEYINPUT43), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n705), .B(new_n525), .C1(KEYINPUT107), .C2(new_n704), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n707), .A2(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n525), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(KEYINPUT106), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n612), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n593), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n703), .B1(new_n714), .B2(KEYINPUT44), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(KEYINPUT44), .B2(new_n714), .ZN(new_n716));
  OAI211_X1 g530(.A(KEYINPUT45), .B(new_n270), .C1(new_n679), .C2(new_n681), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n717), .B(G469), .C1(KEYINPUT45), .C2(new_n292), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(new_n684), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n719), .A2(KEYINPUT46), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n302), .B1(new_n719), .B2(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n401), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(new_n629), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G137), .ZN(G39));
  XOR2_X1   g539(.A(new_n722), .B(KEYINPUT47), .Z(new_n726));
  NOR4_X1   g540(.A1(new_n519), .A2(new_n565), .A3(new_n645), .A4(new_n703), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G140), .ZN(G42));
  OR2_X1    g543(.A1(new_n590), .A2(new_n599), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n521), .A2(new_n347), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n594), .A3(new_n593), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n566), .A2(new_n613), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n566), .A2(new_n613), .A3(new_n732), .A4(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND4_X1   g551(.A1(new_n654), .A2(new_n657), .A3(new_n669), .A4(new_n661), .ZN(new_n738));
  INV_X1    g552(.A(new_n617), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n598), .A2(new_n525), .A3(new_n644), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n703), .A2(new_n619), .A3(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n675), .A2(new_n687), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n701), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT110), .B1(new_n743), .B2(new_n696), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n691), .A2(new_n688), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n692), .A2(new_n693), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(KEYINPUT103), .B2(new_n745), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n738), .A2(new_n742), .A3(new_n701), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n737), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n618), .A2(new_n619), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n739), .B(new_n752), .C1(new_n623), .C2(new_n646), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n641), .A2(new_n640), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n571), .A2(new_n577), .A3(new_n627), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n558), .A2(new_n610), .A3(new_n622), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n401), .A3(new_n685), .A4(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n676), .B(new_n753), .C1(new_n754), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n744), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT54), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n743), .A2(new_n696), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n768), .A3(KEYINPUT53), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n763), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT111), .B1(new_n762), .B2(new_n763), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n767), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n652), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n343), .A3(new_n686), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n712), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n674), .B2(new_n672), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n712), .A2(new_n343), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n668), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n626), .A2(new_n774), .A3(new_n403), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n777), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n779), .B2(new_n703), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n302), .B1(new_n651), .B2(new_n286), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(new_n401), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n790), .B1(new_n726), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n779), .A2(new_n789), .A3(new_n703), .ZN(new_n795));
  OAI221_X1 g609(.A(new_n788), .B1(new_n787), .B2(new_n786), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n754), .A2(new_n565), .A3(new_n775), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT116), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n397), .A3(new_n704), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n796), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n797), .B1(new_n796), .B2(new_n800), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n525), .B(new_n799), .C1(new_n589), .C2(new_n588), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n779), .A2(new_n618), .A3(new_n652), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n712), .A2(new_n678), .A3(new_n775), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT48), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n342), .B(G953), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n808), .A2(KEYINPUT48), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n807), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n805), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n806), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n803), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n801), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n773), .A2(new_n816), .B1(G952), .B2(G953), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n704), .A2(new_n401), .A3(new_n525), .A4(new_n402), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n626), .C1(KEYINPUT49), .C2(new_n791), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(KEYINPUT49), .B2(new_n791), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n754), .A3(new_n565), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT108), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n817), .A2(KEYINPUT119), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(G75));
  NAND2_X1  g642(.A1(new_n762), .A2(new_n763), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n763), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n294), .B1(new_n833), .B2(new_n769), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(G210), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n425), .A2(new_n439), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(new_n437), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT55), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n835), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n835), .B2(new_n836), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n262), .A2(G952), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G51));
  OAI21_X1  g657(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n766), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(KEYINPUT120), .A3(new_n772), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n844), .A2(new_n847), .A3(new_n766), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n684), .B(KEYINPUT57), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n649), .A2(new_n650), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n834), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(new_n718), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n842), .B1(new_n852), .B2(new_n854), .ZN(G54));
  NAND3_X1  g669(.A1(new_n834), .A2(KEYINPUT58), .A3(G475), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n382), .A2(new_n387), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(new_n842), .ZN(G60));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n337), .A2(new_n294), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n586), .A2(new_n846), .A3(new_n848), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n586), .B1(new_n773), .B2(new_n864), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n865), .A2(new_n842), .A3(new_n866), .ZN(G63));
  NAND2_X1  g681(.A1(G217), .A2(G902), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT60), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n844), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n842), .B1(new_n871), .B2(new_n555), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n833), .B2(new_n769), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n606), .B(KEYINPUT122), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n873), .A2(new_n844), .A3(new_n870), .A4(new_n875), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(KEYINPUT61), .B(new_n872), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(G66));
  INV_X1    g696(.A(new_n426), .ZN(new_n883));
  OAI21_X1  g697(.A(G953), .B1(new_n345), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n737), .A2(new_n738), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n886), .B2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n837), .B1(G898), .B2(new_n262), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G69));
  NAND3_X1  g703(.A1(new_n473), .A2(new_n475), .A3(new_n479), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT124), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n371), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n676), .A2(new_n753), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n642), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT62), .Z(new_n895));
  AND2_X1   g709(.A1(new_n730), .A2(new_n686), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n678), .A2(new_n896), .A3(new_n616), .A4(new_n630), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n724), .A2(new_n895), .A3(new_n728), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n892), .B1(new_n898), .B2(G953), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n892), .B1(G900), .B2(G953), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n678), .A2(new_n756), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n723), .B1(new_n716), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n893), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(new_n748), .A3(new_n701), .A4(new_n728), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n900), .B1(new_n905), .B2(G953), .ZN(new_n906));
  INV_X1    g720(.A(G227), .ZN(new_n907));
  OAI21_X1  g721(.A(G953), .B1(new_n907), .B2(new_n621), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n899), .A2(new_n906), .B1(KEYINPUT125), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(KEYINPUT125), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(G72));
  XNOR2_X1  g725(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n636), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n905), .B2(new_n885), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n506), .A2(new_n484), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n842), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n508), .A2(new_n487), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n764), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n506), .A2(new_n484), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n898), .A2(new_n886), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n913), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(G57));
endmodule


