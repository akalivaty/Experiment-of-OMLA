//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(new_n207), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n211), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n221), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(G223), .B1(new_n254), .B2(G77), .ZN(new_n255));
  INV_X1    g0055(.A(G222), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n248), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n264), .A2(G274), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n260), .A2(new_n267), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(G226), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n223), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n274), .A2(KEYINPUT66), .A3(G13), .A4(G20), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G50), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n278), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(G50), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n273), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n208), .A2(G20), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n287), .A2(new_n289), .B1(G150), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n284), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n271), .A2(G200), .B1(new_n293), .B2(KEYINPUT9), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n271), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n293), .B1(new_n271), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n301), .A2(KEYINPUT67), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(KEYINPUT67), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n261), .A2(new_n304), .A3(new_n270), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n213), .A2(G1698), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G226), .B2(G1698), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(new_n254), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(new_n260), .B1(new_n269), .B2(G238), .ZN(new_n313));
  INV_X1    g0113(.A(G274), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n262), .B2(new_n263), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n267), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n313), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n299), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(KEYINPUT73), .A3(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n313), .A2(new_n320), .A3(new_n323), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n313), .B2(new_n320), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n326), .B(G169), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G169), .B1(new_n328), .B2(new_n329), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n328), .A2(new_n329), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(KEYINPUT14), .B1(new_n335), .B2(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n279), .A2(G68), .A3(new_n280), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n289), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n339));
  INV_X1    g0139(.A(new_n290), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n207), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT70), .B(KEYINPUT11), .Z(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(new_n273), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n341), .B2(new_n273), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n282), .A2(KEYINPUT12), .A3(G68), .ZN(new_n346));
  XOR2_X1   g0146(.A(new_n346), .B(KEYINPUT71), .Z(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT12), .B1(new_n282), .B2(G68), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT72), .Z(new_n349));
  AOI21_X1  g0149(.A(new_n345), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n335), .A2(G190), .ZN(new_n353));
  OAI21_X1  g0153(.A(G200), .B1(new_n328), .B2(new_n329), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT7), .B1(new_n254), .B2(new_n224), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NOR4_X1   g0158(.A1(new_n252), .A2(new_n253), .A3(new_n358), .A4(G20), .ZN(new_n359));
  OAI21_X1  g0159(.A(G68), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n290), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n204), .A2(new_n205), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G20), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(KEYINPUT74), .A3(G20), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n360), .A2(new_n361), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n363), .A2(KEYINPUT74), .A3(G20), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT74), .B1(new_n363), .B2(G20), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT16), .A3(new_n360), .A4(new_n361), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n273), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n282), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n286), .B1(new_n274), .B2(G20), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n286), .B1(new_n377), .B2(new_n279), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n268), .B1(G232), .B2(new_n269), .ZN(new_n381));
  OAI211_X1 g0181(.A(G223), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n251), .A2(new_n385), .A3(G226), .ZN(new_n386));
  OAI211_X1 g0186(.A(G226), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n381), .B1(new_n389), .B2(new_n264), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n299), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n381), .B(new_n304), .C1(new_n389), .C2(new_n264), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n379), .A2(new_n380), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n381), .B(new_n296), .C1(new_n389), .C2(new_n264), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n269), .A2(G232), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n316), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n382), .A2(new_n383), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n385), .B1(new_n251), .B2(G226), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n401), .B2(new_n260), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n395), .B1(new_n402), .B2(G200), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n375), .A2(new_n403), .A3(new_n378), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n378), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n284), .B1(new_n368), .B2(new_n369), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n374), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n391), .A2(new_n392), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT18), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n394), .A2(new_n406), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n279), .A2(G77), .A3(new_n280), .ZN(new_n414));
  INV_X1    g0214(.A(G77), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n286), .A2(new_n340), .B1(new_n224), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n289), .B2(new_n418), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n414), .B1(G77), .B2(new_n282), .C1(new_n419), .C2(new_n284), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n268), .B1(G244), .B2(new_n269), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n258), .A2(new_n213), .B1(new_n423), .B2(new_n257), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(G238), .B2(new_n251), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n264), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n299), .ZN(new_n427));
  INV_X1    g0227(.A(new_n304), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(new_n426), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G200), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n421), .B(new_n431), .C1(new_n296), .C2(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n308), .A2(new_n356), .A3(new_n413), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT24), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n224), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT22), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT22), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n257), .A2(new_n438), .A3(new_n224), .A4(G87), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT23), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n224), .B2(G107), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n423), .A2(KEYINPUT23), .A3(G20), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n289), .A2(G116), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(KEYINPUT84), .B(new_n435), .C1(new_n440), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n437), .B2(new_n439), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT84), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT24), .B1(new_n448), .B2(new_n449), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n447), .B(new_n273), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n282), .A2(G107), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT25), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n274), .A2(G33), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n282), .A2(new_n284), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n279), .A2(KEYINPUT77), .A3(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(G107), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G257), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n464));
  OAI211_X1 g0264(.A(G250), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n465));
  INV_X1    g0265(.A(G294), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(new_n465), .C1(new_n288), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n260), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n274), .A2(G45), .ZN(new_n469));
  OR2_X1    g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n315), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n260), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G264), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n468), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G169), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n467), .A2(new_n260), .B1(new_n474), .B2(G264), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G179), .A3(new_n473), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n453), .A2(new_n463), .B1(new_n480), .B2(KEYINPUT85), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT85), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n451), .A2(new_n452), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n447), .A2(new_n273), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n462), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G200), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(G190), .B2(new_n476), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n481), .A2(new_n483), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n423), .A2(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n214), .A2(G107), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT76), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(KEYINPUT6), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(KEYINPUT76), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n491), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(new_n500), .A3(G20), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n290), .A2(G77), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n358), .B1(new_n257), .B2(G20), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n423), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n273), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n459), .A2(G97), .A3(new_n460), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n376), .A2(new_n214), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n266), .A2(G1), .ZN(new_n511));
  INV_X1    g0311(.A(new_n471), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n264), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n473), .B1(new_n515), .B2(new_n215), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n428), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(KEYINPUT78), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  OAI211_X1 g0322(.A(G250), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n518), .C2(new_n519), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT78), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n517), .B1(new_n526), .B2(new_n264), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n510), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n518), .A2(new_n519), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n523), .A2(new_n522), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n520), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n516), .B1(new_n534), .B2(new_n260), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(G169), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT79), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n516), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n526), .B2(new_n264), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n299), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT79), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n510), .A4(new_n527), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n535), .A2(G190), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n487), .C2(new_n535), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n537), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G238), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT80), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n257), .A2(KEYINPUT80), .A3(G238), .A4(new_n248), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n257), .A2(G244), .A3(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n260), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n315), .A2(new_n511), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n264), .A2(G250), .A3(new_n469), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n304), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n554), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n299), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n557), .B1(new_n553), .B2(new_n260), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(KEYINPUT81), .A3(new_n304), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n257), .A2(new_n224), .A3(G68), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n289), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR4_X1   g0369(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT82), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G87), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n423), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n309), .A2(new_n568), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G20), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n566), .B(new_n569), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n273), .B1(new_n376), .B2(new_n417), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n459), .A2(new_n418), .A3(new_n460), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n561), .A2(new_n563), .A3(new_n565), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n459), .A2(G87), .A3(new_n460), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n564), .A2(G190), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n562), .A2(G200), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n272), .A2(new_n223), .B1(G20), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n522), .B(new_n224), .C1(G33), .C2(new_n214), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(KEYINPUT20), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n591), .B2(KEYINPUT20), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n279), .A2(G116), .A3(new_n456), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n376), .A2(new_n588), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n589), .A2(KEYINPUT83), .A3(new_n590), .A4(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n257), .A2(G264), .A3(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n257), .A2(G257), .A3(new_n248), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n254), .A2(G303), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n260), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n514), .A2(G270), .A3(new_n264), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n473), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n598), .A2(new_n607), .A3(G169), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(G200), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n605), .B1(new_n260), .B2(new_n602), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G190), .ZN(new_n613));
  INV_X1    g0413(.A(new_n598), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n598), .A2(new_n612), .A3(G179), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n598), .A2(new_n607), .A3(KEYINPUT21), .A4(G169), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n610), .A2(new_n615), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n587), .A2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n434), .A2(new_n490), .A3(new_n546), .A4(new_n619), .ZN(G372));
  NAND2_X1  g0420(.A1(new_n394), .A2(new_n411), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n421), .A2(new_n429), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n337), .A2(new_n351), .B1(new_n623), .B2(new_n355), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n406), .A2(new_n412), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n306), .B1(new_n626), .B2(new_n298), .ZN(new_n627));
  INV_X1    g0427(.A(new_n434), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n610), .A2(new_n616), .A3(new_n617), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n463), .A2(new_n453), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n480), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n489), .A2(new_n463), .A3(new_n453), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n563), .A2(new_n559), .A3(new_n580), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n634), .A2(new_n586), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n546), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n537), .A2(new_n542), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n581), .A2(new_n586), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(new_n635), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n510), .A2(new_n527), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n540), .A2(new_n586), .A3(new_n643), .A4(new_n635), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n637), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n627), .B1(new_n628), .B2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n274), .A2(new_n224), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n614), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n629), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n618), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n480), .A2(KEYINPUT85), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n631), .A2(new_n483), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n634), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n486), .A2(new_n656), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n663), .B2(new_n656), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  AND4_X1   g0467(.A1(new_n663), .A2(new_n634), .A3(new_n629), .A4(new_n656), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n632), .A2(new_n655), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(G399));
  NAND2_X1  g0471(.A1(new_n574), .A2(new_n588), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n227), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(G1), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n222), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n630), .A2(new_n663), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n546), .A2(new_n636), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n586), .A2(new_n643), .A3(new_n540), .A4(new_n635), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n642), .B1(new_n684), .B2(KEYINPUT26), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n656), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n564), .A2(new_n612), .A3(G179), .A4(new_n478), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n539), .ZN(new_n691));
  AND4_X1   g0491(.A1(G179), .A2(new_n478), .A3(new_n603), .A4(new_n606), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(KEYINPUT30), .A3(new_n535), .A4(new_n564), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n428), .B1(new_n603), .B2(new_n606), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n539), .A2(new_n476), .A3(new_n562), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT31), .B1(new_n696), .B2(new_n655), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n546), .A2(new_n490), .A3(new_n619), .A4(new_n656), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n647), .A2(new_n703), .A3(new_n656), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n688), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n680), .B1(new_n706), .B2(G1), .ZN(G364));
  AND2_X1   g0507(.A1(new_n224), .A2(G13), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n274), .B1(new_n708), .B2(G45), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n675), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n661), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G330), .B2(new_n659), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n711), .B(KEYINPUT86), .Z(new_n714));
  NAND2_X1  g0514(.A1(new_n257), .A2(new_n227), .ZN(new_n715));
  INV_X1    g0515(.A(G355), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n715), .A2(new_n716), .B1(G116), .B2(new_n227), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n254), .A2(new_n227), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT87), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n266), .B2(new_n222), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n246), .A2(G45), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n223), .B1(G20), .B2(new_n299), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT88), .Z(new_n728));
  OAI21_X1  g0528(.A(new_n714), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n224), .A2(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n296), .A3(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n423), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(G190), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(G87), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n296), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n301), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n732), .B(new_n735), .C1(G97), .C2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n224), .A2(G190), .A3(G200), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n428), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n254), .B1(new_n741), .B2(G77), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n304), .A2(new_n224), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(new_n736), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n739), .B(new_n742), .C1(new_n202), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n301), .ZN(new_n747));
  INV_X1    g0547(.A(G159), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT89), .B(KEYINPUT32), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(new_n296), .A3(G200), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n751), .B1(new_n207), .B2(new_n752), .C1(new_n203), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n254), .B1(new_n731), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n744), .B2(G322), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n741), .A2(G311), .B1(G303), .B2(new_n734), .ZN(new_n758));
  INV_X1    g0558(.A(new_n747), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G329), .A2(new_n759), .B1(new_n738), .B2(G294), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G326), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n752), .B1(new_n753), .B2(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n746), .A2(new_n754), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT90), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n726), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n729), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n725), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n659), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n713), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(G396));
  INV_X1    g0574(.A(KEYINPUT96), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n430), .A2(new_n432), .A3(new_n656), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n645), .B1(new_n638), .B2(new_n639), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n635), .B1(new_n684), .B2(KEYINPUT26), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(KEYINPUT95), .B(new_n776), .C1(new_n779), .C2(new_n637), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT95), .ZN(new_n781));
  INV_X1    g0581(.A(new_n776), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n647), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n421), .A2(new_n656), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n623), .B1(new_n785), .B2(new_n432), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n430), .A2(new_n655), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n647), .B2(new_n656), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n702), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n775), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n711), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  OAI211_X1 g0593(.A(KEYINPUT96), .B(new_n702), .C1(new_n784), .C2(new_n789), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n768), .A2(new_n724), .ZN(new_n796));
  INV_X1    g0596(.A(new_n738), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n254), .B1(new_n214), .B2(new_n797), .C1(new_n745), .C2(new_n466), .ZN(new_n798));
  INV_X1    g0598(.A(new_n731), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G311), .A2(new_n759), .B1(new_n799), .B2(G87), .ZN(new_n800));
  INV_X1    g0600(.A(new_n741), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n800), .B1(new_n423), .B2(new_n733), .C1(new_n801), .C2(new_n588), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT91), .B(G283), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n752), .B1(new_n753), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n798), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n744), .A2(G143), .B1(new_n741), .B2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n753), .ZN(new_n809));
  INV_X1    g0609(.A(new_n752), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G137), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n257), .B1(new_n747), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT92), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n731), .A2(new_n203), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n797), .A2(new_n202), .B1(new_n733), .B2(new_n207), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT93), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n806), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n714), .B1(G77), .B2(new_n796), .C1(new_n820), .C2(new_n768), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT94), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n724), .C2(new_n788), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n795), .A2(new_n825), .ZN(G384));
  NAND2_X1  g0626(.A1(new_n495), .A2(new_n500), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT35), .ZN(new_n828));
  OAI211_X1 g0628(.A(G116), .B(new_n225), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT36), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n222), .A2(G77), .A3(new_n362), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n207), .A2(G68), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n274), .B(G13), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n351), .A2(new_n655), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n322), .A2(G179), .A3(new_n324), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n325), .B2(new_n326), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n327), .B2(new_n332), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n355), .B(new_n836), .C1(new_n839), .C2(new_n350), .ZN(new_n840));
  INV_X1    g0640(.A(new_n355), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n351), .B(new_n655), .C1(new_n337), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AND4_X1   g0643(.A1(KEYINPUT40), .A2(new_n701), .A3(new_n843), .A4(new_n788), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n409), .A2(new_n653), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT37), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT97), .B1(new_n409), .B2(new_n410), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT97), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n379), .A2(new_n849), .A3(new_n393), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT37), .B1(new_n409), .B2(new_n403), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n653), .B(KEYINPUT98), .Z(new_n852));
  NAND2_X1  g0652(.A1(new_n379), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n848), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n846), .B1(new_n621), .B2(new_n625), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT38), .ZN(new_n857));
  INV_X1    g0657(.A(new_n852), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n409), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n845), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n854), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n413), .A2(new_n859), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT99), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT38), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT99), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n854), .A2(new_n860), .B1(new_n413), .B2(new_n859), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n865), .B(new_n866), .C1(KEYINPUT38), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n844), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n855), .B2(new_n856), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n857), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n701), .A2(new_n843), .A3(new_n788), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT100), .ZN(new_n876));
  INV_X1    g0676(.A(new_n701), .ZN(new_n877));
  OR3_X1    g0677(.A1(new_n876), .A2(new_n628), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n628), .B2(new_n877), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(G330), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n622), .A2(new_n852), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n857), .A2(new_n871), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n865), .B1(new_n867), .B2(KEYINPUT38), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n352), .A2(new_n655), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n787), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n780), .B2(new_n783), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n843), .C1(new_n857), .C2(new_n871), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n688), .A2(new_n704), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n434), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n627), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n891), .B(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n880), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT101), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n897), .B1(new_n274), .B2(new_n708), .C1(new_n895), .C2(new_n880), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(KEYINPUT101), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n835), .B1(new_n898), .B2(new_n899), .ZN(G367));
  NAND2_X1  g0700(.A1(new_n510), .A2(new_n655), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n546), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n643), .A2(new_n540), .A3(new_n655), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n663), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n656), .B1(new_n904), .B2(new_n638), .ZN(new_n905));
  OR3_X1    g0705(.A1(new_n635), .A2(new_n583), .A3(new_n656), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n586), .B(new_n635), .C1(new_n583), .C2(new_n656), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n902), .A2(new_n903), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n668), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT42), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT42), .B1(new_n910), .B2(new_n668), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n905), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n917), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n913), .A2(new_n914), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n920), .A2(new_n905), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n908), .B(KEYINPUT43), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n918), .A2(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n661), .A2(new_n910), .A3(new_n666), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n675), .B(KEYINPUT41), .Z(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT44), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(new_n929), .C1(new_n910), .C2(new_n670), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n902), .A2(new_n903), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n630), .A2(new_n655), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n490), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n632), .B2(new_n655), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(new_n929), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT45), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n931), .B2(new_n934), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n910), .A2(new_n670), .A3(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n938), .A2(new_n942), .A3(new_n667), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n667), .B1(new_n938), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n933), .B1(new_n666), .B2(new_n932), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n660), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n705), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT105), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT105), .B1(new_n705), .B2(new_n947), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n945), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n927), .B1(new_n952), .B2(new_n706), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n925), .B(new_n926), .C1(new_n953), .C2(new_n710), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n727), .B1(new_n227), .B2(new_n417), .C1(new_n719), .C2(new_n238), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n714), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n804), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n741), .A2(new_n957), .B1(G317), .B2(new_n759), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n799), .A2(G97), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(G311), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n466), .B2(new_n753), .C1(new_n961), .C2(new_n752), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n254), .B1(new_n797), .B2(new_n423), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n733), .A2(new_n588), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n963), .B1(KEYINPUT46), .B2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(KEYINPUT46), .B2(new_n964), .C1(new_n745), .C2(new_n803), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n797), .A2(new_n203), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G137), .B2(new_n759), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n741), .A2(G50), .B1(G58), .B2(new_n734), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n808), .C2(new_n745), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n257), .B1(new_n731), .B2(new_n415), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT106), .Z(new_n972));
  INV_X1    g0772(.A(G143), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n973), .B2(new_n752), .C1(new_n748), .C2(new_n753), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n962), .A2(new_n966), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n956), .B1(new_n771), .B2(new_n908), .C1(new_n976), .C2(new_n768), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n954), .A2(new_n977), .ZN(G387));
  AOI22_X1  g0778(.A1(new_n744), .A2(G317), .B1(new_n741), .B2(G303), .ZN(new_n979));
  XNOR2_X1  g0779(.A(KEYINPUT108), .B(G322), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n979), .B1(new_n961), .B2(new_n753), .C1(new_n752), .C2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT48), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G294), .A2(new_n734), .B1(new_n738), .B2(new_n957), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT109), .Z(new_n987));
  AND2_X1   g0787(.A1(new_n987), .A2(KEYINPUT49), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(KEYINPUT49), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n254), .B1(new_n731), .B2(new_n588), .C1(new_n762), .C2(new_n747), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n257), .B(new_n959), .C1(new_n745), .C2(new_n207), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n747), .A2(new_n808), .B1(new_n733), .B2(new_n415), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n738), .A2(new_n418), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n801), .B2(new_n203), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n810), .A2(G159), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT107), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(new_n286), .C2(new_n753), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n768), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n666), .A2(new_n771), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n235), .A2(new_n266), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n719), .B1(new_n673), .B2(new_n715), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n1005));
  AOI21_X1  g0805(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n673), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1003), .A2(new_n1007), .B1(new_n423), .B2(new_n674), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n714), .B1(new_n1008), .B2(new_n728), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1000), .A2(new_n1001), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n947), .A2(new_n709), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n676), .B1(new_n950), .B2(new_n951), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT110), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n705), .A2(new_n947), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT111), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1012), .B1(new_n1016), .B2(new_n1019), .ZN(G393));
  NAND2_X1  g0820(.A1(new_n945), .A2(new_n710), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n243), .A2(new_n719), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n727), .B1(new_n214), .B2(new_n227), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n714), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n747), .A2(new_n980), .B1(new_n733), .B2(new_n804), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1025), .A2(new_n257), .A3(new_n732), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT113), .Z(new_n1027));
  AOI22_X1  g0827(.A1(new_n741), .A2(G294), .B1(G116), .B2(new_n738), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n803), .C2(new_n753), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n810), .A2(G317), .B1(new_n744), .B2(G311), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT52), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n753), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(G50), .B1(new_n287), .B2(new_n741), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n738), .A2(G77), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n203), .B2(new_n733), .C1(new_n973), .C2(new_n747), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n254), .B(new_n1036), .C1(G87), .C2(new_n799), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n810), .A2(G150), .B1(new_n744), .B2(G159), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1029), .A2(new_n1031), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1024), .B1(new_n1042), .B2(new_n726), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n910), .B2(new_n771), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n952), .A2(new_n675), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1021), .B(new_n1044), .C1(new_n1045), .C2(new_n1046), .ZN(G390));
  OAI21_X1  g0847(.A(new_n714), .B1(new_n287), .B2(new_n796), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n257), .B(new_n735), .C1(new_n744), .C2(G116), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n816), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n741), .A2(G97), .B1(G294), .B2(new_n759), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1035), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n423), .A2(new_n753), .B1(new_n752), .B2(new_n755), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1032), .A2(G137), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n810), .A2(G128), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n759), .A2(G125), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(KEYINPUT54), .B(G143), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n741), .A2(new_n1058), .B1(G50), .B2(new_n799), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n254), .B1(new_n738), .B2(G159), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n733), .A2(new_n808), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(new_n745), .C2(new_n813), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1052), .A2(new_n1053), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1048), .B1(new_n1066), .B2(new_n726), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n885), .B2(new_n724), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n888), .B1(new_n687), .B2(new_n786), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n843), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n886), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n864), .A4(new_n868), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n886), .B1(new_n889), .B2(new_n843), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n885), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n701), .A2(new_n788), .A3(G330), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n843), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1072), .B(new_n1079), .C1(new_n1073), .C2(new_n885), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1068), .B1(new_n1081), .B2(new_n709), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n434), .A2(new_n791), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n893), .A2(new_n627), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OR3_X1    g0886(.A1(new_n1086), .A2(new_n1077), .A3(new_n1069), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n889), .B1(new_n1086), .B2(new_n1077), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1078), .A2(new_n1080), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1089), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n676), .B1(new_n1081), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1082), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G378));
  NAND3_X1  g0894(.A1(new_n869), .A2(new_n874), .A3(G330), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n293), .A2(new_n653), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n308), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n308), .A2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1095), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1107), .A2(new_n869), .A3(G330), .A4(new_n874), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n891), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1106), .A2(new_n887), .A3(new_n1108), .A4(new_n890), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n710), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n711), .B1(G50), .B2(new_n796), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n254), .A2(new_n265), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1115), .B(new_n967), .C1(new_n744), .C2(G107), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G97), .A2(new_n1032), .B1(new_n810), .B2(G116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n747), .A2(new_n755), .B1(new_n733), .B2(new_n415), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n741), .A2(new_n418), .B1(G58), .B2(new_n799), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT58), .ZN(new_n1122));
  AOI21_X1  g0922(.A(G50), .B1(new_n288), .B2(new_n265), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1121), .A2(new_n1122), .B1(new_n1115), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1125), .A2(new_n752), .B1(new_n753), .B2(new_n813), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n741), .A2(G137), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n734), .A2(new_n1058), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n738), .A2(G150), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1126), .B(new_n1130), .C1(G128), .C2(new_n744), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n288), .B(new_n265), .C1(new_n731), .C2(new_n748), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G124), .B2(new_n759), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT59), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1124), .B1(new_n1122), .B2(new_n1121), .C1(new_n1133), .C2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1114), .B1(new_n1138), .B2(new_n726), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1107), .B2(new_n724), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT115), .Z(new_n1141));
  NAND2_X1  g0941(.A1(new_n1113), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1084), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1090), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT116), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT116), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1145), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1090), .A2(new_n1144), .B1(new_n1111), .B2(new_n1110), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n675), .B1(new_n1153), .B2(KEYINPUT57), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1143), .B1(new_n1152), .B2(new_n1154), .ZN(G375));
  NAND2_X1  g0955(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n710), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n714), .B1(G68), .B2(new_n796), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G128), .A2(new_n759), .B1(new_n738), .B2(G50), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n748), .B2(new_n733), .C1(new_n801), .C2(new_n808), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G137), .B2(new_n744), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n257), .B1(new_n731), .B2(new_n202), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT118), .Z(new_n1163));
  AOI22_X1  g0963(.A1(G132), .A2(new_n810), .B1(new_n1032), .B2(new_n1058), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n810), .A2(G294), .B1(G107), .B2(new_n741), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n588), .B2(new_n753), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT117), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n254), .B1(new_n415), .B2(new_n731), .C1(new_n745), .C2(new_n755), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n994), .B1(new_n214), .B2(new_n733), .C1(new_n803), .C2(new_n747), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1158), .B1(new_n1172), .B2(new_n726), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n843), .B2(new_n724), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1157), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1156), .A2(new_n1144), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1089), .A2(new_n927), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(G381));
  AND2_X1   g0979(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1154), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1142), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1093), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1012), .B(new_n773), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1184));
  OR3_X1    g0984(.A1(G381), .A2(G384), .A3(G390), .ZN(new_n1185));
  OR4_X1    g0985(.A1(G387), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(G407));
  OAI211_X1 g0986(.A(G407), .B(G213), .C1(G343), .C2(new_n1183), .ZN(G409));
  INV_X1    g0987(.A(G384), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT119), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT60), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1089), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n1177), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1087), .A2(new_n1088), .A3(new_n1084), .A4(KEYINPUT60), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n675), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1176), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT119), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(G384), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1189), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n654), .A2(G213), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n1197), .A3(new_n1189), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(G2897), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(G2897), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1202), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n1198), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT121), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G378), .B(new_n1143), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1153), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1113), .B(new_n1140), .C1(new_n1211), .C2(new_n927), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1093), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1209), .B1(new_n1214), .B2(new_n1200), .ZN(new_n1215));
  AOI211_X1 g1015(.A(KEYINPUT121), .B(new_n1201), .C1(new_n1210), .C2(new_n1213), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1208), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT122), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(KEYINPUT122), .B(new_n1208), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1201), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(KEYINPUT63), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1184), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n950), .A2(new_n951), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n675), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT110), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n773), .B1(new_n1229), .B2(new_n1012), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1225), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT123), .B1(new_n1233), .B2(new_n1184), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G390), .B1(new_n954), .B2(new_n977), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n954), .A2(new_n977), .A3(G390), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(KEYINPUT124), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT124), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n954), .A2(new_n1241), .A3(new_n977), .A4(G390), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1235), .A2(new_n1236), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1231), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(KEYINPUT123), .A3(new_n1184), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n954), .A2(new_n977), .A3(G390), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1247), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT125), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1239), .B(new_n1238), .C1(new_n1232), .C2(new_n1234), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1243), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1224), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  AND4_X1   g1053(.A1(KEYINPUT120), .A2(new_n1214), .A3(new_n1200), .A4(new_n1223), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT120), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1221), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT127), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1251), .B(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1252), .B1(new_n1222), .B2(new_n1207), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT126), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n1252), .C1(new_n1222), .C2(new_n1207), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT120), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1222), .A2(KEYINPUT120), .A3(new_n1223), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT62), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1261), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1259), .A2(new_n1273), .ZN(G405));
  NOR2_X1   g1074(.A1(new_n1182), .A2(G378), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1210), .ZN(new_n1276));
  OR3_X1    g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1223), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1223), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1261), .B(new_n1279), .ZN(G402));
endmodule


