//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT88), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n211));
  INV_X1    g010(.A(G22gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G15gat), .ZN(new_n213));
  INV_X1    g012(.A(G15gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G22gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n209), .B1(new_n216), .B2(KEYINPUT91), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(G1gat), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI221_X1 g019(.A(new_n216), .B1(KEYINPUT91), .B2(new_n209), .C1(G1gat), .C2(new_n218), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n223), .A2(KEYINPUT89), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n226), .A2(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n229));
  INV_X1    g028(.A(G50gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G43gat), .ZN(new_n231));
  INV_X1    g030(.A(G43gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G50gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT15), .ZN(new_n234));
  NAND2_X1  g033(.A1(G29gat), .A2(G36gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n223), .ZN(new_n238));
  NOR3_X1   g037(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n239));
  OAI22_X1  g038(.A1(new_n237), .A2(KEYINPUT15), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI22_X1  g039(.A1(new_n229), .A2(new_n234), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n240), .A2(new_n236), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n224), .A2(new_n225), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n228), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n234), .B1(new_n248), .B2(new_n235), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n243), .B(new_n244), .C1(new_n245), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n241), .B2(new_n244), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n245), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n222), .A2(KEYINPUT92), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT92), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n220), .A2(new_n257), .A3(new_n221), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n208), .B(new_n242), .C1(new_n253), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n222), .B2(new_n241), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(new_n242), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n208), .B(KEYINPUT13), .Z(new_n265));
  AOI22_X1  g064(.A1(new_n260), .A2(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT90), .B1(new_n254), .B2(KEYINPUT17), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n250), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n256), .A2(new_n258), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(new_n255), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(KEYINPUT18), .A3(new_n208), .A4(new_n242), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n207), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n260), .A2(new_n261), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n271), .A3(new_n274), .A4(new_n207), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT94), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n266), .A2(KEYINPUT94), .A3(new_n271), .A4(new_n207), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  INV_X1    g079(.A(G113gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(G120gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT69), .B(G113gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(G120gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G127gat), .B(G134gat), .Z(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT1), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n284), .A2(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n293), .B2(new_n292), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n289), .A2(new_n291), .B1(new_n287), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT26), .ZN(new_n303));
  INV_X1    g102(.A(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n302), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G183gat), .B(G190gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n302), .A2(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n316), .C1(new_n304), .C2(new_n305), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n309), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(new_n309), .C1(new_n313), .C2(new_n317), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n317), .A2(new_n309), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n298), .A2(G183gat), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G190gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT24), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n328), .B2(new_n311), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n322), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n319), .B(new_n321), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n313), .B(KEYINPUT65), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT66), .B1(new_n333), .B2(new_n322), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n296), .B(new_n308), .C1(new_n332), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(KEYINPUT66), .A3(new_n322), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n330), .A2(new_n331), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n319), .A4(new_n321), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n340), .A2(KEYINPUT71), .A3(new_n296), .A4(new_n308), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n308), .B1(new_n332), .B2(new_n334), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n295), .A2(new_n287), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n286), .A2(new_n288), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n290), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n341), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n280), .B1(new_n350), .B2(KEYINPUT32), .ZN(new_n351));
  XOR2_X1   g150(.A(G71gat), .B(G99gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G15gat), .B(G43gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n347), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(KEYINPUT33), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n337), .A2(new_n346), .A3(new_n341), .A4(new_n348), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT34), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n350), .B(KEYINPUT32), .C1(new_n280), .C2(new_n356), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n358), .B2(new_n361), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT73), .A3(KEYINPUT36), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n361), .ZN(new_n366));
  INV_X1    g165(.A(new_n360), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n371));
  OR2_X1    g170(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G197gat), .B(G204gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT22), .ZN(new_n376));
  INV_X1    g175(.A(G211gat), .ZN(new_n377));
  INV_X1    g176(.A(G218gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G211gat), .B(G218gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT74), .ZN(new_n383));
  INV_X1    g182(.A(new_n381), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n380), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(G148gat), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G141gat), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT80), .B1(new_n392), .B2(G148gat), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n392), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT81), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n391), .A2(new_n394), .A3(new_n397), .A4(new_n393), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(KEYINPUT2), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n401), .A2(KEYINPUT78), .A3(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G141gat), .B(G148gat), .Z(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n407), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n388), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n405), .B1(new_n396), .B2(new_n398), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n412), .A2(new_n414), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT3), .B1(new_n385), .B2(new_n417), .ZN(new_n422));
  OAI211_X1 g221(.A(G228gat), .B(G233gat), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT84), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n383), .A2(new_n387), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT3), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(KEYINPUT29), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n415), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n408), .B1(new_n382), .B2(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n421), .B2(new_n408), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n435), .A2(new_n385), .B1(new_n421), .B2(new_n422), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n429), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n434), .A2(new_n212), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n212), .B1(new_n434), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g238(.A(G78gat), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n418), .A2(new_n423), .A3(KEYINPUT84), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n428), .B1(new_n427), .B2(new_n432), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G22gat), .ZN(new_n444));
  INV_X1    g243(.A(G78gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n434), .A2(new_n212), .A3(new_n437), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  INV_X1    g247(.A(G106gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n440), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n440), .B2(new_n447), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT75), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n342), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n340), .A2(KEYINPUT75), .A3(new_n308), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n417), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G226gat), .A2(G233gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT76), .B(new_n459), .C1(new_n340), .C2(new_n308), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  INV_X1    g261(.A(new_n459), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n342), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n388), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n457), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT75), .B1(new_n340), .B2(new_n308), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n342), .A2(new_n417), .A3(new_n459), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n382), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G8gat), .B(G36gat), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT77), .ZN(new_n474));
  XNOR2_X1  g273(.A(G64gat), .B(G92gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT30), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n479));
  NOR4_X1   g278(.A1(new_n466), .A2(new_n471), .A3(new_n479), .A4(new_n476), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n476), .B1(new_n466), .B2(new_n471), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT0), .ZN(new_n485));
  XNOR2_X1  g284(.A(G57gat), .B(G85gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  OAI21_X1  g286(.A(KEYINPUT3), .B1(new_n419), .B2(new_n420), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n416), .A2(new_n488), .A3(new_n345), .ZN(new_n489));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT4), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n430), .B2(new_n345), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n296), .A2(new_n421), .A3(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT83), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT83), .B1(new_n494), .B2(new_n495), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n430), .A2(new_n345), .A3(new_n493), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT4), .B1(new_n296), .B2(new_n421), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n490), .A4(new_n489), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n489), .A2(new_n494), .A3(new_n490), .A4(new_n495), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n421), .B(new_n345), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT5), .B1(new_n508), .B2(new_n490), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n487), .B(new_n499), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n487), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n503), .B2(new_n506), .ZN(new_n512));
  INV_X1    g311(.A(new_n499), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT6), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n454), .B1(new_n483), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n374), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n460), .A2(new_n465), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n425), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n469), .A2(new_n470), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n385), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n477), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n477), .B1(new_n472), .B2(new_n527), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n522), .A2(new_n425), .B1(new_n524), .B2(new_n385), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT37), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT38), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n523), .A2(new_n527), .A3(new_n525), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT37), .B1(new_n466), .B2(new_n471), .ZN(new_n533));
  AND4_X1   g332(.A1(KEYINPUT38), .A2(new_n532), .A3(new_n476), .A4(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n521), .B(new_n526), .C1(new_n531), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n450), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n438), .A2(new_n439), .A3(G78gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n451), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n526), .A2(new_n479), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n472), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n481), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n489), .B1(new_n497), .B2(new_n498), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT39), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n545), .A3(G225gat), .A4(G233gat), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n508), .B2(new_n490), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n416), .A2(new_n345), .A3(new_n488), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT83), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n500), .B2(new_n501), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(new_n496), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n547), .B1(new_n551), .B2(new_n490), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n552), .A3(new_n487), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT40), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT40), .A4(new_n487), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n555), .A2(new_n514), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n540), .B1(new_n543), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT85), .B1(new_n535), .B2(new_n558), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n520), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n364), .A2(new_n540), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT86), .B1(new_n543), .B2(new_n521), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT35), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT86), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n483), .A2(new_n518), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n454), .A2(new_n370), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n279), .B1(new_n561), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(G57gat), .A2(G64gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G57gat), .A2(G64gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(KEYINPUT95), .A3(new_n577), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(G57gat), .A2(G64gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(G57gat), .A2(G64gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n575), .B(new_n584), .C1(new_n587), .C2(KEYINPUT95), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  AOI21_X1  g396(.A(new_n222), .B1(KEYINPUT21), .B2(new_n589), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G92gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT98), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(G99gat), .A3(G106gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT8), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n609), .B1(new_n608), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n268), .A2(new_n255), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n618), .A2(new_n254), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n621), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT97), .ZN(new_n626));
  XOR2_X1   g425(.A(G134gat), .B(G162gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n620), .B1(new_n619), .B2(new_n623), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n624), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n602), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n588), .B(new_n581), .C1(new_n615), .C2(new_n616), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n608), .A2(new_n614), .ZN(new_n637));
  INV_X1    g436(.A(new_n609), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n608), .A2(new_n614), .A3(new_n609), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n589), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n636), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n635), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n643), .A2(new_n635), .A3(new_n644), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n641), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  XOR2_X1   g452(.A(G120gat), .B(G148gat), .Z(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n644), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n646), .ZN(new_n663));
  AOI211_X1 g462(.A(KEYINPUT102), .B(new_n647), .C1(new_n643), .C2(new_n644), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(new_n653), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n634), .B(new_n660), .C1(new_n666), .C2(new_n658), .ZN(new_n667));
  INV_X1    g466(.A(new_n660), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n658), .B1(new_n665), .B2(new_n653), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n633), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n572), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n518), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n210), .ZN(G1324gat));
  INV_X1    g475(.A(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n543), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT16), .B(G8gat), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT104), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT104), .B(new_n682), .C1(new_n678), .C2(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(G8gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(new_n374), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n674), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n370), .A2(new_n214), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n674), .B2(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n454), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  XNOR2_X1  g491(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(new_n632), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n601), .A2(new_n671), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT105), .Z(new_n696));
  NAND2_X1  g495(.A1(new_n572), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(G29gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n521), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  OR3_X1    g499(.A1(new_n697), .A2(new_n693), .A3(new_n699), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT107), .B1(new_n565), .B2(new_n570), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT86), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n483), .B2(new_n518), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n454), .A2(new_n370), .A3(KEYINPUT87), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n566), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n364), .A2(new_n540), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n709), .A2(new_n518), .A3(new_n483), .A4(new_n567), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT85), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n543), .A2(new_n557), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n454), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n516), .A2(new_n517), .A3(new_n526), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n530), .A2(new_n476), .A3(new_n532), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT38), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n528), .A2(KEYINPUT38), .A3(new_n533), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n712), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n558), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n703), .A2(new_n711), .B1(new_n723), .B2(new_n520), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n702), .B1(new_n724), .B2(new_n632), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n561), .A2(new_n571), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(KEYINPUT44), .A3(new_n694), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n602), .A2(new_n279), .A3(new_n672), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n728), .A2(new_n521), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n700), .B(new_n701), .C1(new_n730), .C2(new_n698), .ZN(G1328gat));
  NAND2_X1  g530(.A1(new_n543), .A2(new_n225), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT46), .B1(new_n697), .B2(new_n732), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n697), .A2(KEYINPUT46), .A3(new_n732), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n728), .A2(new_n543), .A3(new_n729), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n225), .ZN(G1329gat));
  NOR2_X1   g535(.A1(new_n686), .A2(new_n232), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n725), .A2(new_n727), .A3(new_n729), .A4(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n232), .B1(new_n697), .B2(new_n364), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n540), .A3(new_n727), .A4(new_n729), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G50gat), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n572), .A2(new_n230), .A3(new_n540), .A4(new_n696), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(KEYINPUT48), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  NOR3_X1   g548(.A1(new_n565), .A2(KEYINPUT107), .A3(new_n570), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n708), .B1(new_n707), .B2(new_n710), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n561), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n279), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n633), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n672), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n518), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(G57gat), .Z(G1332gat));
  NAND2_X1  g558(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n752), .A2(new_n761), .A3(new_n756), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n483), .A2(KEYINPUT110), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n483), .A2(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n763), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n763), .A2(new_n766), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n767), .ZN(G1333gat));
  NAND4_X1  g570(.A1(new_n760), .A2(G71gat), .A3(new_n374), .A4(new_n762), .ZN(new_n772));
  INV_X1    g571(.A(G71gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n757), .B2(new_n364), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n772), .A2(KEYINPUT50), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT50), .B1(new_n772), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(G1334gat));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n540), .A3(new_n762), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g578(.A1(new_n601), .A2(new_n279), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT111), .Z(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n672), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n728), .A2(new_n521), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G85gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n752), .A2(new_n694), .A3(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n694), .A4(new_n781), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(KEYINPUT112), .A3(new_n786), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n518), .A2(G85gat), .A3(new_n671), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n784), .A2(new_n793), .ZN(G1336gat));
  INV_X1    g593(.A(new_n766), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(G92gat), .A3(new_n671), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n790), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n725), .A2(new_n727), .A3(new_n766), .A4(new_n782), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n787), .A2(new_n789), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n725), .A2(new_n543), .A3(new_n727), .A4(new_n782), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n802), .A2(new_n796), .B1(new_n803), .B2(G92gat), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n797), .A2(new_n801), .B1(new_n804), .B2(new_n800), .ZN(G1337gat));
  NAND3_X1  g604(.A1(new_n728), .A2(new_n374), .A3(new_n782), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n364), .A2(G99gat), .A3(new_n671), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n791), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1338gat));
  NOR3_X1   g609(.A1(new_n454), .A2(G106gat), .A3(new_n671), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n790), .A2(new_n791), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n725), .A2(new_n540), .A3(new_n727), .A4(new_n782), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n802), .A2(new_n811), .B1(new_n813), .B2(G106gat), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n812), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(G1339gat));
  NAND2_X1  g618(.A1(new_n754), .A2(new_n671), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n649), .A2(new_n645), .A3(new_n647), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n643), .A2(new_n647), .A3(new_n644), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT114), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826));
  INV_X1    g625(.A(new_n824), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n651), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n663), .B2(new_n664), .ZN(new_n831));
  INV_X1    g630(.A(new_n658), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT55), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n825), .B2(new_n828), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(new_n668), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n829), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(KEYINPUT115), .A3(new_n660), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n834), .B(new_n279), .C1(new_n838), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n277), .A2(new_n278), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n264), .A2(new_n265), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n208), .B1(new_n270), .B2(new_n242), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n206), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n671), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n834), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT115), .B1(new_n840), .B2(new_n660), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n835), .B(new_n668), .C1(new_n829), .C2(new_n839), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n753), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n672), .A2(new_n843), .A3(new_n846), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(new_n632), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n834), .B1(new_n838), .B2(new_n841), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n847), .A2(new_n632), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n821), .B1(new_n861), .B2(new_n601), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n518), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n709), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n766), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n283), .A3(new_n753), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n602), .B1(new_n857), .B2(new_n860), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT117), .B(new_n454), .C1(new_n867), .C2(new_n821), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n860), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n694), .B1(new_n871), .B2(KEYINPUT116), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(new_n856), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n820), .B1(new_n873), .B2(new_n602), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT117), .B1(new_n874), .B2(new_n454), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n795), .A2(new_n521), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n364), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n753), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n866), .B1(new_n879), .B2(new_n281), .ZN(G1340gat));
  AOI21_X1  g679(.A(G120gat), .B1(new_n865), .B2(new_n672), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n672), .A2(G120gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1341gat));
  NOR3_X1   g682(.A1(new_n864), .A2(new_n601), .A3(new_n766), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(G127gat), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n602), .A2(G127gat), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n886), .A2(new_n887), .B1(new_n878), .B2(new_n888), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n543), .A2(new_n632), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n863), .A2(new_n890), .A3(new_n709), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(KEYINPUT56), .Z(new_n893));
  AND2_X1   g692(.A1(new_n878), .A2(new_n694), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n890), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n374), .A2(new_n454), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n521), .A3(new_n896), .ZN(new_n897));
  NOR4_X1   g696(.A1(new_n897), .A2(G141gat), .A3(new_n279), .A4(new_n766), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n389), .A2(new_n390), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n877), .A2(new_n374), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n874), .B2(new_n540), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n540), .A2(KEYINPUT57), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n753), .A2(new_n660), .A3(new_n850), .A4(new_n840), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n694), .B1(new_n855), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n601), .B1(new_n870), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n905), .B2(new_n820), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n753), .B(new_n900), .C1(new_n901), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n898), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n907), .B2(new_n899), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  AOI221_X4 g711(.A(new_n898), .B1(new_n909), .B2(new_n912), .C1(new_n899), .C2(new_n907), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  NOR4_X1   g713(.A1(new_n897), .A2(G148gat), .A3(new_n671), .A4(new_n766), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT120), .Z(new_n916));
  INV_X1    g715(.A(G148gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n906), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n374), .A3(new_n877), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n917), .C1(new_n919), .C2(new_n672), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n862), .A2(new_n902), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n820), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n540), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n672), .B(new_n900), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n916), .B1(new_n920), .B2(new_n926), .ZN(G1345gat));
  NAND2_X1  g726(.A1(new_n602), .A2(G155gat), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT121), .ZN(new_n929));
  INV_X1    g728(.A(G155gat), .ZN(new_n930));
  INV_X1    g729(.A(new_n897), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n602), .A3(new_n795), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n919), .A2(new_n929), .B1(new_n930), .B2(new_n932), .ZN(G1346gat));
  INV_X1    g732(.A(G162gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n934), .A3(new_n891), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n919), .A2(new_n694), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n862), .A2(new_n521), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n795), .A2(new_n569), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n753), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n483), .A2(new_n521), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n370), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n862), .B2(new_n540), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n946), .B2(new_n868), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n279), .A2(new_n304), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(G1348gat));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n305), .A3(new_n672), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n876), .A2(new_n671), .A3(new_n944), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n305), .ZN(G1349gat));
  AOI21_X1  g751(.A(new_n326), .B1(new_n947), .B2(new_n602), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n602), .A2(new_n297), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n940), .B2(new_n955), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n953), .A2(KEYINPUT60), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT60), .B1(new_n953), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1350gat));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  INV_X1    g759(.A(new_n944), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n694), .B(new_n961), .C1(new_n869), .C2(new_n875), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n632), .A2(G190gat), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n874), .A2(new_n939), .A3(new_n518), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT61), .B1(new_n962), .B2(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n960), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n962), .A2(G190gat), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n972), .A2(KEYINPUT124), .A3(new_n963), .A4(new_n966), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n969), .A2(new_n973), .ZN(G1351gat));
  NAND3_X1  g773(.A1(new_n938), .A2(new_n766), .A3(new_n896), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n975), .A2(G197gat), .A3(new_n279), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT125), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n922), .A2(new_n924), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n686), .A2(new_n943), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n753), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G197gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n977), .A2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(new_n975), .ZN(new_n984));
  INV_X1    g783(.A(G204gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n984), .A2(new_n985), .A3(new_n672), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n978), .A2(new_n671), .A3(new_n979), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n987), .B(new_n988), .C1(new_n985), .C2(new_n989), .ZN(G1353gat));
  NAND3_X1  g789(.A1(new_n984), .A2(new_n377), .A3(new_n602), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n980), .A2(new_n602), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  AOI21_X1  g794(.A(G218gat), .B1(new_n984), .B2(new_n694), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n632), .A2(new_n378), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n996), .B1(new_n980), .B2(new_n998), .ZN(G1355gat));
endmodule


