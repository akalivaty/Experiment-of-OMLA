//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n476), .A2(G137), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n466), .B1(new_n464), .B2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n464), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n478), .A2(new_n482), .B1(G101), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n475), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n474), .A2(new_n482), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT3), .B1(new_n480), .B2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  OAI221_X1 g069(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  INV_X1    g072(.A(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(G2104), .ZN(new_n506));
  AND2_X1   g081(.A1(G126), .A2(G2105), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n501), .A2(new_n506), .B1(new_n482), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  INV_X1    g084(.A(G138), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n471), .A2(new_n472), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n511), .B2(new_n482), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n476), .A2(G138), .A3(new_n477), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n513), .A2(new_n468), .A3(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n508), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n517), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n518), .A2(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n524), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n528), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n518), .A2(new_n519), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n529), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n537), .A2(G89), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n525), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n531), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  XNOR2_X1  g127(.A(KEYINPUT73), .B(G81), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n525), .A2(new_n553), .B1(new_n520), .B2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n531), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n554), .B(KEYINPUT74), .C1(new_n531), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G860), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT76), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  INV_X1    g144(.A(G78), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n541), .A2(new_n569), .B1(new_n570), .B2(new_n517), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n573), .B1(new_n570), .B2(new_n517), .C1(new_n541), .C2(new_n569), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(G651), .A3(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT77), .B(new_n576), .C1(new_n538), .C2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n577), .B1(new_n579), .B2(KEYINPUT9), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n520), .B(new_n580), .C1(new_n579), .C2(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n525), .A2(G91), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n575), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n525), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n520), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n523), .B2(new_n524), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT80), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n525), .A2(G86), .B1(new_n520), .B2(G48), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n598), .B(G651), .C1(new_n591), .C2(new_n593), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n525), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT81), .Z(new_n604));
  AOI22_X1  g179(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n531), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n520), .A2(G54), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n531), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n525), .A2(G92), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT10), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n575), .A2(new_n583), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(G148));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n560), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n616), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g206(.A1(new_n498), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n634), .A2(new_n635), .B1(KEYINPUT84), .B2(G2100), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  OR3_X1    g212(.A1(new_n637), .A2(KEYINPUT84), .A3(G2100), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(KEYINPUT84), .B2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n493), .A2(G135), .ZN(new_n640));
  OAI221_X1 g215(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n487), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT85), .Z(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT15), .B(G2435), .Z(new_n648));
  XOR2_X1   g223(.A(KEYINPUT86), .B(G2438), .Z(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT87), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n650), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(G14), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT89), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n680), .A2(KEYINPUT20), .A3(new_n684), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n685), .B1(new_n684), .B2(new_n681), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G24), .ZN(new_n699));
  INV_X1    g274(.A(G290), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n493), .A2(G131), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n473), .A2(G107), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n488), .A2(G119), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(new_n704), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT91), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n698), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n698), .ZN(new_n719));
  INV_X1    g294(.A(G1971), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n601), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G6), .B2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n698), .A2(G23), .ZN(new_n728));
  INV_X1    g303(.A(G288), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n698), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT33), .B(G1976), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n721), .A2(new_n726), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n703), .B(new_n717), .C1(new_n733), .C2(KEYINPUT34), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(KEYINPUT34), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT36), .ZN(new_n736));
  NAND2_X1  g311(.A1(G164), .A2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G27), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n493), .A2(G141), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(G105), .B2(new_n483), .ZN(new_n746));
  INV_X1    g321(.A(G129), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n741), .B(new_n746), .C1(new_n747), .C2(new_n487), .ZN(new_n748));
  MUX2_X1   g323(.A(G32), .B(new_n748), .S(G29), .Z(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  AOI21_X1  g325(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n698), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n698), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1961), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT24), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G34), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n485), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n739), .B2(new_n738), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n704), .A2(G26), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n493), .A2(G140), .ZN(new_n766));
  OAI221_X1 g341(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n767));
  INV_X1    g342(.A(G128), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n487), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n765), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n698), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n698), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G1966), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n643), .B2(new_n704), .ZN(new_n781));
  INV_X1    g356(.A(new_n773), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n763), .A2(new_n771), .A3(new_n774), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n752), .A2(new_n755), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n704), .A2(G35), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT97), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n496), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT29), .ZN(new_n790));
  INV_X1    g365(.A(G2090), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(G115), .A2(G2104), .ZN(new_n793));
  INV_X1    g368(.A(G127), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n468), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(new_n474), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G139), .ZN(new_n801));
  INV_X1    g376(.A(new_n493), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(KEYINPUT95), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(KEYINPUT95), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G33), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(G2072), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(G2072), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n616), .A2(G16), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G4), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n810), .B1(G1348), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n786), .A2(new_n792), .A3(new_n809), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n698), .A2(G19), .ZN(new_n817));
  INV_X1    g392(.A(new_n560), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n698), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1341), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n790), .A2(new_n791), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n814), .A2(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n698), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G299), .B2(G16), .ZN(new_n827));
  INV_X1    g402(.A(G1956), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OR4_X1    g404(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n736), .A2(new_n816), .A3(new_n830), .ZN(G311));
  XOR2_X1   g406(.A(G311), .B(KEYINPUT99), .Z(G150));
  NAND2_X1  g407(.A1(new_n520), .A2(G55), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT100), .B(G93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n526), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n531), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n556), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n838), .B1(new_n558), .B2(new_n559), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n617), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n561), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n838), .A2(new_n561), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(G145));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n769), .B(new_n515), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n805), .B(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n748), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n712), .B(new_n634), .ZN(new_n856));
  OAI221_X1 g431(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n857));
  INV_X1    g432(.A(G130), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n487), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G142), .B2(new_n493), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n856), .B(new_n860), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n854), .A2(new_n748), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n855), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n855), .A2(new_n862), .ZN(new_n865));
  INV_X1    g440(.A(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n496), .B(new_n485), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n643), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n864), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n867), .A2(new_n863), .ZN(new_n873));
  OAI221_X1 g448(.A(new_n852), .B1(new_n871), .B2(new_n872), .C1(new_n870), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g450(.A1(new_n839), .A2(new_n627), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(G305), .ZN(new_n877));
  XNOR2_X1  g452(.A(G303), .B(G288), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT42), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n629), .B(new_n842), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n616), .A2(G299), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n621), .A2(new_n613), .A3(new_n615), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n882), .A2(KEYINPUT102), .A3(new_n883), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT102), .B1(new_n882), .B2(new_n883), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n887), .B1(new_n881), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n880), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n876), .B1(new_n892), .B2(new_n627), .ZN(G295));
  OAI21_X1  g468(.A(new_n876), .B1(new_n892), .B2(new_n627), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  AOI21_X1  g470(.A(G168), .B1(new_n548), .B2(new_n550), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n548), .A2(G168), .A3(new_n550), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n842), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n900), .A2(new_n896), .B1(new_n841), .B2(new_n840), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT103), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n842), .A2(new_n903), .A3(new_n897), .A4(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n882), .A2(new_n883), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n901), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n905), .A2(new_n906), .B1(new_n886), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n879), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n886), .A2(new_n904), .A3(new_n902), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n901), .B(new_n899), .C1(new_n888), .C2(new_n889), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n879), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n909), .A2(new_n914), .A3(new_n852), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT105), .ZN(new_n918));
  OAI211_X1 g493(.A(KEYINPUT104), .B(new_n852), .C1(new_n908), .C2(new_n879), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n919), .A2(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n852), .B1(new_n908), .B2(new_n879), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n916), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n895), .B1(new_n918), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n923), .A2(new_n916), .A3(new_n909), .A4(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT106), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n920), .A2(new_n928), .A3(new_n916), .A4(new_n923), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n916), .B1(new_n915), .B2(KEYINPUT107), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n909), .A2(new_n914), .A3(new_n852), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n895), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n930), .A2(new_n935), .A3(KEYINPUT108), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT108), .B1(new_n930), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n925), .B1(new_n936), .B2(new_n937), .ZN(G397));
  INV_X1    g513(.A(G8), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT4), .B1(new_n492), .B2(new_n513), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n465), .A2(new_n467), .A3(new_n509), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n511), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n943), .B2(new_n508), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n475), .A2(new_n484), .A3(G40), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n939), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1976), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n729), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n950));
  OAI21_X1  g525(.A(G1981), .B1(new_n596), .B2(new_n600), .ZN(new_n951));
  INV_X1    g526(.A(G1981), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n595), .A2(new_n952), .A3(new_n599), .A4(new_n597), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(KEYINPUT49), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT113), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(KEYINPUT112), .A3(new_n953), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT112), .B1(new_n951), .B2(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n947), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n950), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n954), .B(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n959), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n957), .A3(new_n956), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT114), .A4(new_n947), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n949), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n953), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n947), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n515), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT115), .B1(new_n972), .B2(new_n945), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n974), .B(new_n946), .C1(new_n944), .C2(new_n970), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n515), .A2(new_n970), .A3(new_n971), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n975), .A3(new_n791), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n511), .A2(new_n482), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n978), .A2(KEYINPUT4), .B1(new_n511), .B2(new_n941), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n501), .A2(new_n506), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n482), .A2(new_n507), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n971), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n945), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n944), .A2(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n720), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n977), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n977), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(G8), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G166), .B2(new_n939), .ZN(new_n995));
  NAND3_X1  g570(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n946), .B1(new_n944), .B2(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n983), .A2(new_n984), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n999), .B(new_n783), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n945), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(new_n761), .A3(new_n976), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1966), .B1(new_n985), .B2(new_n986), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n999), .ZN(new_n1007));
  OAI211_X1 g582(.A(G8), .B(G168), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n946), .B1(new_n944), .B2(new_n970), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n976), .A2(new_n791), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1013), .A2(new_n1014), .B1(new_n987), .B2(new_n720), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT109), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1003), .A2(new_n1014), .A3(new_n791), .A4(new_n976), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n988), .A2(new_n1016), .A3(new_n1010), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n995), .A2(new_n1022), .A3(new_n996), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n995), .B2(new_n996), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n998), .A2(new_n1009), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n961), .A2(new_n966), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n947), .B1(new_n948), .B2(G288), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n729), .A2(G1976), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1028), .A2(KEYINPUT52), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(KEYINPUT52), .B2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n969), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT63), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1008), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1027), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT118), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n988), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT110), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(G8), .A4(new_n1019), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n997), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1034), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1033), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G168), .A2(new_n939), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n515), .A2(new_n970), .A3(new_n971), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1049), .A2(new_n972), .A3(new_n945), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1006), .A2(new_n999), .B1(new_n1050), .B2(new_n761), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT117), .B1(new_n1052), .B2(G1966), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1053), .A3(KEYINPUT123), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1046), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n939), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1046), .B1(new_n1056), .B2(KEYINPUT124), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1058), .B(new_n939), .C1(new_n1048), .C2(new_n1054), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT51), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1046), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1055), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n1065));
  NAND3_X1  g640(.A1(G299), .A2(new_n1065), .A3(KEYINPUT57), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(KEYINPUT57), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(KEYINPUT57), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n575), .A2(new_n583), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n828), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1052), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1348), .B1(new_n1003), .B2(new_n976), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n944), .A2(new_n946), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G2067), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n617), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1071), .A2(new_n828), .B1(new_n1052), .B2(new_n1073), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT120), .B1(new_n1082), .B2(new_n1070), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1070), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1072), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1075), .ZN(new_n1089));
  INV_X1    g664(.A(G1996), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1052), .A2(KEYINPUT121), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n987), .B2(G1996), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1079), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n818), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1096), .A2(KEYINPUT122), .A3(KEYINPUT59), .A4(new_n818), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1079), .A2(G2067), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n616), .C1(G1348), .C2(new_n1050), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1081), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1103), .A2(KEYINPUT60), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1089), .A2(new_n1099), .A3(new_n1100), .A4(new_n1106), .ZN(new_n1107));
  AND4_X1   g682(.A1(KEYINPUT61), .A2(new_n1077), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1086), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1039), .A2(new_n1025), .A3(G8), .A4(new_n1019), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1027), .A2(new_n1110), .A3(new_n1031), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n987), .B2(G2078), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1011), .B2(new_n1049), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT53), .A4(new_n739), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1117), .B2(KEYINPUT125), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(G301), .B(KEYINPUT54), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1121), .A2(new_n1122), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n993), .A2(new_n997), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1111), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1109), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1044), .B1(new_n1064), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1044), .B(KEYINPUT126), .C1(new_n1064), .C2(new_n1127), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1063), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1005), .A2(new_n1007), .A3(new_n1047), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT123), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1058), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1056), .A2(KEYINPUT124), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1046), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(new_n1138), .B2(KEYINPUT51), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT62), .B1(new_n1139), .B2(new_n1055), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1055), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1111), .A2(new_n1125), .A3(G301), .A4(new_n1121), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1130), .A2(new_n1131), .A3(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n944), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n713), .A2(new_n715), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n769), .B(G2067), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n748), .B(G1996), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n713), .A2(new_n715), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1149), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(G290), .B(G1986), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1147), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1148), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1152), .A2(new_n713), .A3(new_n715), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n769), .A2(G2067), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1148), .B1(new_n1150), .B2(new_n748), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1158), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT46), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1148), .B2(new_n1090), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1162), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT47), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n1154), .A2(new_n1148), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n700), .A2(new_n702), .A3(new_n1148), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1161), .B(new_n1167), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(new_n918), .A2(new_n924), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n461), .A2(G227), .ZN(new_n1175));
  OAI211_X1 g749(.A(KEYINPUT127), .B(new_n1175), .C1(new_n661), .C2(new_n662), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n661), .B2(new_n662), .ZN(new_n1177));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g753(.A1(new_n874), .A2(new_n696), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1174), .A2(new_n1180), .ZN(G308));
  OR2_X1    g755(.A1(new_n1174), .A2(new_n1180), .ZN(G225));
endmodule


