//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(KEYINPUT80), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n191), .A2(new_n192), .A3(KEYINPUT80), .A4(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n190), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT0), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n202), .B1(new_n207), .B2(new_n205), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n189), .A2(new_n197), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n192), .A2(KEYINPUT80), .A3(G104), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT3), .B1(new_n211), .B2(G107), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n190), .B(new_n196), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT4), .B(new_n213), .C1(new_n197), .C2(KEYINPUT81), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  AOI211_X1 g029(.A(new_n215), .B(new_n190), .C1(new_n195), .C2(new_n196), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n209), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(G137), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(G137), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G134), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n225), .B2(new_n218), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n223), .A2(new_n226), .A3(G131), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n224), .A2(G134), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT64), .B1(new_n224), .B2(G134), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(new_n219), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n218), .B1(new_n220), .B2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n228), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n227), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n223), .B2(new_n226), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n233), .A2(new_n228), .A3(new_n221), .A4(new_n222), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT10), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n192), .A2(KEYINPUT82), .A3(G104), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n192), .A2(G104), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT82), .B1(new_n192), .B2(G104), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n213), .B1(new_n245), .B2(new_n190), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n202), .A2(new_n247), .A3(G128), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n199), .B(new_n201), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n241), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n244), .A2(new_n243), .ZN(new_n253));
  OAI21_X1  g067(.A(G101), .B1(new_n253), .B2(new_n242), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n252), .A2(KEYINPUT10), .A3(new_n213), .A4(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n217), .A2(new_n240), .A3(new_n251), .A4(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n251), .A2(new_n255), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n259), .A2(KEYINPUT83), .A3(new_n217), .A4(new_n240), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n252), .A2(new_n213), .A3(new_n254), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n246), .A2(new_n250), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n236), .A2(new_n238), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(KEYINPUT12), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(new_n264), .A3(new_n268), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G140), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G227), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n277), .B(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n261), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n259), .A2(new_n217), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n275), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n261), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n261), .A2(new_n276), .ZN(new_n286));
  INV_X1    g100(.A(new_n280), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n258), .B2(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n283), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n285), .B1(new_n291), .B2(new_n187), .ZN(new_n292));
  INV_X1    g106(.A(G475), .ZN(new_n293));
  NOR2_X1   g107(.A1(G237), .A2(G953), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n294), .A2(G143), .A3(G214), .ZN(new_n295));
  AOI21_X1  g109(.A(G143), .B1(new_n294), .B2(G214), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT17), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT88), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G125), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G140), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT16), .ZN(new_n304));
  OR3_X1    g118(.A1(new_n302), .A2(KEYINPUT16), .A3(G140), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n304), .A2(G146), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(G146), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n294), .A2(G214), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n200), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n294), .A2(G143), .A3(G214), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n228), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n297), .A2(new_n312), .A3(new_n298), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT17), .A4(G131), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n299), .A2(new_n308), .A3(new_n313), .A4(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(new_n198), .ZN(new_n320));
  AND4_X1   g134(.A1(new_n318), .A2(new_n301), .A3(new_n303), .A4(new_n198), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n320), .A2(new_n321), .B1(new_n198), .B2(new_n319), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n314), .A2(new_n323), .A3(KEYINPUT18), .A4(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(KEYINPUT18), .A3(G131), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n310), .A2(new_n311), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G113), .B(G122), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT87), .B(G104), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n317), .A2(new_n327), .A3(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n293), .B1(new_n335), .B2(new_n188), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G475), .A2(G902), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n297), .A2(new_n312), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT19), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n198), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n304), .A2(new_n305), .A3(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n304), .A2(new_n305), .A3(new_n346), .A4(G146), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n340), .A2(new_n343), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n327), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n332), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n339), .B1(new_n350), .B2(new_n334), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT20), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n337), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n356), .A2(new_n357), .A3(G953), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT89), .B1(new_n204), .B2(G143), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n200), .A3(G128), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n200), .A2(G128), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n220), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G116), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n367), .A2(G122), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(G122), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n192), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(G107), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT13), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT90), .A3(new_n365), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT13), .B1(new_n360), .B2(new_n362), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(new_n364), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n363), .A2(new_n374), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n373), .B1(new_n382), .B2(G134), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n363), .A2(new_n365), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G134), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n366), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n192), .B1(new_n368), .B2(KEYINPUT14), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n387), .A2(new_n370), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n370), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n359), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n364), .B1(new_n363), .B2(new_n374), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n380), .B1(new_n393), .B2(KEYINPUT90), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n220), .B1(new_n394), .B2(new_n379), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n392), .B(new_n358), .C1(new_n395), .C2(new_n373), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n188), .ZN(new_n398));
  INV_X1    g212(.A(G478), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT15), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n391), .B2(new_n396), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(KEYINPUT15), .B2(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G952), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G953), .ZN(new_n406));
  INV_X1    g220(.A(G234), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(new_n188), .B(new_n278), .C1(G234), .C2(G237), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(G898), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n355), .A2(new_n404), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G210), .B1(G237), .B2(G902), .ZN(new_n417));
  INV_X1    g231(.A(new_n246), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n367), .A2(G119), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT2), .B(G113), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT66), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G113), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT2), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G113), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G116), .B(G119), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT66), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n425), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n424), .A2(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n418), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n196), .B1(new_n210), .B2(new_n212), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT81), .B1(new_n439), .B2(G101), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n216), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n422), .A2(new_n423), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT66), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n431), .B1(new_n429), .B2(new_n430), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n197), .A2(new_n189), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n437), .B(new_n438), .C1(new_n442), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(G101), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n215), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n197), .A2(KEYINPUT81), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(KEYINPUT4), .A3(new_n452), .A4(new_n213), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n424), .A2(new_n432), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n454), .A2(new_n443), .B1(new_n189), .B2(new_n197), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n453), .A2(new_n455), .B1(new_n418), .B2(new_n436), .ZN(new_n456));
  INV_X1    g270(.A(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT85), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n449), .B(KEYINPUT6), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n437), .B1(new_n442), .B2(new_n448), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n460), .A2(KEYINPUT85), .A3(new_n461), .A4(new_n457), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n250), .A2(new_n302), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n206), .A2(G125), .A3(new_n208), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G224), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(G953), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n465), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n459), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n438), .B(KEYINPUT8), .Z(new_n470));
  NAND2_X1  g284(.A1(new_n434), .A2(new_n435), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n454), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n246), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n437), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(new_n466), .B2(G953), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n463), .A2(new_n464), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n480), .B2(new_n449), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n417), .B1(new_n469), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n481), .A3(new_n417), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n416), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n292), .A2(new_n414), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT91), .ZN(new_n488));
  INV_X1    g302(.A(new_n486), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n286), .A2(new_n287), .B1(new_n289), .B2(new_n283), .ZN(new_n490));
  OAI21_X1  g304(.A(G469), .B1(new_n490), .B2(G902), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n491), .B2(new_n285), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n414), .A4(new_n485), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT69), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G101), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n294), .A2(G210), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n497), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n225), .A2(new_n222), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G131), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n248), .A2(new_n249), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n504), .A2(new_n238), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n206), .A2(new_n208), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n275), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n446), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT28), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n235), .A2(new_n506), .A3(new_n239), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n504), .A2(new_n238), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n236), .A2(new_n238), .B1(new_n206), .B2(new_n208), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n446), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n501), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n506), .A2(new_n266), .B1(new_n504), .B2(new_n238), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT65), .B1(new_n519), .B2(KEYINPUT30), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n505), .C2(new_n514), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n446), .A4(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n501), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n513), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT31), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(new_n529), .A3(new_n513), .A4(new_n526), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n501), .C1(new_n509), .C2(new_n516), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n518), .A2(new_n528), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT71), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G472), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n507), .B2(new_n508), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT72), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n513), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n509), .B1(new_n543), .B2(KEYINPUT28), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n501), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OR3_X1    g361(.A1(new_n509), .A2(new_n516), .A3(new_n501), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n525), .A2(new_n513), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n501), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n538), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT32), .B1(new_n533), .B2(new_n535), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n537), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n204), .A2(G119), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT23), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n419), .A2(G128), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(G110), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n555), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT24), .B(G110), .Z(new_n567));
  OAI211_X1 g381(.A(new_n561), .B(KEYINPUT74), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n345), .A2(new_n347), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n320), .A2(new_n321), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT74), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n563), .B2(new_n565), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n560), .A2(G110), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n567), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n560), .A2(G110), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n577), .C1(new_n306), .C2(new_n307), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n278), .A2(G221), .A3(G234), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT77), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n575), .A2(new_n578), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n357), .B1(G234), .B2(new_n188), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  INV_X1    g406(.A(new_n587), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n584), .B1(new_n575), .B2(new_n578), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n592), .B(new_n188), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n589), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n588), .B2(new_n188), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT79), .B1(new_n554), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n533), .A2(new_n535), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT32), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n551), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n513), .B1(new_n541), .B2(KEYINPUT72), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n539), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT28), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n509), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n546), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n188), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G472), .B1(new_n603), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n602), .A2(new_n611), .A3(new_n536), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n613));
  INV_X1    g427(.A(new_n598), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n495), .B1(new_n599), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(new_n190), .ZN(G3));
  AOI211_X1 g431(.A(new_n489), .B(new_n598), .C1(new_n491), .C2(new_n285), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n533), .A2(new_n188), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(G472), .ZN(new_n621));
  AOI211_X1 g435(.A(KEYINPUT92), .B(new_n538), .C1(new_n533), .C2(new_n188), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n618), .B(new_n600), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n398), .A2(new_n625), .A3(new_n399), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT93), .B1(new_n402), .B2(G478), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n399), .A2(G902), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n397), .A2(KEYINPUT33), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n391), .B2(new_n396), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n630), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n629), .B1(new_n628), .B2(new_n634), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n355), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n413), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n485), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AOI21_X1  g458(.A(new_n336), .B1(new_n401), .B2(new_n403), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT95), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n354), .B1(new_n353), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n351), .B2(new_n352), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n352), .B2(new_n351), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n645), .A2(new_n639), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n648), .B(new_n354), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n653), .A2(KEYINPUT96), .A3(new_n639), .A4(new_n645), .ZN(new_n654));
  AND4_X1   g468(.A1(KEYINPUT97), .A2(new_n652), .A3(new_n485), .A4(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n469), .A2(new_n417), .A3(new_n481), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n415), .B1(new_n656), .B2(new_n482), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n650), .B2(new_n651), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT97), .B1(new_n658), .B2(new_n654), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n623), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n579), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n590), .ZN(new_n666));
  OAI211_X1 g480(.A(KEYINPUT98), .B(new_n666), .C1(new_n596), .C2(new_n597), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n188), .B1(new_n593), .B2(new_n594), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT25), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n595), .A3(new_n589), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT98), .B1(new_n671), .B2(new_n666), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n488), .A2(new_n494), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n600), .B1(new_n621), .B2(new_n622), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(new_n492), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n554), .A2(new_n657), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n410), .B1(new_n411), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n653), .A2(new_n645), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n673), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n537), .A2(new_n553), .ZN(new_n692));
  INV_X1    g506(.A(new_n549), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n501), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n188), .B1(new_n543), .B2(new_n526), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n691), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n691), .A2(new_n602), .A3(new_n536), .A4(new_n696), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n684), .B(KEYINPUT39), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n492), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n703), .A2(KEYINPUT40), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(KEYINPUT40), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n656), .A2(new_n482), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT38), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n353), .A2(new_n354), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n336), .ZN(new_n709));
  INV_X1    g523(.A(new_n404), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n415), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n674), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n701), .A2(new_n704), .A3(new_n705), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  AOI21_X1  g529(.A(new_n625), .B1(new_n398), .B2(new_n399), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n402), .A2(KEYINPUT93), .A3(G478), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n634), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n635), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n355), .A3(new_n685), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n673), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n682), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  NOR2_X1   g538(.A1(new_n281), .A2(new_n284), .ZN(new_n725));
  OAI21_X1  g539(.A(G469), .B1(new_n725), .B2(G902), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n285), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n489), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n641), .A2(new_n612), .A3(new_n728), .A4(new_n614), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NOR2_X1   g545(.A1(new_n554), .A2(new_n598), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n652), .A2(new_n485), .A3(new_n654), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT97), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n658), .A2(KEYINPUT97), .A3(new_n654), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n737), .A3(new_n728), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NAND4_X1  g553(.A1(new_n726), .A2(new_n485), .A3(new_n486), .A4(new_n285), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n673), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n414), .A3(new_n612), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  INV_X1    g557(.A(KEYINPUT100), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n608), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n606), .A2(KEYINPUT100), .A3(new_n607), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n526), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n528), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT101), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n746), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT100), .B1(new_n606), .B2(new_n607), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n501), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n528), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n754), .A3(new_n530), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n535), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n711), .A2(new_n485), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n727), .A2(new_n757), .A3(new_n413), .A4(new_n489), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n620), .A2(G472), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n756), .A2(new_n758), .A3(new_n614), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  INV_X1    g575(.A(new_n759), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n755), .B2(new_n535), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n709), .B(new_n684), .C1(new_n719), .C2(new_n635), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n741), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NOR3_X1   g580(.A1(new_n656), .A2(new_n482), .A3(new_n416), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n292), .A2(new_n486), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n764), .A3(KEYINPUT42), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT102), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n536), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n533), .A2(KEYINPUT102), .A3(KEYINPUT32), .A4(new_n535), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n602), .A3(new_n611), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n614), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT103), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT103), .A3(new_n614), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n769), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n612), .A2(new_n768), .A3(new_n614), .A4(new_n764), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n778), .A2(KEYINPUT104), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  INV_X1    g597(.A(new_n769), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n773), .A2(KEYINPUT103), .A3(new_n614), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT103), .B1(new_n773), .B2(new_n614), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n779), .A2(new_n780), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NAND4_X1  g605(.A1(new_n612), .A2(new_n768), .A3(new_n614), .A4(new_n686), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n720), .A2(new_n709), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT43), .B1(new_n709), .B2(KEYINPUT105), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n720), .B(new_n709), .C1(KEYINPUT105), .C2(KEYINPUT43), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT106), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n677), .A2(new_n673), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(KEYINPUT44), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n288), .A2(new_n290), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT45), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n802), .B(G469), .C1(new_n804), .C2(G902), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n803), .A2(KEYINPUT45), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n803), .A2(KEYINPUT45), .ZN(new_n807));
  OAI21_X1  g621(.A(G469), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(G469), .A2(G902), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(KEYINPUT46), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n810), .A3(new_n285), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n486), .A3(new_n702), .ZN(new_n812));
  INV_X1    g626(.A(new_n767), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n801), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT44), .B1(new_n799), .B2(new_n800), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n486), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n811), .A2(KEYINPUT47), .A3(new_n486), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n721), .A2(new_n614), .A3(new_n813), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n554), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G140), .ZN(G42));
  XNOR2_X1  g640(.A(new_n727), .B(KEYINPUT49), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n489), .A2(new_n416), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n707), .A2(new_n614), .A3(new_n828), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n701), .A2(new_n794), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT107), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n768), .A2(new_n674), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n762), .B(new_n721), .C1(new_n755), .C2(new_n535), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n336), .A2(new_n684), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n612), .A2(new_n710), .A3(new_n653), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n833), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n488), .A2(new_n494), .A3(new_n674), .ZN(new_n839));
  INV_X1    g653(.A(new_n640), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT108), .B1(new_n709), .B2(new_n404), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n720), .B2(new_n355), .ZN(new_n842));
  AOI211_X1 g656(.A(KEYINPUT108), .B(new_n709), .C1(new_n719), .C2(new_n635), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n839), .A2(new_n676), .B1(new_n844), .B2(new_n623), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n615), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n613), .B1(new_n612), .B2(new_n614), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n494), .B(new_n488), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n838), .A2(new_n846), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n681), .A2(new_n657), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n852), .B(new_n612), .C1(new_n722), .C2(new_n688), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n671), .A2(new_n666), .A3(new_n685), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n681), .A2(new_n757), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n697), .B2(new_n699), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n765), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n765), .A2(new_n856), .A3(KEYINPUT52), .A4(new_n853), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n776), .A2(new_n777), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n781), .B1(new_n863), .B2(new_n784), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n760), .A2(new_n738), .A3(new_n729), .A4(new_n742), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n614), .A2(new_n756), .A3(new_n758), .A4(new_n759), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n612), .A2(new_n728), .A3(new_n614), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n729), .B(new_n742), .C1(new_n660), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n787), .A2(new_n788), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT109), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n841), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n638), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT108), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n720), .A2(new_n876), .A3(new_n355), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n640), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n624), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n849), .A2(new_n678), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n763), .A2(new_n764), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n832), .B1(new_n881), .B2(new_n836), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n880), .A2(new_n865), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n859), .A2(new_n860), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n790), .A2(new_n883), .A3(new_n792), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI221_X4 g700(.A(KEYINPUT54), .B1(new_n861), .B2(new_n873), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n886), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT104), .B1(new_n778), .B2(new_n781), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n787), .A2(new_n783), .A3(new_n788), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n792), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n845), .A2(new_n616), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n870), .A2(new_n893), .A3(new_n838), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n884), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n888), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n409), .B1(new_n796), .B2(new_n797), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n763), .A2(new_n899), .A3(new_n614), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT110), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT50), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n728), .A2(new_n416), .A3(new_n707), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n726), .A2(new_n489), .A3(new_n285), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n821), .A2(new_n822), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n900), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n767), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n726), .A2(new_n486), .A3(new_n285), .A4(new_n767), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT111), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n614), .A2(new_n410), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n720), .A2(new_n355), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n700), .A3(new_n698), .A4(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n763), .A2(new_n899), .A3(new_n913), .A4(new_n674), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n906), .A2(new_n910), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT51), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n906), .A2(new_n910), .A3(new_n920), .A4(KEYINPUT51), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n916), .A2(new_n700), .A3(new_n698), .ZN(new_n925));
  OAI221_X1 g739(.A(new_n406), .B1(new_n740), .B2(new_n900), .C1(new_n925), .C2(new_n638), .ZN(new_n926));
  INV_X1    g740(.A(new_n863), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n899), .A2(new_n913), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n927), .A2(KEYINPUT48), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT48), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n923), .A2(new_n924), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT112), .B1(new_n898), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n895), .B2(new_n884), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n859), .A2(new_n860), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n935), .A2(new_n892), .A3(new_n886), .A4(new_n894), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT54), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n861), .A2(new_n873), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n889), .A2(new_n888), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(KEYINPUT112), .A3(new_n939), .A4(new_n932), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n405), .A2(new_n278), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n831), .B1(new_n933), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(KEYINPUT113), .B(new_n831), .C1(new_n933), .C2(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(G75));
  NAND2_X1  g761(.A1(new_n889), .A2(new_n938), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(G210), .A3(G902), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT56), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n459), .A2(new_n462), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT114), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT55), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n949), .A2(new_n950), .A3(new_n954), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n468), .B(KEYINPUT115), .Z(new_n958));
  AND3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n956), .B2(new_n957), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n278), .A2(G952), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT116), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n959), .A2(new_n960), .A3(new_n963), .ZN(G51));
  NAND2_X1  g778(.A1(new_n948), .A2(KEYINPUT54), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n939), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n809), .B(KEYINPUT57), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n725), .B(KEYINPUT117), .Z(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g784(.A1(new_n885), .A2(new_n886), .B1(new_n873), .B2(new_n861), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n188), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(G469), .A3(new_n804), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n961), .B1(new_n970), .B2(new_n973), .ZN(G54));
  NAND3_X1  g788(.A1(new_n972), .A2(KEYINPUT58), .A3(G475), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n350), .A2(new_n334), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n978), .A3(new_n961), .ZN(G60));
  OR2_X1    g793(.A1(new_n631), .A2(new_n633), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n937), .A2(new_n939), .ZN(new_n981));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT59), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n980), .A2(new_n983), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n963), .B(new_n984), .C1(new_n966), .C2(new_n985), .ZN(G63));
  INV_X1    g800(.A(KEYINPUT118), .ZN(new_n987));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT60), .Z(new_n989));
  NAND3_X1  g803(.A1(new_n948), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT118), .B1(new_n971), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n665), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT119), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT61), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n963), .B1(new_n993), .B2(new_n665), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n990), .A2(new_n992), .A3(new_n587), .A4(new_n586), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT119), .B1(new_n993), .B2(new_n665), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n998), .B(new_n997), .C1(new_n1001), .C2(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n412), .B2(new_n466), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT120), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n880), .A2(new_n865), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT121), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n953), .B1(G898), .B2(new_n278), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(G69));
  AOI21_X1  g824(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n765), .A2(new_n853), .ZN(new_n1012));
  OR3_X1    g826(.A1(new_n927), .A2(new_n812), .A3(new_n757), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n817), .A2(new_n825), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n278), .B1(new_n1014), .B2(new_n892), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n341), .A2(new_n342), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT122), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1016), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n683), .A2(G953), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT125), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1012), .A2(new_n714), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT123), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT62), .ZN(new_n1025));
  XOR2_X1   g839(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n813), .B(new_n703), .C1(new_n877), .C2(new_n875), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n848), .B2(new_n847), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1027), .A2(new_n817), .A3(new_n825), .A4(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1019), .A2(new_n278), .ZN(new_n1031));
  AOI22_X1  g845(.A1(new_n1015), .A2(new_n1022), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT126), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1011), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1033), .B1(new_n1032), .B2(KEYINPUT124), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  INV_X1    g852(.A(new_n1006), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1038), .B1(new_n1030), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n961), .B1(new_n1040), .B2(new_n694), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1014), .A2(new_n892), .A3(new_n1039), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1038), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n693), .B(new_n501), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1043), .B1(new_n550), .B2(new_n527), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT127), .Z(new_n1047));
  AOI21_X1  g861(.A(new_n1047), .B1(new_n889), .B2(new_n896), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1045), .A2(new_n1048), .ZN(G57));
endmodule


