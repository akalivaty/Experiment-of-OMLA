//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n602, new_n604, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n465), .B2(G101), .ZN(new_n466));
  AND4_X1   g041(.A1(new_n463), .A2(new_n459), .A3(G101), .A4(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n470), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AOI211_X1 g051(.A(KEYINPUT69), .B(new_n459), .C1(new_n473), .C2(new_n474), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n469), .B(new_n471), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n459), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n460), .A2(new_n461), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n459), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n480), .A2(new_n494), .A3(G138), .A4(new_n459), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n461), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n459), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n507), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n511), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT73), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n530));
  AND3_X1   g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n508), .A2(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(G89), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n510), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n518), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n521), .ZN(new_n541));
  OR3_X1    g116(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT75), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n539), .B2(new_n541), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n534), .A2(G81), .B1(new_n510), .B2(G43), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT76), .Z(new_n546));
  AOI22_X1  g121(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G860), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n510), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT5), .B(G543), .Z(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(G91), .B2(new_n534), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  OR2_X1    g142(.A1(new_n517), .A2(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(new_n510), .B2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n534), .A2(G87), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G288));
  AOI22_X1  g147(.A1(new_n534), .A2(G86), .B1(new_n510), .B2(G48), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n515), .B2(new_n516), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n510), .A2(G47), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n518), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n521), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(new_n534), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n560), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(G868), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g170(.A(new_n594), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G299), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G280));
  INV_X1    g175(.A(new_n593), .ZN(new_n601));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n549), .A2(new_n597), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n593), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n597), .B2(new_n605), .ZN(G323));
  XOR2_X1   g181(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  NAND2_X1  g183(.A1(new_n480), .A2(new_n465), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n488), .A2(G123), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  OR3_X1    g193(.A1(new_n459), .A2(KEYINPUT79), .A3(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT79), .B1(new_n459), .B2(G111), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n617), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n482), .B2(G135), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n612), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(G2096), .ZN(new_n627));
  NAND4_X1  g202(.A1(new_n613), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(G156));
  XOR2_X1   g203(.A(G1341), .B(G1348), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT82), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n632), .B(new_n638), .Z(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n642), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n647), .B(KEYINPUT17), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n650), .B(KEYINPUT84), .Z(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(new_n649), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n649), .B1(new_n654), .B2(new_n647), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI22_X1  g233(.A1(new_n658), .A2(KEYINPUT85), .B1(new_n654), .B2(new_n653), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(KEYINPUT85), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n664), .A2(new_n665), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(new_n666), .ZN(new_n674));
  MUX2_X1   g249(.A(new_n674), .B(new_n673), .S(new_n669), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n684), .A3(new_n682), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G23), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n571), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT33), .B(G1976), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n689), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1971), .ZN(new_n696));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G305), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  NOR3_X1   g276(.A1(new_n693), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n482), .A2(G131), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(G107), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G2105), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n488), .B2(G119), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n707), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G24), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n585), .B(KEYINPUT88), .Z(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1986), .Z(new_n721));
  NAND4_X1  g296(.A1(new_n704), .A2(new_n705), .A3(new_n717), .A4(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(KEYINPUT36), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n726), .B(new_n727), .C1(KEYINPUT36), .C2(new_n722), .ZN(new_n729));
  NOR2_X1   g304(.A1(G4), .A2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n601), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1348), .ZN(new_n732));
  NOR2_X1   g307(.A1(G164), .A2(new_n706), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G27), .B2(new_n706), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n623), .A2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n740));
  OR2_X1    g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  NAND2_X1  g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n732), .A2(new_n736), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n689), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  INV_X1    g322(.A(G299), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n689), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n706), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n745), .B(new_n751), .C1(G2084), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G171), .B2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT95), .Z(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(G168), .A2(G16), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(KEYINPUT94), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT94), .B2(new_n764), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1966), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n762), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n706), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n488), .A2(G128), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n482), .A2(G140), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n459), .A2(G116), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n774), .B(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2067), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  AOI22_X1  g358(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n459), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n482), .B2(G139), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT93), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G33), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT92), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n781), .B1(new_n791), .B2(G2072), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G35), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G162), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n794), .B(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n735), .B2(new_n734), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n792), .B(new_n799), .C1(G2072), .C2(new_n791), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n482), .A2(G141), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n488), .A2(G129), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT26), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n465), .A2(G105), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G32), .B(new_n806), .S(G29), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G19), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n546), .A2(new_n548), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G16), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n812), .A2(G1341), .B1(G2084), .B2(new_n756), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n813), .C1(G1341), .C2(new_n812), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n757), .A2(new_n769), .A3(new_n800), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n728), .A2(new_n729), .A3(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n510), .A2(G55), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n518), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n521), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n549), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n593), .A2(new_n602), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n828), .B(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n550), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n825), .A2(G860), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT98), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n490), .B(new_n623), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G160), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n500), .B2(new_n503), .ZN(new_n844));
  OAI221_X1 g419(.A(KEYINPUT99), .B1(new_n501), .B2(new_n502), .C1(new_n487), .C2(new_n497), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n496), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n496), .A2(new_n845), .A3(new_n844), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n778), .B(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n806), .Z(new_n852));
  INV_X1    g427(.A(new_n786), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n806), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n787), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n482), .A2(G142), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n459), .A2(G118), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n858), .B2(KEYINPUT101), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n859), .A2(new_n861), .B1(new_n488), .B2(G130), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n610), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n714), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n854), .A2(new_n856), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n854), .B2(new_n856), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(KEYINPUT102), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n854), .A2(new_n869), .A3(new_n865), .A4(new_n856), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n842), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n841), .B(KEYINPUT103), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n874), .B2(new_n867), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(G395));
  NAND2_X1  g453(.A1(new_n825), .A2(new_n597), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n827), .B(new_n605), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n593), .A2(new_n748), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n593), .A2(new_n748), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n881), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n890), .A2(new_n891), .B1(new_n881), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(new_n571), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n698), .B(new_n585), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n894), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n879), .B1(new_n899), .B2(new_n597), .ZN(G295));
  OAI21_X1  g475(.A(new_n879), .B1(new_n899), .B2(new_n597), .ZN(G331));
  XNOR2_X1  g476(.A(G171), .B(G168), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n827), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n827), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n885), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n897), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n893), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n893), .ZN(new_n911));
  INV_X1    g486(.A(new_n905), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n897), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n893), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n903), .A2(new_n904), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n916), .A2(KEYINPUT105), .A3(new_n906), .A4(new_n905), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n910), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n885), .A2(new_n891), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n888), .A2(new_n892), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n903), .A2(new_n904), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n905), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n897), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT43), .A2(new_n927), .A3(new_n910), .A4(new_n917), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n927), .A2(new_n910), .A3(new_n919), .A4(new_n917), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  XNOR2_X1  g510(.A(new_n778), .B(new_n780), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n806), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n716), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n939), .A2(new_n940), .B1(G2067), .B2(new_n778), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n847), .A2(new_n942), .A3(new_n849), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G40), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n478), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n937), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  INV_X1    g528(.A(new_n936), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n949), .B1(new_n954), .B2(new_n806), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n957));
  XOR2_X1   g532(.A(new_n713), .B(new_n716), .Z(new_n958));
  NOR2_X1   g533(.A1(new_n939), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n948), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n948), .A2(G1986), .A3(G290), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT48), .ZN(new_n963));
  OAI221_X1 g538(.A(new_n951), .B1(new_n956), .B2(new_n957), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n956), .B2(new_n957), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n480), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT69), .B1(new_n966), .B2(new_n459), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n475), .A2(new_n472), .A3(G2105), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(G40), .A3(new_n469), .A4(new_n471), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n846), .A2(new_n942), .ZN(new_n971));
  OAI21_X1  g546(.A(G8), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT111), .B(G8), .C1(new_n970), .C2(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n510), .A2(G48), .ZN(new_n977));
  INV_X1    g552(.A(G86), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n518), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n578), .ZN(new_n980));
  OAI21_X1  g555(.A(G1981), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n984));
  INV_X1    g559(.A(G1981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n573), .A2(new_n985), .A3(new_n578), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n573), .A2(KEYINPUT113), .A3(new_n985), .A4(new_n578), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n983), .A2(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT49), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n984), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n989), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n990), .A2(KEYINPUT115), .A3(KEYINPUT49), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n976), .B(new_n991), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(new_n571), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n994), .B(KEYINPUT116), .Z(new_n1002));
  OAI21_X1  g577(.A(new_n976), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n505), .A2(new_n942), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n496), .B2(new_n504), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT107), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n1008), .ZN(new_n1012));
  INV_X1    g587(.A(G2084), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .A4(new_n947), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n971), .A2(new_n944), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1007), .A2(KEYINPUT45), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n947), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1966), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  NOR2_X1   g596(.A1(G286), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n970), .B1(new_n944), .B2(new_n1004), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n942), .A4(new_n849), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1010), .A2(new_n1012), .A3(new_n796), .A4(new_n947), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1021), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n1030));
  OAI221_X1 g605(.A(G8), .B1(new_n1030), .B2(KEYINPUT55), .C1(new_n519), .C2(new_n522), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G166), .A2(new_n1021), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1020), .B(new_n1022), .C1(new_n1029), .C2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n571), .A2(G1976), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT112), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n947), .A2(new_n1011), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT111), .B1(new_n1038), .B2(G8), .ZN(new_n1039));
  INV_X1    g614(.A(new_n975), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1000), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n976), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n999), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT63), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1003), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n947), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1008), .B1(new_n846), .B2(new_n942), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n970), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1027), .B1(G2090), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1034), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(KEYINPUT63), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1034), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT109), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1028), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1971), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1071), .A2(KEYINPUT110), .A3(G8), .A4(new_n1065), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1045), .B1(new_n1061), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1047), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1014), .A2(new_n1019), .A3(G168), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(G168), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1080), .A3(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT62), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1034), .B1(new_n1055), .B2(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1045), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1079), .A2(new_n1081), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1004), .A2(new_n944), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1024), .A2(new_n947), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n735), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1010), .A2(new_n947), .A3(new_n1012), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1091), .B1(new_n761), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(G2078), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n947), .A2(new_n1015), .A3(new_n1016), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(G301), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1085), .A2(new_n1087), .A3(new_n1073), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1083), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1042), .A2(new_n1044), .A3(new_n999), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n1073), .A2(new_n1100), .A3(new_n1058), .A4(new_n1096), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT124), .B1(new_n1101), .B2(new_n1087), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1075), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1038), .A2(G2067), .ZN(new_n1104));
  INV_X1    g679(.A(G1348), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1092), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n593), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G299), .B(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1054), .A2(new_n750), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1024), .A2(new_n947), .A3(new_n1088), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n970), .A2(new_n1051), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1114), .A2(new_n1049), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1956), .B1(new_n1115), .B2(new_n1052), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1109), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1107), .A2(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(new_n601), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(KEYINPUT60), .B2(new_n1106), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n750), .B2(new_n1054), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1113), .B2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1038), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1024), .A2(new_n937), .A3(new_n947), .A4(new_n1088), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n811), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT119), .B(new_n549), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT59), .B(new_n1130), .C1(new_n1131), .C2(new_n1129), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1128), .A2(new_n811), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT118), .B(new_n1133), .C1(new_n1134), .C2(KEYINPUT119), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1124), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1110), .A2(KEYINPUT120), .A3(new_n1112), .A4(new_n1109), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1054), .A2(new_n750), .B1(new_n1089), .B2(new_n1111), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT61), .B1(new_n1141), .B2(new_n1109), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1136), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1121), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(KEYINPUT122), .B(new_n1136), .C1(new_n1143), .C2(new_n1146), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1118), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1152));
  XOR2_X1   g727(.A(G171), .B(KEYINPUT54), .Z(new_n1153));
  INV_X1    g728(.A(new_n945), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n946), .B1(new_n475), .B2(G2105), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n469), .A2(new_n471), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1156), .A2(KEYINPUT123), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(KEYINPUT123), .ZN(new_n1158));
  AND4_X1   g733(.A1(new_n1024), .A2(new_n1157), .A3(new_n1094), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1153), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1152), .A2(new_n1153), .B1(new_n1160), .B2(new_n1093), .ZN(new_n1161));
  AND4_X1   g736(.A1(new_n1073), .A2(new_n1085), .A3(new_n1082), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1103), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n585), .B(G1986), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n948), .B1(new_n959), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n965), .B1(new_n1163), .B2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g741(.A1(new_n871), .A2(new_n875), .ZN(new_n1168));
  INV_X1    g742(.A(new_n457), .ZN(new_n1169));
  OR3_X1    g743(.A1(new_n645), .A2(new_n1169), .A3(G227), .ZN(new_n1170));
  NOR2_X1   g744(.A1(G229), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1171), .A3(new_n932), .ZN(G225));
  INV_X1    g746(.A(G225), .ZN(G308));
endmodule


