//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n580, new_n581,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n642, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR3_X1   g034(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n453), .B2(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n458), .B1(new_n454), .B2(new_n459), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(KEYINPUT68), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n470), .A3(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n465), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n468), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT66), .B1(new_n480), .B2(new_n472), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(G2104), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n471), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n478), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(G113), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n471), .A2(new_n482), .A3(new_n483), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n483), .B1(new_n471), .B2(new_n482), .ZN(new_n492));
  OAI21_X1  g067(.A(G125), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n477), .B1(new_n490), .B2(new_n495), .ZN(G160));
  INV_X1    g071(.A(new_n476), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  OR2_X1    g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n500));
  INV_X1    g075(.A(G124), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n473), .A2(new_n475), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n498), .B(new_n500), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G162));
  NAND2_X1  g084(.A1(new_n465), .A2(G138), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n491), .B2(new_n492), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT68), .B1(new_n479), .B2(G2104), .ZN(new_n515));
  OAI211_X1 g090(.A(G126), .B(new_n475), .C1(new_n515), .C2(new_n480), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT71), .A2(G114), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT71), .A2(G114), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(G2104), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G2105), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n465), .A2(G102), .A3(G2104), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n475), .A4(new_n511), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n514), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G164));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .A3(G62), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n527), .A2(new_n529), .ZN(new_n534));
  INV_X1    g109(.A(G62), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n539), .A2(KEYINPUT6), .A3(G651), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT6), .B1(new_n539), .B2(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n534), .ZN(new_n543));
  OAI21_X1  g118(.A(G543), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(G88), .A2(new_n543), .B1(new_n545), .B2(G50), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n538), .A2(new_n546), .ZN(G303));
  INV_X1    g122(.A(G303), .ZN(G166));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n530), .B1(new_n541), .B2(new_n540), .ZN(new_n551));
  INV_X1    g126(.A(G89), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n545), .A2(G51), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(G286));
  INV_X1    g133(.A(G286), .ZN(G168));
  NAND2_X1  g134(.A1(G77), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G64), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n534), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n543), .A2(G90), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n545), .A2(G52), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G301));
  INV_X1    g143(.A(G301), .ZN(G171));
  NAND2_X1  g144(.A1(G68), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G56), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n534), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n545), .A2(G43), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n543), .A2(G81), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  AND3_X1   g152(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G36), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G188));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n545), .A2(new_n583), .A3(G53), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n545), .A2(new_n583), .A3(new_n586), .A4(G53), .ZN(new_n587));
  NAND2_X1  g162(.A1(G78), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G65), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n534), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n585), .A2(new_n587), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n543), .A2(KEYINPUT77), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n551), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G91), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(G299));
  NAND2_X1  g172(.A1(new_n545), .A2(G49), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n595), .B2(G87), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G288));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n592), .B2(new_n594), .ZN(new_n604));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n534), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n545), .A2(G48), .B1(new_n607), .B2(G651), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G305));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n534), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n545), .A2(G47), .B1(new_n614), .B2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n543), .A2(G85), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G651), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G66), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(G66), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n530), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n595), .A2(G92), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n595), .A2(KEYINPUT10), .A3(G92), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(G54), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n618), .B1(new_n635), .B2(G868), .ZN(G284));
  OAI21_X1  g211(.A(new_n618), .B1(new_n635), .B2(G868), .ZN(G321));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(G299), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G168), .B2(new_n638), .ZN(G297));
  XOR2_X1   g215(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n635), .B1(new_n642), .B2(G860), .ZN(G148));
  NAND2_X1  g218(.A1(new_n575), .A2(new_n638), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n634), .A2(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n481), .A2(new_n484), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(new_n467), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n497), .A2(G135), .ZN(new_n653));
  OAI21_X1  g228(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n656), .B(new_n657), .C1(G111), .C2(new_n465), .ZN(new_n658));
  INV_X1    g233(.A(G123), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n653), .B(new_n658), .C1(new_n659), .C2(new_n503), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2096), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n652), .A2(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT82), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XOR2_X1   g240(.A(G2443), .B(G2446), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1341), .B(G1348), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT15), .B(G2435), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(G2438), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2427), .B(G2430), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT14), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n669), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT84), .ZN(G401));
  XNOR2_X1  g253(.A(G2084), .B(G2090), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT85), .ZN(new_n680));
  XOR2_X1   g255(.A(G2067), .B(G2678), .Z(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT17), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT18), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(KEYINPUT18), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n688), .B(new_n690), .Z(G227));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT20), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n692), .A2(new_n693), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(KEYINPUT20), .ZN(new_n705));
  INV_X1    g280(.A(new_n694), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n698), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n702), .A2(new_n704), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1986), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1991), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n710), .B(new_n713), .ZN(G229));
  INV_X1    g289(.A(KEYINPUT97), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT23), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(G20), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n716), .B(new_n718), .C1(G299), .C2(G16), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n716), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1956), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n717), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1966), .ZN(new_n725));
  OR2_X1    g300(.A1(G5), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G301), .B2(new_n717), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n717), .A2(G19), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n576), .B2(new_n717), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1341), .ZN(new_n732));
  INV_X1    g307(.A(G28), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n660), .B2(new_n736), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G1341), .B2(new_n731), .ZN(new_n739));
  OR2_X1    g314(.A1(G29), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n497), .A2(G139), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n648), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n743), .C1(new_n744), .C2(new_n465), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n729), .A2(new_n732), .A3(new_n739), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n725), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT91), .B1(G4), .B2(G16), .ZN(new_n751));
  OR3_X1    g326(.A1(KEYINPUT91), .A2(G4), .A3(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n751), .B(new_n752), .C1(new_n634), .C2(new_n717), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n722), .A2(new_n750), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n736), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n736), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n758), .B(new_n760), .C1(G162), .C2(new_n736), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT96), .Z(new_n766));
  NOR2_X1   g341(.A1(G29), .A2(G32), .ZN(new_n767));
  INV_X1    g342(.A(new_n503), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n497), .A2(G141), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n467), .A2(G105), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n767), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT27), .B(G1996), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n779));
  INV_X1    g354(.A(G26), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G29), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(G29), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n497), .A2(G140), .ZN(new_n783));
  OR2_X1    g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n785));
  INV_X1    g360(.A(G128), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n785), .C1(new_n786), .C2(new_n503), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n782), .B1(new_n787), .B2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n781), .B1(new_n788), .B2(new_n779), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  OAI211_X1 g365(.A(G1961), .B(new_n726), .C1(G301), .C2(new_n717), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n746), .A2(new_n747), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n778), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G34), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT24), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT24), .ZN(new_n797));
  AOI21_X1  g372(.A(G29), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G160), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(G2084), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT92), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT94), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n794), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n762), .A2(new_n764), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n763), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n757), .A2(new_n766), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n736), .A2(G27), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n736), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2078), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n715), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n756), .A2(new_n806), .A3(new_n809), .ZN(new_n816));
  INV_X1    g391(.A(new_n814), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n816), .A2(KEYINPUT97), .A3(new_n817), .A4(new_n766), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n736), .A2(G25), .ZN(new_n820));
  OR2_X1    g395(.A1(G95), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n822));
  INV_X1    g397(.A(G131), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n476), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n768), .B2(G119), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n825), .B2(new_n736), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n717), .A2(G23), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n601), .B2(new_n717), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT33), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT33), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G1976), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n717), .A2(G6), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n610), .B2(new_n717), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT32), .B(G1981), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n831), .A2(G1976), .A3(new_n832), .ZN(new_n840));
  INV_X1    g415(.A(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT89), .B1(new_n841), .B2(G16), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n841), .A2(KEYINPUT89), .A3(G16), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(G166), .C2(new_n717), .ZN(new_n844));
  INV_X1    g419(.A(G1971), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n835), .A2(new_n839), .A3(new_n840), .A4(new_n846), .ZN(new_n847));
  AOI211_X1 g422(.A(new_n819), .B(new_n828), .C1(new_n847), .C2(KEYINPUT34), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n717), .A2(G24), .ZN(new_n849));
  INV_X1    g424(.A(G290), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n717), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT88), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G1986), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n848), .B(new_n853), .C1(KEYINPUT34), .C2(new_n847), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT36), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(KEYINPUT36), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n815), .A2(new_n818), .B1(new_n855), .B2(new_n856), .ZN(G311));
  NAND2_X1  g432(.A1(new_n815), .A2(new_n818), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(G150));
  NAND2_X1  g435(.A1(new_n635), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n619), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n543), .A2(G93), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n545), .A2(G55), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n865), .A2(KEYINPUT98), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT98), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n576), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n575), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT39), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n862), .B(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(G860), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT99), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(G860), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G145));
  XNOR2_X1  g454(.A(new_n508), .B(new_n660), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n799), .ZN(new_n881));
  INV_X1    g456(.A(new_n825), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n774), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n650), .B(new_n745), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n787), .B(new_n524), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n884), .A2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n883), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n768), .A2(G130), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n497), .A2(G142), .ZN(new_n894));
  OR2_X1    g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n889), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n889), .B2(new_n892), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n881), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n881), .B(KEYINPUT100), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n881), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n899), .A2(new_n900), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n881), .A2(new_n906), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g487(.A(new_n645), .B(new_n872), .ZN(new_n913));
  INV_X1    g488(.A(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n634), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n630), .A2(G299), .A3(new_n633), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n635), .A2(KEYINPUT102), .A3(G299), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n925), .B2(new_n913), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(G166), .B(new_n601), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(G305), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(G305), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n929), .A2(new_n850), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n850), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n935), .B(new_n921), .C1(new_n925), .C2(new_n913), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n927), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n927), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n869), .A2(new_n638), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(G295));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n940), .ZN(G331));
  AOI21_X1  g517(.A(G171), .B1(G286), .B2(KEYINPUT104), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n555), .A2(new_n945), .A3(new_n556), .A4(new_n557), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n870), .A2(new_n946), .A3(new_n871), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n870), .B2(new_n871), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n949), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n943), .B1(new_n951), .B2(new_n947), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n924), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n943), .A3(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n955), .A2(new_n956), .B1(new_n918), .B2(new_n919), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n933), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n924), .B2(new_n953), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n933), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT43), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n915), .A2(new_n917), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT41), .A4(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n950), .A2(new_n952), .A3(new_n922), .ZN(new_n967));
  INV_X1    g542(.A(new_n920), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n933), .B(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G37), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n969), .B(new_n970), .C1(new_n962), .C2(new_n933), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT44), .B1(new_n964), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n961), .B2(new_n963), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n510), .B1(new_n481), .B2(new_n484), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n522), .B(new_n523), .C1(new_n981), .C2(KEYINPUT4), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n465), .B1(new_n516), .B2(new_n519), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n477), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT67), .B1(new_n494), .B2(G2105), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n489), .B(new_n465), .C1(new_n493), .C2(new_n486), .ZN(new_n991));
  OAI211_X1 g566(.A(G40), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(G290), .A2(KEYINPUT106), .A3(G1986), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n996));
  INV_X1    g571(.A(G1986), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n850), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n850), .A2(new_n997), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT107), .Z(new_n1002));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n994), .B2(G1996), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n993), .A2(KEYINPUT108), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n775), .ZN(new_n1008));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n787), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1005), .B2(new_n775), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n993), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n882), .A2(new_n827), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n882), .A2(new_n827), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n993), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1008), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1002), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n984), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT109), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT50), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(G40), .A3(G160), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n728), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT124), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1020), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT109), .B1(new_n524), .B2(new_n980), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n524), .B2(new_n980), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n992), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT124), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n728), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n984), .A2(new_n986), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n524), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(G160), .A3(G40), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1036), .B1(new_n1039), .B2(G2078), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1036), .A2(G2078), .ZN(new_n1041));
  AND4_X1   g616(.A1(G40), .A2(new_n1038), .A3(new_n989), .A4(new_n488), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n988), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1035), .A2(G301), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1038), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n992), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1019), .A2(new_n986), .A3(new_n1020), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n1041), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1024), .A2(new_n1040), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1044), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1029), .A2(new_n1031), .A3(new_n801), .ZN(new_n1058));
  NAND3_X1  g633(.A1(G160), .A2(G40), .A3(new_n1038), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n986), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1058), .B(G168), .C1(new_n1061), .C2(G1966), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1057), .B1(new_n1062), .B2(G8), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1065));
  INV_X1    g640(.A(G1966), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(G168), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(new_n1062), .C1(new_n1068), .C2(new_n1057), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n538), .B2(new_n546), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1072), .A2(KEYINPUT111), .A3(KEYINPUT55), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT111), .B1(new_n1072), .B2(KEYINPUT55), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1072), .A2(KEYINPUT110), .A3(KEYINPUT55), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT110), .B1(new_n1072), .B2(KEYINPUT55), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1073), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1026), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n992), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1019), .A2(KEYINPUT50), .A3(new_n1020), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n763), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1039), .A2(new_n845), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1077), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(G40), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1086), .B(new_n477), .C1(new_n490), .C2(new_n495), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n601), .A2(G1976), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(G8), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT52), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n992), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n1071), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT49), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n543), .A2(G86), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n608), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G1981), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1094), .B(new_n1097), .C1(G305), .C2(G1981), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n604), .A2(new_n609), .A3(G1981), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1097), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT49), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(G288), .B2(new_n834), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1088), .A2(G8), .A3(new_n1089), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1091), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1029), .A2(new_n1031), .A3(new_n763), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1083), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(G8), .A3(new_n1077), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1071), .B1(new_n1107), .B2(new_n1083), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(KEYINPUT112), .A3(new_n1077), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1085), .B(new_n1106), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1033), .B1(new_n1032), .B2(new_n728), .ZN(new_n1115));
  AOI211_X1 g690(.A(KEYINPUT124), .B(G1961), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1043), .B(new_n1040), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G171), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1049), .A2(G171), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT54), .A3(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1056), .A2(new_n1070), .A3(new_n1114), .A4(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n591), .A2(KEYINPUT57), .A3(new_n596), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n591), .B2(new_n596), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n721), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1046), .A2(new_n1037), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1956), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n1087), .A2(new_n1037), .A3(new_n1038), .A4(new_n1128), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1124), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT119), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT61), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1127), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT120), .B1(new_n1142), .B2(KEYINPUT119), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1137), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1145), .A2(G1348), .B1(G2067), .B2(new_n1088), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT121), .B(new_n634), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1150));
  INV_X1    g725(.A(G1348), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1032), .A2(new_n1151), .B1(new_n1009), .B2(new_n1092), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n635), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n634), .A2(KEYINPUT121), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1148), .A2(new_n1150), .A3(new_n1156), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT115), .B(G1996), .Z(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1087), .A2(new_n1037), .A3(new_n1038), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT116), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT58), .B(G1341), .Z(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1162), .B(new_n1163), .C1(new_n1092), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1088), .A2(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1163), .B1(new_n1168), .B2(new_n1162), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n1171));
  XNOR2_X1  g746(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n576), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1162), .B1(new_n1092), .B2(new_n1165), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT116), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1175), .A2(new_n576), .A3(new_n1166), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1175), .A2(new_n576), .A3(new_n1166), .A4(new_n1172), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT118), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1173), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1144), .A2(new_n1157), .A3(new_n1159), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1146), .A2(new_n635), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1182), .A2(KEYINPUT114), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1141), .B1(new_n1182), .B2(KEYINPUT114), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1140), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1121), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1085), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1091), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1112), .A2(KEYINPUT112), .A3(new_n1077), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT112), .B1(new_n1112), .B2(new_n1077), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1188), .B(new_n1189), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1058), .B1(new_n1061), .B2(G1966), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1193), .A2(G8), .A3(G168), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1187), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1106), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1194), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1112), .A2(new_n1077), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1196), .A2(KEYINPUT63), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1057), .B1(new_n1193), .B2(G286), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1062), .A2(G8), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT62), .B1(new_n1203), .B2(new_n1063), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1064), .A2(new_n1069), .A3(new_n1206), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1204), .A2(new_n1114), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1111), .A2(new_n1189), .A3(new_n1113), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n601), .A2(new_n834), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT113), .Z(new_n1211));
  NOR2_X1   g786(.A1(new_n1211), .A2(new_n1102), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1093), .B1(new_n1212), .B2(new_n1099), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1200), .A2(new_n1208), .A3(new_n1209), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1017), .B1(new_n1186), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1010), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n993), .B1(new_n774), .B2(new_n1216), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1004), .A2(KEYINPUT46), .A3(new_n1006), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT46), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1220), .B(new_n1221), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n787), .A2(G2067), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n993), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1016), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1008), .A2(KEYINPUT126), .A3(new_n1012), .A4(new_n1015), .ZN(new_n1228));
  XNOR2_X1  g803(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n999), .B(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  AND3_X1   g806(.A1(new_n1222), .A2(new_n1225), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1215), .A2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g808(.A(new_n963), .ZN(new_n1235));
  OAI21_X1  g809(.A(new_n970), .B1(new_n962), .B2(new_n933), .ZN(new_n1236));
  OAI21_X1  g810(.A(KEYINPUT43), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g811(.A1(new_n959), .A2(new_n960), .ZN(new_n1238));
  NAND4_X1  g812(.A1(new_n1238), .A2(new_n972), .A3(new_n970), .A4(new_n969), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g814(.A1(G229), .A2(new_n463), .ZN(new_n1241));
  INV_X1    g815(.A(G227), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n677), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1243), .B1(new_n905), .B2(new_n910), .ZN(new_n1244));
  AND3_X1   g818(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .ZN(G308));
  NAND3_X1  g819(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .ZN(G225));
endmodule


