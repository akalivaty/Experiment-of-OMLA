

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n734), .ZN(n696) );
  AND2_X1 U553 ( .A1(n773), .A2(n518), .ZN(n774) );
  INV_X1 U554 ( .A(KEYINPUT102), .ZN(n705) );
  OR2_X1 U555 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U556 ( .A1(G543), .A2(n540), .ZN(n541) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n520) );
  NAND2_X1 U558 ( .A1(G286), .A2(G8), .ZN(n517) );
  OR2_X1 U559 ( .A1(n781), .A2(n772), .ZN(n518) );
  OR2_X1 U560 ( .A1(n754), .A2(KEYINPUT33), .ZN(n519) );
  XNOR2_X1 U561 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n697) );
  XNOR2_X1 U562 ( .A(n698), .B(n697), .ZN(n700) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n715) );
  XNOR2_X1 U564 ( .A(n716), .B(n715), .ZN(n720) );
  OR2_X1 U565 ( .A1(n744), .A2(n517), .ZN(n741) );
  XNOR2_X1 U566 ( .A(n742), .B(KEYINPUT32), .ZN(n749) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n758) );
  NOR2_X1 U568 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U569 ( .A1(G651), .A2(n637), .ZN(n645) );
  NOR2_X2 U570 ( .A1(n524), .A2(n523), .ZN(n875) );
  XNOR2_X1 U571 ( .A(KEYINPUT15), .B(n596), .ZN(n966) );
  NAND2_X1 U572 ( .A1(n879), .A2(G137), .ZN(n531) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XNOR2_X2 U574 ( .A(n521), .B(n520), .ZN(n879) );
  NAND2_X1 U575 ( .A1(n879), .A2(G138), .ZN(n530) );
  INV_X1 U576 ( .A(G2105), .ZN(n523) );
  NOR2_X4 U577 ( .A1(G2104), .A2(n523), .ZN(n874) );
  NAND2_X1 U578 ( .A1(G126), .A2(n874), .ZN(n522) );
  XNOR2_X1 U579 ( .A(KEYINPUT89), .B(n522), .ZN(n528) );
  INV_X1 U580 ( .A(G2104), .ZN(n524) );
  NAND2_X1 U581 ( .A1(G114), .A2(n875), .ZN(n526) );
  NOR2_X4 U582 ( .A1(G2105), .A2(n524), .ZN(n878) );
  NAND2_X1 U583 ( .A1(G102), .A2(n878), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  AND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(G164) );
  XNOR2_X1 U587 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U588 ( .A(n531), .B(KEYINPUT64), .ZN(n756) );
  NAND2_X1 U589 ( .A1(G101), .A2(n878), .ZN(n532) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(n532), .Z(n536) );
  NAND2_X1 U591 ( .A1(G125), .A2(n874), .ZN(n534) );
  NAND2_X1 U592 ( .A1(G113), .A2(n875), .ZN(n533) );
  AND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n684) );
  AND2_X1 U595 ( .A1(n756), .A2(n684), .ZN(G160) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U597 ( .A1(G85), .A2(n644), .ZN(n539) );
  XNOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n537), .B(KEYINPUT65), .ZN(n637) );
  INV_X1 U600 ( .A(G651), .ZN(n540) );
  NOR2_X1 U601 ( .A1(n637), .A2(n540), .ZN(n648) );
  NAND2_X1 U602 ( .A1(G72), .A2(n648), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n545) );
  NAND2_X1 U604 ( .A1(G47), .A2(n645), .ZN(n543) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n541), .Z(n643) );
  NAND2_X1 U606 ( .A1(G60), .A2(n643), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U608 ( .A1(n545), .A2(n544), .ZN(G290) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  NAND2_X1 U612 ( .A1(n643), .A2(G62), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n645), .A2(G50), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n644), .A2(G88), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT82), .ZN(n550) );
  NAND2_X1 U617 ( .A1(G75), .A2(n648), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT83), .B(n551), .Z(n552) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(G166) );
  NAND2_X1 U621 ( .A1(G64), .A2(n643), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT66), .B(n554), .Z(n561) );
  NAND2_X1 U623 ( .A1(G90), .A2(n644), .ZN(n556) );
  NAND2_X1 U624 ( .A1(G77), .A2(n648), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n557), .B(KEYINPUT9), .ZN(n559) );
  NAND2_X1 U627 ( .A1(G52), .A2(n645), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U629 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G51), .A2(n645), .ZN(n563) );
  NAND2_X1 U631 ( .A1(G63), .A2(n643), .ZN(n562) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U633 ( .A(KEYINPUT6), .B(n564), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G89), .A2(n644), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT4), .B(n565), .Z(n566) );
  XNOR2_X1 U636 ( .A(n566), .B(KEYINPUT75), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G76), .A2(n648), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U639 ( .A(n569), .B(KEYINPUT5), .Z(n570) );
  NOR2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U641 ( .A(KEYINPUT76), .B(n572), .Z(n573) );
  XNOR2_X1 U642 ( .A(KEYINPUT7), .B(n573), .ZN(G168) );
  XOR2_X1 U643 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U645 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U646 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n576) );
  INV_X1 U647 ( .A(G223), .ZN(n826) );
  NAND2_X1 U648 ( .A1(G567), .A2(n826), .ZN(n575) );
  XNOR2_X1 U649 ( .A(n576), .B(n575), .ZN(G234) );
  NAND2_X1 U650 ( .A1(n644), .A2(G81), .ZN(n577) );
  XNOR2_X1 U651 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G68), .A2(n648), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n580), .B(KEYINPUT13), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G43), .A2(n645), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n643), .A2(G56), .ZN(n583) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n583), .Z(n584) );
  NOR2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n586), .ZN(n984) );
  INV_X1 U661 ( .A(n984), .ZN(n613) );
  NAND2_X1 U662 ( .A1(G860), .A2(n613), .ZN(n587) );
  XNOR2_X1 U663 ( .A(n587), .B(KEYINPUT72), .ZN(G153) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G92), .A2(n644), .ZN(n588) );
  XNOR2_X1 U667 ( .A(n588), .B(KEYINPUT74), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G79), .A2(n648), .ZN(n590) );
  NAND2_X1 U669 ( .A1(G54), .A2(n645), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U671 ( .A1(G66), .A2(n643), .ZN(n591) );
  XNOR2_X1 U672 ( .A(KEYINPUT73), .B(n591), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U674 ( .A(n966), .ZN(n611) );
  INV_X1 U675 ( .A(G868), .ZN(n655) );
  NAND2_X1 U676 ( .A1(n611), .A2(n655), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G53), .A2(n645), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n599), .B(KEYINPUT68), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G91), .A2(n644), .ZN(n601) );
  NAND2_X1 U681 ( .A1(G78), .A2(n648), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G65), .A2(n643), .ZN(n602) );
  XNOR2_X1 U684 ( .A(KEYINPUT67), .B(n602), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(G299) );
  NAND2_X1 U687 ( .A1(G868), .A2(G286), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G299), .A2(n655), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(G297) );
  INV_X1 U690 ( .A(G860), .ZN(n628) );
  NAND2_X1 U691 ( .A1(n628), .A2(G559), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n609), .A2(n966), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U695 ( .A1(n655), .A2(n612), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n613), .A2(G868), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U698 ( .A(KEYINPUT77), .B(n616), .ZN(G282) );
  XNOR2_X1 U699 ( .A(G2100), .B(KEYINPUT79), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n874), .A2(G123), .ZN(n617) );
  XNOR2_X1 U701 ( .A(n617), .B(KEYINPUT18), .ZN(n619) );
  NAND2_X1 U702 ( .A1(G135), .A2(n879), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT78), .B(n620), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G111), .A2(n875), .ZN(n622) );
  NAND2_X1 U706 ( .A1(G99), .A2(n878), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n925) );
  XNOR2_X1 U709 ( .A(n925), .B(G2096), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U711 ( .A1(G559), .A2(n966), .ZN(n627) );
  XOR2_X1 U712 ( .A(n984), .B(n627), .Z(n663) );
  NAND2_X1 U713 ( .A1(n628), .A2(n663), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G93), .A2(n644), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G55), .A2(n645), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n648), .A2(G80), .ZN(n631) );
  XOR2_X1 U718 ( .A(KEYINPUT80), .B(n631), .Z(n632) );
  NOR2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n643), .A2(G67), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n636), .B(n657), .ZN(G145) );
  NAND2_X1 U723 ( .A1(G49), .A2(n645), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G87), .A2(n637), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U726 ( .A1(n643), .A2(n640), .ZN(n642) );
  NAND2_X1 U727 ( .A1(G651), .A2(G74), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U729 ( .A1(n643), .A2(G61), .ZN(n653) );
  NAND2_X1 U730 ( .A1(G86), .A2(n644), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G48), .A2(n645), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n648), .A2(G73), .ZN(n649) );
  XOR2_X1 U734 ( .A(KEYINPUT2), .B(n649), .Z(n650) );
  NOR2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U737 ( .A(KEYINPUT81), .B(n654), .Z(G305) );
  NAND2_X1 U738 ( .A1(n655), .A2(n657), .ZN(n656) );
  XNOR2_X1 U739 ( .A(n656), .B(KEYINPUT84), .ZN(n666) );
  XNOR2_X1 U740 ( .A(G290), .B(n657), .ZN(n661) );
  XNOR2_X1 U741 ( .A(G288), .B(KEYINPUT19), .ZN(n659) );
  INV_X1 U742 ( .A(G299), .ZN(n969) );
  XNOR2_X1 U743 ( .A(G166), .B(n969), .ZN(n658) );
  XNOR2_X1 U744 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(G305), .ZN(n899) );
  XNOR2_X1 U747 ( .A(n899), .B(n663), .ZN(n664) );
  NAND2_X1 U748 ( .A1(G868), .A2(n664), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U754 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U756 ( .A1(G120), .A2(G69), .ZN(n671) );
  NOR2_X1 U757 ( .A1(G237), .A2(n671), .ZN(n672) );
  XNOR2_X1 U758 ( .A(KEYINPUT86), .B(n672), .ZN(n673) );
  NAND2_X1 U759 ( .A1(n673), .A2(G108), .ZN(n831) );
  NAND2_X1 U760 ( .A1(G567), .A2(n831), .ZN(n674) );
  XNOR2_X1 U761 ( .A(n674), .B(KEYINPUT87), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G219), .A2(G220), .ZN(n675) );
  XOR2_X1 U763 ( .A(KEYINPUT85), .B(n675), .Z(n676) );
  XNOR2_X1 U764 ( .A(KEYINPUT22), .B(n676), .ZN(n677) );
  NAND2_X1 U765 ( .A1(n677), .A2(G96), .ZN(n678) );
  OR2_X1 U766 ( .A1(G218), .A2(n678), .ZN(n832) );
  AND2_X1 U767 ( .A1(G2106), .A2(n832), .ZN(n679) );
  NOR2_X1 U768 ( .A1(n680), .A2(n679), .ZN(G319) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n682) );
  INV_X1 U770 ( .A(G319), .ZN(n681) );
  NOR2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U772 ( .A(n683), .B(KEYINPUT88), .ZN(n829) );
  NAND2_X1 U773 ( .A1(G36), .A2(n829), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  AND2_X1 U775 ( .A1(n684), .A2(G40), .ZN(n755) );
  AND2_X1 U776 ( .A1(n755), .A2(n756), .ZN(n685) );
  NAND2_X2 U777 ( .A1(n685), .A2(n758), .ZN(n734) );
  NAND2_X1 U778 ( .A1(G8), .A2(n734), .ZN(n781) );
  XNOR2_X1 U779 ( .A(KEYINPUT100), .B(G1996), .ZN(n947) );
  NAND2_X1 U780 ( .A1(n696), .A2(n947), .ZN(n686) );
  XNOR2_X1 U781 ( .A(n686), .B(KEYINPUT26), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G1341), .A2(n734), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n690) );
  INV_X1 U784 ( .A(KEYINPUT101), .ZN(n689) );
  XNOR2_X1 U785 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U786 ( .A1(n691), .A2(n984), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n704), .A2(n966), .ZN(n695) );
  NOR2_X1 U788 ( .A1(G2067), .A2(n734), .ZN(n693) );
  NOR2_X1 U789 ( .A1(n696), .A2(G1348), .ZN(n692) );
  NOR2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n703) );
  NAND2_X1 U792 ( .A1(G2072), .A2(n696), .ZN(n698) );
  AND2_X1 U793 ( .A1(n734), .A2(G1956), .ZN(n699) );
  NOR2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n710) );
  NOR2_X1 U795 ( .A1(n710), .A2(n969), .ZN(n702) );
  XNOR2_X1 U796 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n702), .B(n701), .ZN(n709) );
  AND2_X1 U798 ( .A1(n703), .A2(n709), .ZN(n708) );
  NOR2_X1 U799 ( .A1(n704), .A2(n966), .ZN(n706) );
  XNOR2_X1 U800 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n714) );
  INV_X1 U802 ( .A(n709), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n969), .A2(n710), .ZN(n711) );
  OR2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U806 ( .A1(G1961), .A2(n734), .ZN(n718) );
  XOR2_X1 U807 ( .A(KEYINPUT25), .B(G2078), .Z(n948) );
  NAND2_X1 U808 ( .A1(n696), .A2(n948), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G301), .A2(n721), .ZN(n719) );
  NOR2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n731) );
  NAND2_X1 U812 ( .A1(G301), .A2(n721), .ZN(n722) );
  XNOR2_X1 U813 ( .A(n722), .B(KEYINPUT103), .ZN(n728) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n781), .ZN(n723) );
  XOR2_X1 U815 ( .A(KEYINPUT97), .B(n723), .Z(n745) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n734), .ZN(n743) );
  NOR2_X1 U817 ( .A1(n745), .A2(n743), .ZN(n724) );
  NAND2_X1 U818 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U819 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U820 ( .A1(G168), .A2(n726), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(KEYINPUT31), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U824 ( .A(n732), .B(KEYINPUT104), .ZN(n744) );
  INV_X1 U825 ( .A(G8), .ZN(n739) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n781), .ZN(n733) );
  XNOR2_X1 U827 ( .A(KEYINPUT105), .B(n733), .ZN(n737) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U829 ( .A1(G166), .A2(n735), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n738) );
  OR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(G8), .A2(n743), .ZN(n747) );
  NOR2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U837 ( .A(n750), .B(KEYINPUT106), .ZN(n779) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n771) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n771), .A2(n751), .ZN(n982) );
  NAND2_X1 U841 ( .A1(n779), .A2(n982), .ZN(n752) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n967) );
  NAND2_X1 U843 ( .A1(n752), .A2(n967), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n781), .A2(n753), .ZN(n754) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n976) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n820) );
  NAND2_X1 U848 ( .A1(n875), .A2(G116), .ZN(n759) );
  XNOR2_X1 U849 ( .A(n759), .B(KEYINPUT90), .ZN(n761) );
  NAND2_X1 U850 ( .A1(G128), .A2(n874), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT35), .ZN(n767) );
  NAND2_X1 U853 ( .A1(G104), .A2(n878), .ZN(n764) );
  NAND2_X1 U854 ( .A1(G140), .A2(n879), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U856 ( .A(KEYINPUT34), .B(n765), .Z(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U858 ( .A(n768), .B(KEYINPUT36), .Z(n888) );
  XNOR2_X1 U859 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  OR2_X1 U860 ( .A1(n888), .A2(n818), .ZN(n769) );
  XNOR2_X1 U861 ( .A(KEYINPUT91), .B(n769), .ZN(n940) );
  NAND2_X1 U862 ( .A1(n820), .A2(n940), .ZN(n770) );
  XNOR2_X1 U863 ( .A(n770), .B(KEYINPUT92), .ZN(n817) );
  AND2_X1 U864 ( .A1(n976), .A2(n817), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n771), .A2(KEYINPUT33), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n519), .A2(n774), .ZN(n788) );
  INV_X1 U867 ( .A(n817), .ZN(n786) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U869 ( .A(n775), .B(KEYINPUT96), .Z(n776) );
  XNOR2_X1 U870 ( .A(KEYINPUT24), .B(n776), .ZN(n777) );
  OR2_X1 U871 ( .A1(n781), .A2(n777), .ZN(n784) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G8), .A2(n778), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n809) );
  NAND2_X1 U878 ( .A1(G129), .A2(n874), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G117), .A2(n875), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n878), .A2(G105), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U884 ( .A(KEYINPUT95), .B(n794), .Z(n796) );
  NAND2_X1 U885 ( .A1(n879), .A2(G141), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n892) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n892), .ZN(n806) );
  NAND2_X1 U888 ( .A1(n874), .A2(G119), .ZN(n797) );
  XOR2_X1 U889 ( .A(KEYINPUT93), .B(n797), .Z(n799) );
  NAND2_X1 U890 ( .A1(n875), .A2(G107), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT94), .B(n800), .Z(n804) );
  NAND2_X1 U893 ( .A1(n878), .A2(G95), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G131), .A2(n879), .ZN(n801) );
  AND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n860) );
  NAND2_X1 U897 ( .A1(G1991), .A2(n860), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n813) );
  INV_X1 U899 ( .A(n813), .ZN(n931) );
  XOR2_X1 U900 ( .A(G1986), .B(G290), .Z(n968) );
  NAND2_X1 U901 ( .A1(n931), .A2(n968), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n807), .A2(n820), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n824) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n892), .ZN(n933) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n860), .ZN(n929) );
  NOR2_X1 U907 ( .A1(n810), .A2(n929), .ZN(n811) );
  XOR2_X1 U908 ( .A(KEYINPUT107), .B(n811), .Z(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n933), .A2(n814), .ZN(n815) );
  XNOR2_X1 U911 ( .A(KEYINPUT39), .B(n815), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n888), .A2(n818), .ZN(n926) );
  NAND2_X1 U914 ( .A1(n819), .A2(n926), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT108), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U918 ( .A(KEYINPUT40), .B(n825), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U921 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n828) );
  XOR2_X1 U923 ( .A(KEYINPUT109), .B(n828), .Z(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G188) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(G325) );
  XOR2_X1 U926 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  XOR2_X1 U932 ( .A(KEYINPUT43), .B(G2678), .Z(n834) );
  XNOR2_X1 U933 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2072), .Z(n836) );
  XNOR2_X1 U936 ( .A(G2090), .B(G2067), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U938 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2100), .B(G2096), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U941 ( .A(G2078), .B(G2084), .Z(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1986), .B(G1976), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1956), .B(G1971), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n845), .B(G2474), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U949 ( .A(KEYINPUT41), .B(G1981), .Z(n849) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G124), .A2(n874), .ZN(n852) );
  XOR2_X1 U954 ( .A(KEYINPUT44), .B(n852), .Z(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(KEYINPUT113), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G112), .A2(n875), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G100), .A2(n878), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G136), .A2(n879), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U961 ( .A1(n859), .A2(n858), .ZN(G162) );
  XNOR2_X1 U962 ( .A(n925), .B(n860), .ZN(n895) );
  NAND2_X1 U963 ( .A1(G103), .A2(n878), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G139), .A2(n879), .ZN(n861) );
  NAND2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n875), .A2(G115), .ZN(n863) );
  XOR2_X1 U967 ( .A(KEYINPUT115), .B(n863), .Z(n865) );
  NAND2_X1 U968 ( .A1(n874), .A2(G127), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n918) );
  XOR2_X1 U972 ( .A(KEYINPUT116), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U975 ( .A(n871), .B(KEYINPUT114), .Z(n873) );
  XNOR2_X1 U976 ( .A(G164), .B(KEYINPUT46), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n873), .B(n872), .ZN(n886) );
  NAND2_X1 U978 ( .A1(G130), .A2(n874), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G118), .A2(n875), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G106), .A2(n878), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G142), .A2(n879), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(n882), .B(KEYINPUT45), .Z(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n887) );
  XOR2_X1 U987 ( .A(n887), .B(G162), .Z(n890) );
  XOR2_X1 U988 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n918), .B(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U994 ( .A(G286), .B(KEYINPUT119), .ZN(n898) );
  XNOR2_X1 U995 ( .A(G171), .B(n966), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n901) );
  XOR2_X1 U997 ( .A(n984), .B(n899), .Z(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2430), .Z(n904) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2443), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n910) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n906) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2427), .Z(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n911) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n911), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1018 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n923) );
  XOR2_X1 U1019 ( .A(G2072), .B(n918), .Z(n920) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(n921), .B(KEYINPUT50), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(n923), .B(n922), .ZN(n938) );
  XOR2_X1 U1024 ( .A(G2084), .B(G160), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT51), .B(n934), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n962) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n962), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n957) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(n947), .B(G32), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1056 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n965), .ZN(n1021) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1060 ( .A(G1348), .B(n966), .ZN(n975) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(G1956), .B(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT122), .B(n978), .Z(n979) );
  XNOR2_X1 U1070 ( .A(KEYINPUT57), .B(n979), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(G171), .B(G1961), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G1341), .B(n984), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1019) );
  INV_X1 U1078 ( .A(G16), .ZN(n1017) );
  XOR2_X1 U1079 ( .A(G1986), .B(G24), .Z(n993) );
  XNOR2_X1 U1080 ( .A(G1971), .B(KEYINPUT127), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(G22), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(KEYINPUT58), .B(n996), .Z(n1014) );
  XOR2_X1 U1086 ( .A(G1961), .B(G5), .Z(n1009) );
  XOR2_X1 U1087 ( .A(KEYINPUT124), .B(G4), .Z(n998) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n998), .B(n997), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT123), .B(G1956), .Z(n999) );
  XNOR2_X1 U1091 ( .A(G20), .B(n999), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G6), .B(G1981), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(KEYINPUT125), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT60), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1012), .Z(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

