//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  XNOR2_X1  g000(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT18), .A2(G131), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT70), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G237), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT85), .A2(G143), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n194), .A2(G214), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G214), .ZN(new_n198));
  AOI211_X1 g012(.A(new_n198), .B(G953), .C1(new_n191), .C2(new_n193), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT85), .B(G143), .Z(new_n200));
  OAI211_X1 g014(.A(new_n189), .B(new_n197), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT87), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(G214), .A3(new_n195), .ZN(new_n204));
  INV_X1    g018(.A(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n206), .A2(KEYINPUT87), .A3(new_n189), .A4(new_n197), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G125), .B(G140), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n212));
  INV_X1    g026(.A(new_n189), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT86), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n212), .A2(KEYINPUT86), .A3(new_n213), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n208), .B(new_n211), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n197), .ZN(new_n217));
  AOI21_X1  g031(.A(G953), .B1(new_n191), .B2(new_n193), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n200), .B1(G214), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n222), .A3(new_n197), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G125), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(KEYINPUT16), .A3(G140), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n209), .A2(KEYINPUT16), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G125), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT74), .B1(new_n230), .B2(KEYINPUT16), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n210), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(G146), .A3(new_n231), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n212), .A2(KEYINPUT17), .A3(G131), .ZN(new_n237));
  AOI21_X1  g051(.A(G146), .B1(new_n228), .B2(new_n231), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n227), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n225), .A2(G140), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n240), .A3(KEYINPUT16), .ZN(new_n241));
  AND4_X1   g055(.A1(G146), .A2(new_n239), .A3(new_n231), .A4(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT89), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n224), .A2(new_n236), .A3(new_n237), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G113), .B(G122), .ZN(new_n245));
  INV_X1    g059(.A(G104), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT88), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n216), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n216), .A2(new_n244), .A3(new_n251), .A4(new_n248), .ZN(new_n252));
  INV_X1    g066(.A(new_n247), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n220), .A2(new_n223), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n209), .B(KEYINPUT19), .Z(new_n255));
  OAI211_X1 g069(.A(new_n254), .B(new_n234), .C1(G146), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n216), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n250), .A2(new_n252), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G475), .ZN(new_n259));
  INV_X1    g073(.A(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n188), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n250), .A2(new_n252), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n253), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n259), .A3(new_n260), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n262), .B1(new_n266), .B2(KEYINPUT20), .ZN(new_n267));
  INV_X1    g081(.A(G952), .ZN(new_n268));
  AOI211_X1 g082(.A(G953), .B(new_n268), .C1(G234), .C2(G237), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n260), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT21), .B(G898), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n216), .A2(new_n244), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT91), .B1(new_n274), .B2(new_n253), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT91), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n277), .B(new_n247), .C1(new_n216), .C2(new_n244), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n263), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT92), .A3(new_n260), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G475), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n275), .A2(new_n278), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n283), .B2(new_n263), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT92), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n267), .B(new_n273), .C1(new_n282), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT97), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G116), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n291), .A3(G122), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n288), .A2(G122), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(KEYINPUT14), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT14), .ZN(new_n296));
  OAI21_X1  g110(.A(G107), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G107), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n299), .A3(new_n293), .ZN(new_n300));
  INV_X1    g114(.A(G143), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G128), .ZN(new_n302));
  INV_X1    g116(.A(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G143), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G134), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n300), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT93), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n292), .A2(new_n299), .A3(new_n293), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n299), .B1(new_n292), .B2(new_n293), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n294), .A2(G107), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT93), .A3(new_n300), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT13), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT94), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n302), .B2(new_n319), .ZN(new_n321));
  AOI211_X1 g135(.A(KEYINPUT94), .B(KEYINPUT13), .C1(new_n301), .C2(G128), .ZN(new_n322));
  OAI221_X1 g136(.A(new_n304), .B1(new_n319), .B2(new_n302), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n307), .B1(new_n323), .B2(G134), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n318), .A2(KEYINPUT95), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT95), .B1(new_n318), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n311), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT9), .B(G234), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(G217), .A3(new_n195), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n311), .B(new_n332), .C1(new_n325), .C2(new_n326), .ZN(new_n333));
  AOI21_X1  g147(.A(G902), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT96), .ZN(new_n335));
  INV_X1    g149(.A(G478), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT15), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n334), .B2(new_n335), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n287), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n335), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n337), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(KEYINPUT97), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n286), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G210), .B1(G237), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n210), .A2(G143), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n301), .A2(G146), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT0), .A2(G128), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G143), .B(G146), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G128), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G125), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n351), .A2(new_n352), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n303), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT1), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n351), .A2(new_n352), .A3(new_n361), .A4(G128), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n301), .A2(KEYINPUT1), .A3(G146), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n360), .A2(new_n362), .A3(new_n225), .A4(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n350), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G224), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G953), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT80), .B1(new_n357), .B2(G125), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n358), .A2(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT7), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n369), .A2(KEYINPUT7), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G119), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  OAI21_X1  g191(.A(G113), .B1(new_n377), .B2(KEYINPUT5), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n289), .A2(new_n291), .A3(G119), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT67), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n288), .B2(G119), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT66), .B(G116), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT67), .A3(G119), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n378), .B1(new_n386), .B2(KEYINPUT5), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT2), .B(G113), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n383), .B2(new_n385), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n299), .B2(G104), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n299), .A2(G104), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n246), .A2(KEYINPUT77), .A3(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G101), .ZN(new_n395));
  INV_X1    g209(.A(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n246), .A2(G107), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n299), .A2(KEYINPUT3), .A3(G104), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT3), .B1(new_n299), .B2(G104), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n387), .A2(new_n389), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n389), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT5), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n381), .B1(new_n384), .B2(G119), .ZN(new_n405));
  AND4_X1   g219(.A1(KEYINPUT67), .A2(new_n289), .A3(new_n291), .A4(G119), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT68), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n383), .A2(new_n385), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n404), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n403), .B1(new_n410), .B2(new_n378), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n402), .B1(new_n411), .B2(new_n401), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G122), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT8), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n375), .B(KEYINPUT82), .C1(new_n412), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n388), .A3(new_n409), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT69), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n389), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G101), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n424), .A3(G101), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n407), .A2(new_n418), .A3(new_n409), .A4(new_n388), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n395), .A2(new_n400), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n403), .B(new_n429), .C1(new_n410), .C2(new_n378), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n413), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n416), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n383), .A2(new_n385), .A3(new_n408), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n408), .B1(new_n383), .B2(new_n385), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT5), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n378), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n429), .B1(new_n437), .B2(new_n403), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n414), .B1(new_n438), .B2(new_n402), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT82), .B1(new_n439), .B2(new_n375), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n260), .B1(new_n432), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n428), .A2(new_n430), .ZN(new_n442));
  INV_X1    g256(.A(new_n413), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n365), .A2(new_n368), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(new_n367), .Z(new_n447));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n349), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n375), .B1(new_n412), .B2(new_n415), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n431), .A3(new_n416), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n260), .A4(new_n348), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(KEYINPUT83), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(new_n349), .C1(new_n441), .C2(new_n450), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G472), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT64), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n357), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n306), .B2(G137), .ZN(new_n469));
  INV_X1    g283(.A(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT11), .A3(G134), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n306), .A2(G137), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G131), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(new_n471), .A3(new_n222), .A4(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n354), .B(KEYINPUT64), .C1(new_n355), .C2(new_n356), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n360), .A2(new_n363), .A3(new_n362), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT65), .B1(new_n306), .B2(G137), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n306), .A2(KEYINPUT65), .A3(G137), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n475), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n420), .A2(new_n485), .A3(new_n427), .ZN(new_n486));
  INV_X1    g300(.A(new_n357), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n484), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n420), .B2(new_n427), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n465), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n218), .A2(G210), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT27), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G101), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n420), .A2(new_n427), .ZN(new_n496));
  INV_X1    g310(.A(new_n489), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n491), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n485), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n488), .A2(new_n484), .A3(KEYINPUT30), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n504), .A2(new_n420), .A3(new_n427), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n498), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n501), .B(new_n502), .C1(new_n495), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n490), .A2(KEYINPUT28), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n420), .A2(new_n489), .A3(new_n427), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n498), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n510), .B1(new_n512), .B2(KEYINPUT28), .ZN(new_n513));
  INV_X1    g327(.A(new_n495), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n502), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n464), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n495), .A3(new_n498), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT31), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n506), .A2(new_n521), .A3(new_n498), .A4(new_n495), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n495), .B1(new_n491), .B2(new_n500), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT32), .ZN(new_n526));
  INV_X1    g340(.A(new_n465), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n420), .A2(new_n485), .A3(new_n427), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n498), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n514), .B1(new_n529), .B2(new_n510), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n520), .A3(new_n522), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n518), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n517), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n303), .A2(G119), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n376), .A2(G128), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT24), .B(G110), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n376), .A2(G128), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT73), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n536), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n539), .B1(new_n547), .B2(G110), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n242), .B2(new_n238), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n537), .A2(new_n538), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n547), .B2(G110), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n209), .A2(new_n210), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n234), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n553), .A3(KEYINPUT75), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  INV_X1    g369(.A(G221), .ZN(new_n556));
  INV_X1    g370(.A(G234), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n556), .A2(new_n557), .A3(G953), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n555), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT75), .B1(new_n549), .B2(new_n553), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g376(.A(KEYINPUT75), .B(new_n559), .C1(new_n549), .C2(new_n553), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n260), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT25), .B(new_n260), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G217), .B1(new_n557), .B2(G902), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(KEYINPUT72), .Z(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n260), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT76), .Z(new_n572));
  OR2_X1    g386(.A1(new_n562), .A2(new_n563), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n568), .A2(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n534), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n556), .B1(new_n329), .B2(new_n260), .ZN(new_n577));
  XNOR2_X1  g391(.A(G110), .B(G140), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n195), .A2(G227), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT78), .ZN(new_n582));
  AOI21_X1  g396(.A(G128), .B1(new_n351), .B2(new_n352), .ZN(new_n583));
  INV_X1    g397(.A(new_n363), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n363), .B(KEYINPUT78), .C1(new_n355), .C2(G128), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n362), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n429), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n476), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n423), .A2(new_n487), .A3(new_n425), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n429), .A2(KEYINPUT10), .A3(new_n479), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n401), .A2(new_n360), .A3(new_n363), .A4(new_n362), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT12), .B1(new_n596), .B2(new_n476), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT12), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n598), .B(new_n591), .C1(new_n588), .C2(new_n595), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(KEYINPUT79), .B(new_n594), .C1(new_n597), .C2(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n581), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n594), .A2(new_n581), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n362), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n363), .B1(new_n355), .B2(G128), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n582), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n401), .B1(new_n610), .B2(new_n586), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n592), .B(new_n593), .C1(new_n611), .C2(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n476), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(G469), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G469), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n597), .A2(new_n599), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n606), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n581), .B1(new_n613), .B2(new_n594), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n616), .B(new_n260), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(G469), .A2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n577), .B1(new_n615), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n347), .A2(new_n463), .A3(new_n576), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  AOI21_X1  g440(.A(new_n464), .B1(new_n531), .B2(new_n260), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n627), .A2(KEYINPUT98), .ZN(new_n628));
  INV_X1    g442(.A(new_n518), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n520), .A2(new_n522), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n530), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n628), .A2(new_n632), .A3(new_n624), .A4(new_n574), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n459), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n635), .B(new_n272), .C1(new_n451), .C2(new_n457), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n331), .A2(new_n333), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n318), .A2(new_n324), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT95), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n318), .A2(KEYINPUT95), .A3(new_n324), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n310), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n642), .B2(KEYINPUT99), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n637), .A2(new_n643), .ZN(new_n645));
  OAI21_X1  g459(.A(G478), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n334), .A2(new_n336), .ZN(new_n647));
  NAND2_X1  g461(.A1(G478), .A2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n259), .B1(new_n284), .B2(KEYINPUT92), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n280), .A2(new_n260), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT92), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n649), .B1(new_n654), .B2(new_n267), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n634), .A2(new_n636), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  NAND4_X1  g472(.A1(new_n265), .A2(new_n259), .A3(new_n260), .A4(new_n187), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n262), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n346), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n634), .A2(new_n661), .A3(new_n636), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n568), .A2(new_n570), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n549), .A2(new_n553), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n572), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n628), .A2(new_n632), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n347), .A2(new_n463), .A3(new_n672), .A4(new_n624), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AND3_X1   g489(.A1(new_n531), .A2(new_n532), .A3(new_n518), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n532), .B1(new_n531), .B2(new_n518), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n509), .A2(new_n516), .ZN(new_n678));
  OAI22_X1  g492(.A1(new_n676), .A2(new_n677), .B1(new_n678), .B2(new_n464), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n635), .B1(new_n451), .B2(new_n457), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n679), .A2(new_n680), .A3(new_n624), .A4(new_n671), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n270), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n269), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n346), .A2(new_n654), .A3(new_n660), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n526), .A2(new_n533), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n498), .A2(new_n511), .ZN(new_n691));
  AOI21_X1  g505(.A(G902), .B1(new_n691), .B2(new_n514), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n507), .A2(new_n495), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n464), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n689), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(KEYINPUT101), .B(new_n694), .C1(new_n526), .C2(new_n533), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n635), .A3(new_n671), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n267), .B1(new_n282), .B2(new_n285), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n458), .A2(new_n461), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n699), .A2(new_n346), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n685), .B(KEYINPUT39), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n624), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT40), .Z(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  INV_X1    g525(.A(new_n649), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n700), .A2(new_n712), .A3(new_n685), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n679), .A2(new_n680), .A3(new_n624), .A4(new_n671), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n210), .ZN(G48));
  OR2_X1    g530(.A1(new_n597), .A2(new_n599), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n613), .A2(new_n594), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n717), .A2(new_n607), .B1(new_n718), .B2(new_n580), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  INV_X1    g534(.A(new_n577), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n620), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n534), .A2(new_n575), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n636), .A3(new_n655), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND3_X1  g540(.A1(new_n661), .A2(new_n723), .A3(new_n636), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  INV_X1    g542(.A(new_n286), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n635), .B(new_n722), .C1(new_n451), .C2(new_n457), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n669), .B1(new_n568), .B2(new_n570), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n534), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n341), .A2(new_n345), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n730), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND2_X1  g549(.A1(new_n531), .A2(new_n260), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G472), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n500), .B1(new_n691), .B2(new_n499), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n514), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n630), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n518), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n574), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n720), .A2(new_n721), .A3(new_n620), .A4(new_n273), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n346), .A3(new_n700), .A4(new_n680), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  AOI21_X1  g560(.A(new_n629), .B1(new_n630), .B2(new_n739), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n731), .A2(new_n627), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n655), .A2(new_n730), .A3(new_n685), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  AND3_X1   g564(.A1(new_n700), .A2(new_n712), .A3(new_n685), .ZN(new_n751));
  INV_X1    g565(.A(new_n614), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n604), .A2(new_n616), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n721), .B1(new_n753), .B2(new_n622), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n635), .B(new_n754), .C1(new_n458), .C2(new_n461), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(KEYINPUT42), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n751), .A2(new_n755), .A3(new_n576), .A4(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n635), .B1(new_n458), .B2(new_n461), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n576), .A3(new_n624), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n713), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n346), .A2(new_n654), .A3(new_n660), .A4(new_n685), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT104), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n755), .A2(new_n686), .A3(new_n768), .A4(new_n576), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  INV_X1    g585(.A(new_n760), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n712), .A2(new_n267), .A3(new_n654), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT43), .Z(new_n774));
  AOI21_X1  g588(.A(new_n731), .B1(new_n628), .B2(new_n632), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n605), .A2(KEYINPUT45), .A3(new_n614), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n604), .B2(new_n752), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(G469), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n782), .B2(new_n621), .ZN(new_n783));
  INV_X1    g597(.A(new_n620), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n621), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n577), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n707), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n778), .B(new_n789), .C1(new_n777), .C2(new_n776), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  NAND2_X1  g605(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n787), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n751), .A2(new_n575), .A3(new_n534), .A4(new_n760), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NAND3_X1  g612(.A1(new_n574), .A2(new_n459), .A3(new_n721), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT106), .ZN(new_n800));
  INV_X1    g614(.A(new_n720), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n784), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT49), .Z(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n703), .ZN(new_n805));
  INV_X1    g619(.A(new_n773), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n698), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT107), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n634), .A2(new_n463), .A3(new_n273), .A4(new_n655), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n625), .A3(new_n673), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n727), .A2(new_n734), .A3(new_n724), .A4(new_n745), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n339), .B2(new_n340), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n343), .A2(KEYINPUT109), .A3(new_n344), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n286), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT110), .B1(new_n817), .B2(new_n463), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n462), .A2(new_n286), .A3(new_n819), .A4(new_n816), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n634), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n650), .A2(new_n653), .B1(new_n262), .B2(new_n659), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n685), .A3(new_n816), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n760), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT111), .B1(new_n772), .B2(new_n824), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n534), .A2(new_n754), .A3(new_n731), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n751), .A2(new_n755), .A3(new_n748), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n764), .A2(new_n770), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n835));
  INV_X1    g649(.A(new_n685), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n754), .A2(new_n671), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n696), .B2(new_n697), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n700), .A2(new_n346), .A3(new_n680), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n615), .A2(new_n623), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n721), .A3(new_n731), .A4(new_n685), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n695), .B1(new_n676), .B2(new_n677), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n690), .A2(new_n689), .A3(new_n695), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n700), .A2(new_n346), .A3(new_n680), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT112), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n829), .A2(new_n680), .A3(new_n655), .A4(new_n685), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n687), .A2(new_n850), .A3(new_n749), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n834), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n700), .A2(new_n748), .A3(new_n712), .A4(new_n685), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n680), .A2(new_n721), .A3(new_n802), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n853), .A2(new_n854), .B1(new_n714), .B2(new_n766), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n715), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n848), .A4(new_n840), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n852), .A2(new_n857), .B1(KEYINPUT52), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n833), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n810), .A2(new_n821), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n852), .A2(new_n857), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n811), .B(KEYINPUT108), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n764), .A2(new_n770), .A3(new_n830), .A4(new_n831), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n859), .B1(new_n864), .B2(KEYINPUT53), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n867), .A3(KEYINPUT53), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n724), .A2(new_n745), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT108), .A3(new_n727), .A4(new_n734), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT108), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n811), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n872), .A3(new_n810), .A4(new_n821), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n832), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n858), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT113), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n861), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n876), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n868), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n866), .B1(new_n880), .B2(KEYINPUT54), .ZN(new_n881));
  INV_X1    g695(.A(new_n742), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n774), .A2(new_n269), .A3(new_n882), .ZN(new_n883));
  OR4_X1    g697(.A1(new_n459), .A2(new_n883), .A3(new_n703), .A4(new_n722), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n884), .A2(KEYINPUT50), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(KEYINPUT50), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n772), .A2(new_n684), .A3(new_n722), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n774), .A2(new_n748), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n574), .A3(new_n698), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n889), .A2(new_n700), .A3(new_n712), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n885), .A2(new_n886), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n802), .A2(new_n577), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n772), .B(new_n883), .C1(new_n795), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT114), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n894), .A2(KEYINPUT51), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(KEYINPUT51), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n268), .A2(G953), .ZN(new_n897));
  INV_X1    g711(.A(new_n655), .ZN(new_n898));
  OAI221_X1 g712(.A(new_n897), .B1(new_n889), .B2(new_n898), .C1(new_n883), .C2(new_n854), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n774), .A2(new_n576), .A3(new_n887), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n901), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n902));
  XOR2_X1   g716(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n903));
  AOI211_X1 g717(.A(new_n899), .B(new_n902), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n881), .A2(new_n895), .A3(new_n896), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n808), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n195), .A2(G952), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT53), .B1(new_n874), .B2(new_n861), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n833), .A2(new_n858), .ZN(new_n910));
  OAI211_X1 g724(.A(G210), .B(G902), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n445), .A2(new_n449), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n447), .Z(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(KEYINPUT56), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n908), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n865), .A2(KEYINPUT117), .A3(G210), .A4(G902), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n915), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n922), .B2(new_n915), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(KEYINPUT119), .B(new_n917), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G51));
  XNOR2_X1  g744(.A(new_n865), .B(KEYINPUT54), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n621), .B(KEYINPUT57), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n719), .B1(new_n933), .B2(KEYINPUT120), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(KEYINPUT120), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n865), .A2(G902), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(new_n782), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n908), .B1(new_n935), .B2(new_n937), .ZN(G54));
  INV_X1    g752(.A(new_n908), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT58), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n936), .A2(new_n940), .A3(new_n259), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n265), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n265), .B2(new_n941), .ZN(G60));
  XOR2_X1   g757(.A(new_n648), .B(KEYINPUT59), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n863), .A2(new_n862), .A3(new_n860), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n838), .A2(new_n835), .A3(new_n839), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT112), .B1(new_n846), .B2(new_n847), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT52), .B1(new_n949), .B2(new_n856), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n849), .A2(new_n834), .A3(new_n851), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n876), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n953), .A2(new_n867), .B1(new_n864), .B2(KEYINPUT53), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n878), .A2(KEYINPUT113), .A3(new_n876), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT54), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n944), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n644), .A2(new_n645), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT121), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n961));
  INV_X1    g775(.A(new_n959), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n961), .B(new_n962), .C1(new_n881), .C2(new_n944), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n944), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n908), .B1(new_n931), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n960), .A2(new_n963), .A3(KEYINPUT122), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  AND2_X1   g786(.A1(new_n865), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n939), .B1(new_n973), .B2(new_n573), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n668), .B2(new_n973), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g790(.A(G953), .B1(new_n271), .B2(new_n366), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT123), .ZN(new_n978));
  INV_X1    g792(.A(new_n873), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT124), .Z(new_n981));
  OAI21_X1  g795(.A(new_n912), .B1(G898), .B2(new_n195), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G69));
  NAND2_X1  g797(.A1(new_n504), .A2(new_n505), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(new_n255), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n790), .A2(new_n770), .A3(new_n797), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n789), .A2(new_n576), .A3(new_n847), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n764), .A3(new_n856), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n195), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n682), .A2(G953), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n989), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n710), .A2(new_n856), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n898), .B1(new_n700), .B2(new_n816), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n998), .A2(new_n576), .A3(new_n707), .A4(new_n755), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n790), .A2(new_n797), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n996), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n985), .A2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n994), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(G72));
  NOR3_X1   g820(.A1(new_n986), .A2(new_n873), .A3(new_n988), .ZN(new_n1007));
  XOR2_X1   g821(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1008));
  NOR2_X1   g822(.A1(new_n464), .A2(new_n260), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OR3_X1    g824(.A1(new_n1007), .A2(KEYINPUT127), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n507), .A2(new_n495), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT127), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1010), .B1(new_n1002), .B2(new_n979), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1014), .B(new_n939), .C1(new_n693), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n693), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1017), .A2(new_n1012), .A3(new_n1010), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1016), .B1(new_n880), .B2(new_n1018), .ZN(G57));
endmodule


