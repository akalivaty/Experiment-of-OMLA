//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT21), .B(G898), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G214), .B1(G237), .B2(G902), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT9), .B(G234), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT9), .B(G234), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT75), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n198), .A2(G217), .A3(new_n188), .A4(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT89), .B1(new_n202), .B2(G143), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G122), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G122), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n215), .A3(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n203), .A2(new_n206), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n209), .B1(new_n221), .B2(KEYINPUT13), .ZN(new_n222));
  AOI211_X1 g036(.A(KEYINPUT90), .B(KEYINPUT13), .C1(new_n203), .C2(new_n206), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT13), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n207), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n222), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n220), .B1(new_n227), .B2(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n213), .A2(KEYINPUT14), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n217), .A2(new_n229), .A3(G107), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n213), .B(new_n215), .C1(KEYINPUT14), .C2(new_n218), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(G134), .B1(new_n221), .B2(new_n209), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n211), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n201), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n234), .ZN(new_n236));
  INV_X1    g050(.A(new_n201), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT90), .B1(new_n221), .B2(KEYINPUT13), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n207), .A2(new_n224), .A3(new_n225), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n208), .B1(new_n240), .B2(new_n222), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n236), .B(new_n237), .C1(new_n241), .C2(new_n220), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G902), .ZN(new_n244));
  INV_X1    g058(.A(G478), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n245), .A2(KEYINPUT15), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(G902), .B1(new_n235), .B2(new_n242), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(new_n246), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G140), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G125), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G140), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT72), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n188), .A3(G214), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n205), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT18), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n268), .A2(KEYINPUT86), .A3(new_n272), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT86), .B1(new_n268), .B2(new_n272), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n262), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(KEYINPUT66), .A2(G131), .ZN(new_n278));
  NOR2_X1   g092(.A1(KEYINPUT66), .A2(G131), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n268), .A2(KEYINPUT17), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(KEYINPUT87), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n268), .A2(new_n281), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT17), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n265), .A2(new_n280), .A3(new_n267), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n253), .A2(KEYINPUT16), .A3(G140), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT16), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n255), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n259), .ZN(new_n292));
  OAI211_X1 g106(.A(G146), .B(new_n289), .C1(new_n255), .C2(new_n290), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n283), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G113), .B(G122), .ZN(new_n296));
  INV_X1    g110(.A(G104), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n298), .B(new_n277), .C1(new_n283), .C2(new_n294), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n244), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G475), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT19), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n257), .A2(new_n258), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n255), .A2(KEYINPUT19), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n259), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n284), .A2(new_n286), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n293), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n277), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n299), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n301), .ZN(new_n313));
  NOR2_X1   g127(.A1(G475), .A2(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT20), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n313), .A2(KEYINPUT88), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n314), .ZN(new_n320));
  AOI211_X1 g134(.A(KEYINPUT20), .B(new_n320), .C1(new_n312), .C2(new_n301), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(KEYINPUT88), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n250), .B(new_n304), .C1(new_n319), .C2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G210), .B1(G237), .B2(G902), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT85), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n297), .A2(G107), .ZN(new_n328));
  AND2_X1   g142(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n329));
  NOR2_X1   g143(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G101), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n328), .B(KEYINPUT77), .C1(new_n330), .C2(new_n329), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n218), .B2(G104), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n218), .A2(G104), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n333), .A2(new_n334), .A3(new_n335), .A4(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n218), .A2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n328), .B2(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n340), .B2(new_n343), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n214), .A2(KEYINPUT5), .A3(G119), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT83), .ZN(new_n347));
  INV_X1    g161(.A(G113), .ZN(new_n348));
  XNOR2_X1  g162(.A(G116), .B(G119), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(KEYINPUT5), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT2), .B(G113), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n349), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n344), .A2(new_n345), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n331), .A2(new_n332), .B1(new_n338), .B2(new_n337), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n334), .B1(new_n358), .B2(new_n335), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n361));
  OR2_X1    g175(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n338), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n339), .B1(new_n364), .B2(KEYINPUT77), .ZN(new_n365));
  INV_X1    g179(.A(new_n335), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n361), .B(G101), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n349), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n352), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n354), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n327), .B1(new_n356), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n340), .A2(new_n343), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n351), .A2(new_n354), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n365), .B2(new_n366), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n370), .A3(new_n367), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n381), .A3(new_n326), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(new_n327), .C1(new_n356), .C2(new_n372), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT65), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n205), .B2(G146), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n259), .A2(KEYINPUT65), .A3(G143), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n205), .A2(G146), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT0), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n202), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n259), .A2(G143), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n394), .A2(new_n389), .B1(KEYINPUT0), .B2(G128), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n391), .A3(new_n202), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G125), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n388), .A2(new_n389), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n387), .A4(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n387), .A2(new_n388), .A3(new_n405), .A4(new_n389), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT67), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n394), .A2(new_n389), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n202), .B1(new_n394), .B2(KEYINPUT1), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n402), .B1(new_n414), .B2(G125), .ZN(new_n415));
  INV_X1    g229(.A(G224), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n383), .A2(new_n385), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n355), .A2(new_n374), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n378), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n326), .B(KEYINPUT8), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n417), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT7), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n415), .B(new_n426), .C1(KEYINPUT84), .C2(new_n417), .ZN(new_n427));
  INV_X1    g241(.A(new_n426), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n390), .A2(new_n392), .B1(new_n395), .B2(new_n399), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n253), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n412), .B1(new_n406), .B2(new_n408), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(new_n253), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n417), .A2(KEYINPUT84), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n382), .A2(new_n427), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n244), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n325), .B1(new_n419), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n382), .A2(new_n427), .A3(new_n434), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  INV_X1    g253(.A(new_n325), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n383), .A2(new_n385), .A3(new_n418), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n195), .B(new_n323), .C1(new_n437), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n198), .A2(new_n200), .ZN(new_n444));
  OAI21_X1  g258(.A(G221), .B1(new_n444), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n367), .A2(new_n429), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT78), .B1(new_n360), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n401), .B1(new_n359), .B2(new_n361), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n380), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n344), .A2(new_n345), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT10), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n431), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n407), .B(new_n404), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n390), .A2(new_n411), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n340), .B(new_n343), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n454), .A2(new_n456), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT11), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n208), .B2(G137), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n208), .A2(G137), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT11), .A3(G134), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G131), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n280), .A2(new_n463), .A3(new_n462), .A4(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n453), .A2(new_n460), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  INV_X1    g286(.A(G227), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G953), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n472), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT80), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n453), .A2(new_n460), .A3(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n459), .A2(new_n455), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n375), .A2(new_n456), .A3(new_n376), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n450), .A2(new_n380), .A3(new_n451), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n451), .B1(new_n450), .B2(new_n380), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n470), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n478), .A2(new_n480), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n459), .B1(new_n454), .B2(new_n414), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n490), .A2(KEYINPUT12), .A3(new_n469), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n490), .B2(new_n469), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n471), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(new_n475), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n447), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n484), .A2(new_n485), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n483), .A2(new_n482), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n487), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n469), .A3(new_n481), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n471), .A2(new_n479), .A3(new_n476), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n479), .B1(new_n471), .B2(new_n476), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n475), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n446), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n476), .B1(new_n499), .B2(new_n471), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n471), .B(new_n476), .C1(new_n491), .C2(new_n492), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n446), .B(new_n244), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(G469), .A2(G902), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n443), .B(new_n445), .C1(new_n505), .C2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n503), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT82), .B1(new_n502), .B2(new_n503), .ZN(new_n517));
  OAI21_X1  g331(.A(G469), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(KEYINPUT91), .A3(new_n445), .A4(new_n443), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n292), .A2(new_n293), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n202), .A2(G119), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT71), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT24), .B(G110), .Z(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n535));
  INV_X1    g349(.A(new_n528), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n527), .B(new_n535), .C1(new_n536), .C2(KEYINPUT23), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G110), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n525), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(G110), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(new_n531), .B2(new_n532), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n293), .B(new_n260), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n539), .A2(KEYINPUT73), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT73), .B1(new_n539), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n524), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n542), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n523), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n244), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n545), .A2(KEYINPUT25), .A3(new_n244), .A4(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G217), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(G234), .B2(new_n244), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n545), .A2(new_n548), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT74), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n429), .A2(new_n469), .ZN(new_n563));
  INV_X1    g377(.A(new_n370), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n464), .A2(G134), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n463), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G131), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n468), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n409), .B2(new_n413), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT68), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n370), .B1(new_n429), .B2(new_n469), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT68), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n573), .C1(new_n431), .C2(new_n569), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n266), .A2(G210), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n571), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT69), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT30), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n568), .B(new_n468), .C1(new_n457), .C2(new_n412), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(new_n563), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n563), .B(new_n582), .C1(new_n431), .C2(new_n569), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n370), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT69), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n571), .A2(new_n574), .A3(new_n588), .A4(new_n578), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n580), .A2(new_n581), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n565), .A2(new_n570), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT28), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n563), .B1(new_n431), .B2(new_n569), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n370), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n571), .A2(new_n574), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n592), .B1(new_n595), .B2(KEYINPUT28), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n590), .B1(new_n578), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n587), .A2(new_n589), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n581), .B1(new_n598), .B2(new_n580), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n562), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n580), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n587), .A2(new_n589), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT31), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n596), .ZN(new_n604));
  INV_X1    g418(.A(new_n578), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT70), .A4(new_n590), .ZN(new_n607));
  NOR2_X1   g421(.A1(G472), .A2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT32), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n600), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n593), .A2(KEYINPUT30), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n564), .B1(new_n613), .B2(new_n585), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n571), .A2(new_n574), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT29), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n578), .B2(new_n596), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n596), .A2(KEYINPUT29), .A3(new_n578), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n244), .ZN(new_n621));
  OAI21_X1  g435(.A(G472), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n600), .A2(new_n608), .A3(new_n607), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n610), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n561), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n514), .A2(new_n520), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  NAND3_X1  g442(.A1(new_n600), .A2(new_n244), .A3(new_n607), .ZN(new_n629));
  INV_X1    g443(.A(G472), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(KEYINPUT92), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n561), .ZN(new_n636));
  INV_X1    g450(.A(new_n445), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n515), .B2(new_n518), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n437), .A2(KEYINPUT93), .A3(new_n442), .ZN(new_n640));
  INV_X1    g454(.A(new_n194), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT93), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n640), .A2(new_n644), .A3(new_n193), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n201), .B(KEYINPUT94), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n228), .B2(new_n234), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n227), .A2(G134), .ZN(new_n652));
  INV_X1    g466(.A(new_n220), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n234), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n651), .B1(new_n654), .B2(new_n237), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n647), .B(KEYINPUT95), .C1(new_n228), .C2(new_n234), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n650), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n243), .A2(new_n651), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n245), .A2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n657), .A2(KEYINPUT96), .A3(new_n658), .A4(new_n659), .ZN(new_n663));
  INV_X1    g477(.A(new_n248), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT97), .B(G478), .Z(new_n665));
  AOI22_X1  g479(.A1(new_n662), .A2(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(KEYINPUT88), .B2(new_n321), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT88), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n315), .B2(KEYINPUT20), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n668), .A2(new_n670), .B1(G475), .B2(new_n303), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n646), .B1(new_n666), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n662), .A2(new_n663), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n664), .A2(new_n665), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n304), .B1(new_n319), .B2(new_n322), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(KEYINPUT98), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n645), .B1(new_n672), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n639), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n297), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  OAI21_X1  g496(.A(new_n304), .B1(new_n321), .B2(new_n667), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(new_n250), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n645), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n639), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NOR2_X1   g502(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n546), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n557), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT100), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n556), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n632), .A2(new_n633), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n514), .A2(new_n520), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  AOI21_X1  g512(.A(new_n693), .B1(new_n623), .B2(new_n625), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n640), .A2(new_n644), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n189), .B(KEYINPUT101), .Z(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(G900), .B2(new_n192), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n700), .A2(new_n684), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n638), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  INV_X1    g520(.A(new_n442), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n642), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT38), .Z(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n601), .A2(new_n602), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n605), .B2(new_n595), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n712), .B2(G902), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n625), .A2(new_n612), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n250), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n676), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n693), .A2(new_n194), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n710), .A2(new_n715), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n702), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n638), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n675), .A2(new_n676), .A3(new_n702), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n700), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n666), .A2(new_n671), .A3(new_n703), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n640), .A4(new_n644), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n638), .A3(new_n699), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  NAND3_X1  g548(.A1(new_n625), .A2(new_n612), .A3(new_n622), .ZN(new_n735));
  INV_X1    g549(.A(new_n509), .ZN(new_n736));
  INV_X1    g550(.A(new_n471), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n488), .B2(new_n481), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n507), .B1(new_n738), .B2(new_n476), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n446), .B1(new_n739), .B2(new_n244), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n736), .A2(new_n740), .A3(new_n637), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n678), .A2(new_n735), .A3(new_n741), .A4(new_n636), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT104), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n742), .B(new_n744), .ZN(G15));
  NAND4_X1  g559(.A1(new_n741), .A2(new_n735), .A3(new_n685), .A4(new_n636), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  OAI21_X1  g561(.A(new_n244), .B1(new_n506), .B2(new_n508), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n445), .A2(new_n749), .A3(new_n509), .A4(new_n193), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n700), .A2(new_n323), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n699), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  INV_X1    g567(.A(new_n597), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n609), .B1(new_n754), .B2(new_n603), .ZN(new_n755));
  AOI211_X1 g569(.A(new_n755), .B(new_n561), .C1(new_n629), .C2(G472), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n700), .A2(new_n717), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NOR2_X1   g573(.A1(new_n700), .A2(new_n728), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n736), .A2(new_n740), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n445), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n755), .B1(new_n629), .B2(G472), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n694), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT105), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n755), .B(new_n693), .C1(G472), .C2(new_n629), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n741), .A3(new_n767), .A4(new_n760), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NOR2_X1   g584(.A1(new_n637), .A2(new_n641), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n708), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n502), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT106), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n446), .B(new_n494), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n773), .B(new_n730), .C1(new_n777), .C2(new_n511), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n624), .A2(new_n610), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n612), .A2(new_n622), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n636), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT107), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT42), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n478), .A2(new_n480), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT106), .B1(new_n784), .B2(new_n499), .ZN(new_n785));
  INV_X1    g599(.A(new_n776), .ZN(new_n786));
  OAI211_X1 g600(.A(G469), .B(new_n503), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n772), .B1(new_n515), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n626), .A2(new_n788), .A3(new_n789), .A4(new_n730), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n782), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n778), .A2(new_n783), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n781), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n626), .A2(KEYINPUT108), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  NOR2_X1   g612(.A1(new_n684), .A2(new_n703), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n626), .A2(new_n788), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G134), .ZN(G36));
  NAND2_X1  g615(.A1(new_n675), .A2(new_n671), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(KEYINPUT109), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n634), .A2(new_n694), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT110), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n708), .A2(new_n194), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n807), .B2(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT45), .B(new_n503), .C1(new_n785), .C2(new_n786), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n495), .A2(new_n504), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n814), .B(G469), .C1(new_n815), .C2(KEYINPUT45), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT46), .B1(new_n816), .B2(new_n510), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n736), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(KEYINPUT46), .A3(new_n510), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n637), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n721), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n464), .ZN(G39));
  XNOR2_X1  g637(.A(new_n820), .B(KEYINPUT47), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n735), .A2(new_n811), .A3(new_n636), .A4(new_n728), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NAND2_X1  g641(.A1(new_n636), .A2(new_n771), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n709), .A2(new_n802), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n761), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n715), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  INV_X1    g648(.A(new_n701), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n806), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT114), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n741), .A3(new_n756), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n710), .A2(new_n641), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n811), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n741), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n764), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT118), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n842), .A2(new_n834), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n839), .A2(new_n840), .B1(KEYINPUT116), .B2(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n845), .A2(new_n561), .A3(new_n189), .A4(new_n714), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n671), .A3(new_n666), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n843), .A2(new_n848), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n838), .A2(new_n756), .A3(new_n844), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n830), .A2(new_n445), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n824), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n839), .A2(new_n700), .ZN(new_n858));
  INV_X1    g672(.A(G952), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n677), .A2(new_n672), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n859), .B(G953), .C1(new_n851), .C2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n858), .A2(KEYINPUT119), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n794), .A2(new_n795), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n846), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT48), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT119), .B1(new_n858), .B2(new_n861), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n855), .B(KEYINPUT115), .Z(new_n868));
  OAI21_X1  g682(.A(new_n854), .B1(new_n824), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n857), .B(new_n867), .C1(new_n870), .C2(KEYINPUT51), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n323), .B1(new_n675), .B2(new_n671), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n708), .A3(new_n195), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n635), .A2(new_n638), .A3(new_n636), .A4(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n627), .A2(new_n696), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n752), .A2(new_n742), .A3(new_n758), .A4(new_n746), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n811), .A2(new_n716), .A3(new_n683), .A4(new_n703), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n699), .A2(new_n638), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n788), .A2(new_n766), .A3(new_n730), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n800), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n881), .A3(new_n797), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT111), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT111), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n875), .A2(new_n881), .A3(new_n797), .A4(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n638), .B(new_n699), .C1(new_n732), .C2(new_n704), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n515), .A2(new_n787), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n694), .A2(new_n637), .A3(new_n703), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n714), .A3(new_n889), .A4(new_n757), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n769), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n769), .A2(new_n887), .A3(KEYINPUT112), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(KEYINPUT52), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT53), .B1(new_n886), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n883), .A2(new_n885), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n891), .A2(KEYINPUT52), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n895), .B2(new_n896), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n900), .A2(KEYINPUT54), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n886), .B2(new_n899), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT52), .B1(new_n893), .B2(new_n894), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n909), .A2(new_n882), .A3(new_n902), .A4(new_n904), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT113), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n906), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n906), .B2(new_n912), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n871), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n859), .A2(new_n188), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT120), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n833), .B1(new_n916), .B2(new_n918), .ZN(G75));
  AND3_X1   g733(.A1(new_n893), .A2(KEYINPUT52), .A3(new_n894), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n909), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n921), .B2(new_n901), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n910), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n244), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n325), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n383), .A2(new_n385), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n418), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  NOR2_X1   g742(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n925), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n188), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n928), .B1(new_n925), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(G51));
  XNOR2_X1  g751(.A(new_n923), .B(new_n908), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n510), .B(KEYINPUT57), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n739), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n923), .A2(new_n244), .A3(new_n816), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n932), .B1(new_n941), .B2(new_n942), .ZN(G54));
  NAND3_X1  g757(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n944));
  INV_X1    g758(.A(new_n313), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n947), .A3(new_n932), .ZN(G60));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT59), .Z(new_n951));
  AOI21_X1  g765(.A(new_n904), .B1(new_n921), .B2(new_n901), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n908), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n922), .A2(KEYINPUT54), .A3(new_n910), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT113), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n906), .A2(new_n912), .A3(new_n913), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n657), .A2(new_n658), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n949), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n951), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n914), .B2(new_n915), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(KEYINPUT122), .A3(new_n959), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n959), .A2(new_n951), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n932), .B1(new_n938), .B2(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  XOR2_X1   g783(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n923), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n560), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n923), .A2(new_n971), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n690), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n933), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G66));
  OAI21_X1  g792(.A(G953), .B1(new_n190), .B2(new_n416), .ZN(new_n979));
  INV_X1    g793(.A(new_n876), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n875), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n979), .B1(new_n982), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n926), .B1(G898), .B2(new_n188), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  NOR2_X1   g799(.A1(new_n584), .A2(new_n586), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n306), .A2(new_n307), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n989));
  NOR4_X1   g803(.A1(new_n722), .A2(new_n781), .A3(new_n811), .A4(new_n872), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n822), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n769), .A2(new_n887), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n725), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(new_n826), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n988), .B(new_n989), .C1(new_n996), .C2(new_n188), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n473), .A2(G900), .A3(G953), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n992), .B1(new_n813), .B2(new_n821), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT126), .Z(new_n1000));
  OR4_X1    g814(.A1(new_n700), .A2(new_n821), .A3(new_n717), .A4(new_n863), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n797), .A2(new_n1001), .A3(new_n800), .A4(new_n826), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n998), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n997), .B1(new_n1004), .B2(new_n988), .ZN(G72));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  INV_X1    g821(.A(new_n616), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n711), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n952), .A2(new_n953), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1007), .B1(new_n996), .B2(new_n981), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1011), .B(new_n578), .C1(new_n615), .C2(new_n614), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n933), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1000), .A2(new_n982), .A3(new_n1002), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n1007), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1014), .A2(KEYINPUT127), .A3(new_n1007), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n614), .A2(new_n615), .A3(new_n578), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n1010), .B(new_n1013), .C1(new_n1019), .C2(new_n1020), .ZN(G57));
endmodule


