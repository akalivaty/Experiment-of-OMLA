//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  AND2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(KEYINPUT3), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT68), .B(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(new_n464), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n463), .B(G2104), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G2105), .B1(G101), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n474), .A2(new_n482), .ZN(G160));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n467), .B2(new_n472), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  INV_X1    g061(.A(G100), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n487), .A2(new_n484), .A3(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n487), .B2(new_n484), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G112), .B2(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G136), .B2(new_n473), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR4_X1   g068(.A1(new_n478), .A2(KEYINPUT4), .A3(new_n493), .A4(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI211_X1 g070(.A(new_n493), .B(G2105), .C1(new_n467), .C2(new_n472), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n484), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT72), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT71), .B(G114), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n508), .A2(new_n509), .A3(new_n484), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n499), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n505), .B1(new_n508), .B2(new_n484), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n502), .A2(G114), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n514));
  OAI211_X1 g089(.A(KEYINPUT72), .B(G2105), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n512), .A2(KEYINPUT73), .A3(new_n515), .A4(G2104), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n511), .A2(new_n516), .B1(G126), .B2(new_n485), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n498), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n525), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  INV_X1    g108(.A(new_n529), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n534), .A2(G51), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n522), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n526), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G168));
  INV_X1    g119(.A(new_n527), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G52), .Z(new_n546));
  AOI22_X1  g121(.A1(G90), .A2(new_n545), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT75), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n524), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n540), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n524), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(new_n556), .B2(new_n555), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT77), .B(G43), .ZN(new_n559));
  AOI22_X1  g134(.A1(G81), .A2(new_n545), .B1(new_n534), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(new_n534), .A2(G53), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n545), .A2(G91), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(G78), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G78), .ZN(new_n574));
  INV_X1    g149(.A(G543), .ZN(new_n575));
  NOR3_X1   g150(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT78), .ZN(new_n576));
  AOI211_X1 g151(.A(new_n573), .B(new_n576), .C1(G65), .C2(new_n522), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n571), .B1(new_n577), .B2(new_n524), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G299));
  INV_X1    g155(.A(G168), .ZN(G286));
  OAI21_X1  g156(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n529), .B2(new_n583), .C1(new_n584), .C2(new_n527), .ZN(G288));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n520), .B2(new_n521), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n522), .A2(new_n526), .A3(G86), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n524), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n527), .A2(new_n595), .B1(new_n529), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(new_n545), .A2(G92), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT10), .Z(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n540), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n534), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G321));
  NOR2_X1   g185(.A1(G168), .A2(new_n607), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(G299), .B2(new_n607), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT79), .Z(G297));
  XNOR2_X1  g188(.A(new_n612), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g189(.A(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n561), .A2(new_n607), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n606), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n473), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n485), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n484), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n484), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n627), .A2(new_n628), .A3(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(G401));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n650), .A2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n651), .B1(new_n657), .B2(KEYINPUT17), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n652), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n659), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n655), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n670), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n673), .B(new_n676), .C1(new_n667), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n685));
  OR2_X1    g260(.A1(G288), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(G288), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(G23), .B(new_n688), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  NAND4_X1  g276(.A1(new_n692), .A2(new_n693), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT89), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n702), .A2(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(KEYINPUT89), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(KEYINPUT34), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G24), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n598), .B(KEYINPUT86), .Z(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n473), .A2(G131), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n485), .A2(G119), .ZN(new_n716));
  OR2_X1    g291(.A1(G95), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G107), .C2(new_n484), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n713), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT85), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n721), .B(new_n723), .Z(new_n724));
  NOR2_X1   g299(.A1(new_n712), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n705), .A2(new_n708), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT36), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n705), .A2(new_n728), .A3(new_n708), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT97), .ZN(new_n731));
  NOR2_X1   g306(.A1(G171), .A2(new_n694), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G5), .B2(new_n694), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT93), .Z(new_n736));
  NOR2_X1   g311(.A1(new_n626), .A2(new_n713), .ZN(new_n737));
  INV_X1    g312(.A(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n740));
  OR2_X1    g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  NAND2_X1  g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G168), .A2(new_n694), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n694), .B2(G21), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n737), .B(new_n747), .C1(new_n746), .C2(new_n745), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n736), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT94), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n713), .A2(G32), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n485), .A2(G129), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT26), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(G105), .B2(new_n481), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n473), .A2(G141), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n751), .B1(new_n761), .B2(new_n713), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT27), .Z(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G1996), .ZN(new_n764));
  NOR2_X1   g339(.A1(G29), .A2(G35), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G162), .B2(G29), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2090), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  OR3_X1    g346(.A1(new_n764), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n562), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G16), .B2(G19), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n713), .B1(new_n776), .B2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G160), .B2(G29), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n774), .A2(new_n775), .B1(G2084), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n694), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT23), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n579), .B2(new_n694), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n780), .B(new_n786), .C1(G2084), .C2(new_n779), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n733), .A2(new_n734), .ZN(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT90), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n606), .B2(new_n694), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1348), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n788), .B(new_n792), .C1(new_n775), .C2(new_n774), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n787), .B(new_n793), .C1(G1996), .C2(new_n763), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n713), .A2(G26), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n473), .A2(G140), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n485), .A2(G128), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n484), .A2(G116), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NOR2_X1   g378(.A1(G27), .A2(G29), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G164), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G2078), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n794), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G29), .A2(G33), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n473), .A2(G139), .ZN(new_n810));
  INV_X1    g385(.A(G127), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n478), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G115), .B2(G2104), .ZN(new_n813));
  NAND2_X1  g388(.A1(G103), .A2(G2104), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(G2105), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(KEYINPUT25), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n814), .A2(new_n817), .A3(G2105), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n810), .B1(new_n484), .B2(new_n813), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT91), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT92), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n809), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2072), .ZN(new_n823));
  NOR4_X1   g398(.A1(new_n750), .A2(new_n772), .A3(new_n808), .A4(new_n823), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n730), .A2(new_n731), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n731), .B1(new_n730), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n730), .A2(new_n824), .ZN(G150));
  XNOR2_X1  g403(.A(KEYINPUT98), .B(G93), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n527), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n524), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n830), .B(new_n832), .C1(G55), .C2(new_n534), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n561), .B1(new_n833), .B2(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n615), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n834), .B1(new_n842), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n836), .B1(new_n845), .B2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n518), .B(new_n801), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n761), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n820), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n821), .B2(new_n849), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n719), .B(KEYINPUT103), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n630), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n484), .A2(KEYINPUT102), .A3(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT102), .B1(new_n484), .B2(G118), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  AND4_X1   g431(.A1(G2104), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n473), .A2(G142), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT101), .Z(new_n859));
  AOI211_X1 g434(.A(new_n857), .B(new_n859), .C1(G130), .C2(new_n485), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n853), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n851), .A2(new_n861), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n626), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n862), .A2(new_n865), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n869), .B(new_n870), .C1(new_n868), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g448(.A(new_n839), .B(new_n619), .Z(new_n874));
  NOR2_X1   g449(.A1(new_n615), .A2(G299), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n606), .A2(new_n579), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n875), .A2(new_n880), .A3(new_n876), .ZN(new_n881));
  INV_X1    g456(.A(new_n875), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n876), .B1(new_n882), .B2(KEYINPUT105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(KEYINPUT105), .B2(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n884), .B2(new_n880), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n885), .B2(new_n874), .ZN(new_n886));
  XNOR2_X1  g461(.A(G303), .B(G305), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n688), .B(new_n598), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(KEYINPUT106), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(KEYINPUT106), .B2(new_n889), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n889), .A2(KEYINPUT106), .A3(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT42), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n886), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G868), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G868), .B2(new_n833), .ZN(G295));
  XOR2_X1   g472(.A(G295), .B(KEYINPUT107), .Z(G331));
  XNOR2_X1  g473(.A(G301), .B(G286), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n839), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n878), .B2(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(new_n893), .ZN(new_n903));
  AOI21_X1  g478(.A(G37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n893), .B(KEYINPUT108), .Z(new_n905));
  AND2_X1   g480(.A1(new_n900), .A2(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n884), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n905), .B(new_n907), .C1(new_n878), .C2(new_n906), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n905), .B(new_n901), .C1(new_n878), .C2(new_n900), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n912), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT44), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n904), .A2(new_n911), .A3(new_n909), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n904), .A2(new_n908), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n917), .B(new_n918), .C1(new_n909), .C2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n914), .B1(new_n920), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n485), .A2(G126), .ZN(new_n923));
  OAI21_X1  g498(.A(G2105), .B1(new_n513), .B2(new_n514), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n464), .B1(new_n924), .B2(new_n505), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT73), .B1(new_n925), .B2(new_n515), .ZN(new_n926));
  AND4_X1   g501(.A1(KEYINPUT73), .A2(new_n512), .A3(G2104), .A4(new_n515), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n932), .B2(G2104), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n466), .A2(KEYINPUT69), .A3(new_n464), .ZN(new_n934));
  OAI211_X1 g509(.A(G138), .B(new_n484), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n494), .B1(new_n935), .B2(KEYINPUT4), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n922), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n474), .A2(G40), .A3(new_n482), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(G1996), .A3(new_n760), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n801), .B(G2067), .Z(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(G1996), .B2(new_n760), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n942), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n719), .B(new_n723), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(G290), .A2(G1986), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n942), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n951), .B2(G1996), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT125), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n945), .B(new_n761), .C1(new_n959), .C2(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n942), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n961), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  NAND2_X1  g542(.A1(new_n720), .A2(new_n723), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n949), .A2(new_n968), .B1(G2067), .B2(new_n801), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n958), .B(new_n967), .C1(new_n942), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT124), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n498), .B2(new_n517), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n940), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(KEYINPUT50), .B(G1384), .C1(new_n498), .C2(new_n517), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n785), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n977));
  NAND2_X1  g552(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n579), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n570), .C2(new_n578), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n518), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT56), .B(G2072), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n939), .A2(new_n940), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n976), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n982), .B1(new_n976), .B2(new_n985), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT61), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n985), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n941), .B1(new_n937), .B2(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n518), .A2(new_n973), .A3(new_n922), .ZN(new_n992));
  AOI21_X1  g567(.A(G1956), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n981), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n976), .A2(new_n982), .A3(new_n985), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT61), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n940), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n939), .A2(new_n983), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n518), .A2(new_n922), .A3(new_n940), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT58), .B(G1341), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n562), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(KEYINPUT117), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(KEYINPUT118), .A3(new_n562), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1010), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT118), .B1(new_n1005), .B2(new_n562), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n1007), .B(new_n561), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n997), .A2(new_n998), .A3(new_n1012), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n988), .B1(new_n986), .B2(new_n987), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n994), .A2(KEYINPUT61), .A3(new_n995), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT119), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1348), .B1(new_n991), .B2(new_n992), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1002), .A2(G2067), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1024), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n974), .A2(new_n975), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n1027), .C1(new_n1028), .C2(G1348), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n606), .B1(new_n1030), .B2(KEYINPUT60), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1032), .B(new_n615), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1031), .A2(new_n1033), .B1(KEYINPUT60), .B2(new_n1030), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1017), .A2(new_n1022), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n994), .B1(new_n1030), .B2(new_n606), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n995), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT120), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G168), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n1044), .B2(KEYINPUT121), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n939), .A2(new_n940), .A3(new_n983), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n940), .A3(new_n992), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1047), .A2(G1966), .B1(G2084), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(new_n1046), .C1(new_n1050), .C2(G286), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1044), .ZN(new_n1052));
  INV_X1    g627(.A(G2084), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n939), .A2(new_n940), .A3(new_n983), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1028), .A2(new_n1053), .B1(new_n1054), .B2(new_n746), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1052), .B(new_n1045), .C1(new_n1055), .C2(new_n1043), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(new_n1044), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n939), .A2(new_n806), .A3(new_n983), .A4(new_n940), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1049), .A2(new_n734), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1064));
  OAI21_X1  g639(.A(G171), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1047), .A2(new_n1066), .A3(KEYINPUT53), .A4(new_n806), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1060), .A2(new_n1059), .B1(new_n1049), .B2(new_n734), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1059), .A2(KEYINPUT122), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(G301), .A4(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1070), .A3(KEYINPUT54), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1048), .A2(new_n769), .A3(new_n992), .A4(new_n940), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT111), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n991), .A2(new_n1074), .A3(new_n769), .A4(new_n992), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1054), .A2(new_n697), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G303), .A2(G8), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT55), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(G8), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n686), .A2(G1976), .A3(new_n687), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1002), .A2(G8), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1090));
  INV_X1    g665(.A(G1981), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n589), .B2(KEYINPUT113), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n589), .A2(new_n1093), .A3(new_n590), .A4(new_n591), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1002), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1043), .B1(new_n972), .B2(new_n940), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n1086), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1085), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1002), .A2(G8), .A3(new_n1086), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n1089), .A4(new_n1098), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1084), .A2(new_n1079), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1058), .A2(new_n1071), .A3(new_n1082), .A4(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1068), .B(G301), .C1(new_n1060), .C2(new_n1059), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT54), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1028), .A2(new_n769), .B1(new_n1054), .B2(new_n697), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1079), .B1(new_n1114), .B2(new_n1043), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1082), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1044), .B1(new_n1050), .B2(G8), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1118), .A2(new_n1045), .B1(new_n1050), .B2(new_n1044), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(new_n1051), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .A4(new_n1071), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1113), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1039), .A2(new_n1041), .A3(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1117), .A2(new_n1110), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI211_X1 g706(.A(G1976), .B(G288), .C1(new_n1101), .C2(new_n1097), .ZN(new_n1132));
  NOR2_X1   g707(.A1(G305), .A2(G1981), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1101), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1105), .A2(new_n1089), .A3(new_n1098), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1082), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1050), .A2(G8), .A3(G168), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1117), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1138), .A2(new_n1137), .A3(new_n1135), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1077), .A2(G8), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1079), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1082), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1136), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1127), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n954), .ZN(new_n1147));
  NAND2_X1  g722(.A1(G290), .A2(G1986), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n951), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n953), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n971), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1150), .ZN(new_n1152));
  AOI211_X1 g727(.A(KEYINPUT124), .B(new_n1152), .C1(new_n1127), .C2(new_n1145), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n970), .B1(new_n1151), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g729(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1156));
  AND2_X1   g730(.A1(new_n913), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n1157), .A2(new_n872), .ZN(G225));
  INV_X1    g732(.A(G225), .ZN(G308));
endmodule


