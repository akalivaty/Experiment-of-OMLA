

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594;

  XNOR2_X1 U329 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U330 ( .A(n418), .B(KEYINPUT123), .ZN(n419) );
  XNOR2_X1 U331 ( .A(n420), .B(n419), .ZN(n442) );
  NOR2_X1 U332 ( .A1(n472), .A2(n578), .ZN(n443) );
  XNOR2_X1 U333 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U334 ( .A(n461), .B(KEYINPUT58), .ZN(n462) );
  XNOR2_X1 U335 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT74), .B(G85GAT), .Z(n298) );
  XNOR2_X1 U337 ( .A(G99GAT), .B(G106GAT), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n380) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n324) );
  XOR2_X1 U340 ( .A(n380), .B(n324), .Z(n300) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U342 ( .A(n300), .B(n299), .Z(n317) );
  XOR2_X1 U343 ( .A(KEYINPUT79), .B(KEYINPUT9), .Z(n302) );
  XNOR2_X1 U344 ( .A(KEYINPUT11), .B(KEYINPUT80), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n304) );
  INV_X1 U346 ( .A(KEYINPUT78), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n308) );
  INV_X1 U348 ( .A(n308), .ZN(n306) );
  XOR2_X1 U349 ( .A(G43GAT), .B(G134GAT), .Z(n456) );
  XNOR2_X1 U350 ( .A(n456), .B(KEYINPUT10), .ZN(n307) );
  INV_X1 U351 ( .A(n307), .ZN(n305) );
  NAND2_X1 U352 ( .A1(n306), .A2(n305), .ZN(n310) );
  NAND2_X1 U353 ( .A1(n308), .A2(n307), .ZN(n309) );
  NAND2_X1 U354 ( .A1(n310), .A2(n309), .ZN(n315) );
  XNOR2_X1 U355 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n311), .B(KEYINPUT7), .ZN(n365) );
  XNOR2_X1 U357 ( .A(n365), .B(KEYINPUT64), .ZN(n313) );
  INV_X1 U358 ( .A(KEYINPUT65), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U360 ( .A(KEYINPUT81), .B(G92GAT), .Z(n319) );
  XNOR2_X1 U361 ( .A(G190GAT), .B(G218GAT), .ZN(n318) );
  XNOR2_X1 U362 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U363 ( .A(G36GAT), .B(n320), .Z(n349) );
  XNOR2_X1 U364 ( .A(n321), .B(n349), .ZN(n565) );
  XNOR2_X1 U365 ( .A(KEYINPUT82), .B(n565), .ZN(n548) );
  XOR2_X1 U366 ( .A(G106GAT), .B(G218GAT), .Z(n323) );
  XOR2_X1 U367 ( .A(G22GAT), .B(G155GAT), .Z(n404) );
  XOR2_X1 U368 ( .A(KEYINPUT73), .B(G148GAT), .Z(n377) );
  XNOR2_X1 U369 ( .A(n404), .B(n377), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U371 ( .A(n325), .B(n324), .Z(n330) );
  XOR2_X1 U372 ( .A(KEYINPUT24), .B(G204GAT), .Z(n327) );
  NAND2_X1 U373 ( .A1(G228GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U375 ( .A(KEYINPUT93), .B(n328), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U377 ( .A(G211GAT), .B(KEYINPUT22), .Z(n332) );
  XNOR2_X1 U378 ( .A(G78GAT), .B(KEYINPUT23), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U380 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U381 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n336) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n335) );
  XNOR2_X1 U383 ( .A(n336), .B(n335), .ZN(n434) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n337), .B(KEYINPUT91), .ZN(n350) );
  XNOR2_X1 U386 ( .A(n434), .B(n350), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n472) );
  XNOR2_X1 U388 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n340), .B(KEYINPUT18), .ZN(n341) );
  XOR2_X1 U390 ( .A(n341), .B(KEYINPUT17), .Z(n343) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G176GAT), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n450) );
  XOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT75), .Z(n378) );
  XOR2_X1 U394 ( .A(KEYINPUT98), .B(n378), .Z(n345) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n348) );
  XOR2_X1 U397 ( .A(G64GAT), .B(G211GAT), .Z(n347) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n396) );
  XOR2_X1 U400 ( .A(n348), .B(n396), .Z(n352) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U402 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U403 ( .A(n450), .B(n353), .Z(n526) );
  XOR2_X1 U404 ( .A(KEYINPUT122), .B(n526), .Z(n417) );
  XOR2_X1 U405 ( .A(G141GAT), .B(G22GAT), .Z(n355) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G15GAT), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U408 ( .A(KEYINPUT67), .B(KEYINPUT71), .Z(n357) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G1GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U412 ( .A(KEYINPUT70), .B(G8GAT), .Z(n361) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U415 ( .A(KEYINPUT30), .B(n362), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U417 ( .A(G50GAT), .B(G36GAT), .Z(n367) );
  XNOR2_X1 U418 ( .A(n365), .B(G113GAT), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U420 ( .A(n369), .B(n368), .Z(n374) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n371) );
  XNOR2_X1 U422 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n372), .B(G43GAT), .ZN(n373) );
  XOR2_X1 U425 ( .A(n374), .B(n373), .Z(n556) );
  INV_X1 U426 ( .A(n556), .ZN(n581) );
  XOR2_X1 U427 ( .A(KEYINPUT13), .B(G57GAT), .Z(n376) );
  XNOR2_X1 U428 ( .A(G71GAT), .B(G78GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n397) );
  XNOR2_X1 U430 ( .A(n377), .B(n397), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U432 ( .A(n380), .B(KEYINPUT33), .Z(n382) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U435 ( .A(n384), .B(n383), .Z(n392) );
  XOR2_X1 U436 ( .A(G64GAT), .B(G92GAT), .Z(n386) );
  XNOR2_X1 U437 ( .A(G176GAT), .B(G120GAT), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U439 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n388) );
  XNOR2_X1 U440 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n392), .B(n391), .ZN(n585) );
  NAND2_X1 U444 ( .A1(n581), .A2(n585), .ZN(n409) );
  XOR2_X1 U445 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n394) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U448 ( .A(n395), .B(KEYINPUT83), .Z(n399) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U451 ( .A(KEYINPUT84), .B(KEYINPUT15), .Z(n401) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(KEYINPUT85), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U454 ( .A(n403), .B(n402), .Z(n406) );
  XOR2_X1 U455 ( .A(G15GAT), .B(G127GAT), .Z(n453) );
  XNOR2_X1 U456 ( .A(n453), .B(n404), .ZN(n405) );
  XOR2_X1 U457 ( .A(n406), .B(n405), .Z(n562) );
  INV_X1 U458 ( .A(n562), .ZN(n589) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(n548), .ZN(n592) );
  NOR2_X1 U460 ( .A1(n589), .A2(n592), .ZN(n407) );
  XOR2_X1 U461 ( .A(n407), .B(KEYINPUT45), .Z(n408) );
  NOR2_X1 U462 ( .A1(n409), .A2(n408), .ZN(n415) );
  XOR2_X1 U463 ( .A(n562), .B(KEYINPUT116), .Z(n576) );
  NAND2_X1 U464 ( .A1(n565), .A2(n576), .ZN(n412) );
  XNOR2_X1 U465 ( .A(n585), .B(KEYINPUT41), .ZN(n558) );
  INV_X1 U466 ( .A(n558), .ZN(n572) );
  NOR2_X1 U467 ( .A1(n581), .A2(n572), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n410), .B(KEYINPUT46), .ZN(n411) );
  OR2_X1 U469 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U470 ( .A(KEYINPUT47), .B(n413), .ZN(n414) );
  NOR2_X1 U471 ( .A1(n415), .A2(n414), .ZN(n416) );
  XOR2_X1 U472 ( .A(KEYINPUT48), .B(n416), .Z(n553) );
  NAND2_X1 U473 ( .A1(n417), .A2(n553), .ZN(n420) );
  XNOR2_X1 U474 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n418) );
  XOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n422) );
  XNOR2_X1 U476 ( .A(KEYINPUT94), .B(G57GAT), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n427) );
  XNOR2_X1 U478 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(G120GAT), .ZN(n455) );
  XOR2_X1 U480 ( .A(n455), .B(KEYINPUT1), .Z(n425) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U484 ( .A(KEYINPUT96), .B(G148GAT), .Z(n429) );
  XNOR2_X1 U485 ( .A(G127GAT), .B(G155GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U487 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n431) );
  XNOR2_X1 U488 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U490 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U491 ( .A(G85GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U492 ( .A(G134GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(G29GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n552) );
  NAND2_X1 U497 ( .A1(n442), .A2(n552), .ZN(n578) );
  XNOR2_X1 U498 ( .A(KEYINPUT55), .B(n443), .ZN(n459) );
  XOR2_X1 U499 ( .A(G183GAT), .B(G71GAT), .Z(n445) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n446), .B(KEYINPUT87), .Z(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n448) );
  XNOR2_X1 U504 ( .A(G190GAT), .B(G99GAT), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n454) );
  XOR2_X1 U508 ( .A(n454), .B(n453), .Z(n458) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U510 ( .A(n458), .B(n457), .Z(n466) );
  BUF_X1 U511 ( .A(n466), .Z(n536) );
  NOR2_X1 U512 ( .A1(n459), .A2(n536), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT125), .ZN(n575) );
  NOR2_X1 U514 ( .A1(n548), .A2(n575), .ZN(n463) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n585), .A2(n556), .ZN(n497) );
  NOR2_X1 U517 ( .A1(n526), .A2(n466), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n472), .A2(n464), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n465), .B(KEYINPUT25), .ZN(n469) );
  XOR2_X1 U520 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n468) );
  NAND2_X1 U521 ( .A1(n472), .A2(n466), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n468), .B(n467), .ZN(n579) );
  XOR2_X1 U523 ( .A(KEYINPUT27), .B(n526), .Z(n475) );
  NAND2_X1 U524 ( .A1(n579), .A2(n475), .ZN(n551) );
  NAND2_X1 U525 ( .A1(n469), .A2(n551), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT101), .B(n470), .Z(n471) );
  NAND2_X1 U527 ( .A1(n471), .A2(n552), .ZN(n479) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT66), .ZN(n491) );
  XNOR2_X1 U529 ( .A(n491), .B(KEYINPUT28), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n552), .A2(n473), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n535) );
  XNOR2_X1 U532 ( .A(KEYINPUT99), .B(n535), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n536), .B(KEYINPUT90), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(KEYINPUT102), .ZN(n494) );
  XOR2_X1 U537 ( .A(KEYINPUT86), .B(KEYINPUT16), .Z(n482) );
  NAND2_X1 U538 ( .A1(n548), .A2(n562), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n494), .A2(n483), .ZN(n510) );
  OR2_X1 U541 ( .A1(n497), .A2(n510), .ZN(n492) );
  NOR2_X1 U542 ( .A1(n552), .A2(n492), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT103), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n526), .A2(n492), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT104), .B(n487), .Z(n488) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U549 ( .A1(n536), .A2(n492), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  XOR2_X1 U552 ( .A(n491), .B(KEYINPUT28), .Z(n532) );
  NOR2_X1 U553 ( .A1(n532), .A2(n492), .ZN(n493) );
  XOR2_X1 U554 ( .A(G22GAT), .B(n493), .Z(G1327GAT) );
  XNOR2_X1 U555 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n589), .A2(n494), .ZN(n495) );
  NOR2_X1 U557 ( .A1(n592), .A2(n495), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n496), .ZN(n522) );
  NOR2_X1 U559 ( .A1(n522), .A2(n497), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT105), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT38), .ZN(n508) );
  NOR2_X1 U562 ( .A1(n552), .A2(n508), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n504) );
  NOR2_X1 U566 ( .A1(n526), .A2(n508), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NOR2_X1 U568 ( .A1(n508), .A2(n536), .ZN(n506) );
  XNOR2_X1 U569 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U571 ( .A(G43GAT), .B(n507), .Z(G1330GAT) );
  NOR2_X1 U572 ( .A1(n508), .A2(n532), .ZN(n509) );
  XOR2_X1 U573 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  NAND2_X1 U574 ( .A1(n581), .A2(n558), .ZN(n521) );
  NOR2_X1 U575 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(KEYINPUT109), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n552), .A2(n518), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U580 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n518), .ZN(n515) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n536), .A2(n518), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n532), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n531) );
  NOR2_X1 U590 ( .A1(n552), .A2(n531), .ZN(n524) );
  XNOR2_X1 U591 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n531), .ZN(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n536), .A2(n531), .ZN(n530) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n537), .A2(n553), .ZN(n538) );
  XOR2_X1 U605 ( .A(n538), .B(KEYINPUT117), .Z(n547) );
  INV_X1 U606 ( .A(n547), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n556), .A2(n541), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n539), .B(KEYINPUT118), .ZN(n540) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U611 ( .A1(n541), .A2(n558), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U613 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  NOR2_X1 U614 ( .A1(n576), .A2(n547), .ZN(n545) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(n545), .Z(n546) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  NOR2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT120), .B(n555), .ZN(n566) );
  INV_X1 U623 ( .A(n566), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n563), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U627 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n581), .A2(n575), .ZN(n569) );
  XOR2_X1 U636 ( .A(G169GAT), .B(n569), .Z(G1348GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n571) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT126), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n574) );
  NOR2_X1 U640 ( .A1(n572), .A2(n575), .ZN(n573) );
  XOR2_X1 U641 ( .A(n574), .B(n573), .Z(G1349GAT) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G183GAT), .B(n577), .Z(G1350GAT) );
  INV_X1 U644 ( .A(n578), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n591) );
  NOR2_X1 U646 ( .A1(n581), .A2(n591), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(n584), .ZN(G1352GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n591), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U653 ( .A(G204GAT), .B(n588), .Z(G1353GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n591), .ZN(n590) );
  XOR2_X1 U655 ( .A(G211GAT), .B(n590), .Z(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

