//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(G134gat), .B(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT15), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(G50gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n207), .A2(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n208), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT91), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n206), .B1(new_n221), .B2(new_n204), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n203), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(KEYINPUT17), .B(new_n213), .C1(new_n220), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT92), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT15), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n229), .A2(new_n217), .A3(new_n219), .A4(new_n214), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT17), .A4(new_n213), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT7), .ZN(new_n235));
  NOR2_X1   g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(KEYINPUT8), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT100), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n237), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n243), .A3(new_n238), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n244), .A2(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n213), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT102), .ZN(new_n252));
  AND2_X1   g051(.A1(G232gat), .A2(G233gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n249), .A2(new_n247), .B1(KEYINPUT41), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n251), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n202), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(new_n202), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G190gat), .B(G218gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT101), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n253), .A2(KEYINPUT41), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n261), .A3(new_n266), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(G71gat), .A2(G78gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  XOR2_X1   g071(.A(G57gat), .B(G64gat), .Z(new_n273));
  AOI211_X1 g072(.A(new_n271), .B(new_n272), .C1(new_n273), .C2(KEYINPUT9), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(KEYINPUT9), .B2(new_n272), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT98), .B(G57gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G64gat), .ZN(new_n277));
  INV_X1    g076(.A(G64gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G57gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(KEYINPUT21), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G155gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT16), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(G1gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G1gat), .B2(new_n285), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G8gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(KEYINPUT21), .B2(new_n281), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n284), .B(new_n290), .Z(new_n291));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT99), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n291), .B(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n270), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT103), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n247), .B2(new_n281), .ZN(new_n301));
  INV_X1    g100(.A(new_n281), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n302), .A2(new_n245), .A3(KEYINPUT103), .A4(new_n246), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n281), .A2(new_n244), .A3(new_n241), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G230gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT104), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n301), .A2(new_n310), .A3(new_n303), .A4(new_n304), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n281), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n306), .ZN(new_n314));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(KEYINPUT104), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n309), .A2(new_n314), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(new_n308), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT105), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G169gat), .B(G197gat), .Z(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT89), .ZN(new_n330));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT88), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n330), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT12), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n289), .B1(new_n249), .B2(new_n248), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n233), .A2(new_n337), .B1(new_n249), .B2(new_n289), .ZN(new_n338));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT93), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT18), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT97), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(KEYINPUT18), .A3(new_n340), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n288), .B(G8gat), .Z(new_n347));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n213), .A4(new_n230), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT95), .B1(new_n249), .B2(new_n289), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n249), .A2(new_n289), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT96), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n340), .B(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n355), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT96), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n343), .A2(new_n346), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n345), .B(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n299), .A2(KEYINPUT105), .A3(new_n325), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n328), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT35), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT27), .B(G183gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G183gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT27), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G183gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT67), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n371), .B2(new_n373), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(KEYINPUT28), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n369), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT68), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  INV_X1    g185(.A(G169gat), .ZN(new_n387));
  INV_X1    g186(.A(G176gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT65), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(G169gat), .B2(G176gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(KEYINPUT24), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G183gat), .B(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT24), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT23), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n382), .A2(KEYINPUT64), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT23), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(G169gat), .B2(G176gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(G169gat), .A3(G176gat), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n403), .A2(new_n405), .A3(new_n407), .A4(KEYINPUT25), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n401), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n370), .A2(G190gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n367), .A2(G183gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n397), .B1(new_n412), .B2(KEYINPUT24), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT23), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n405), .A3(new_n382), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT25), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n380), .A2(new_n396), .B1(new_n409), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G127gat), .B(G134gat), .Z(new_n419));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(KEYINPUT1), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G120gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G113gat), .ZN(new_n423));
  INV_X1    g222(.A(G113gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G120gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G127gat), .B(G134gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT1), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n395), .B(new_n394), .C1(new_n432), .C2(new_n369), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n428), .B2(new_n426), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT25), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n401), .B2(new_n415), .ZN(new_n438));
  INV_X1    g237(.A(new_n408), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT23), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n413), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n365), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n364), .B1(new_n444), .B2(KEYINPUT33), .ZN(new_n445));
  XNOR2_X1  g244(.A(G15gat), .B(G43gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n365), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n433), .A2(new_n436), .A3(new_n442), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n436), .B1(new_n433), .B2(new_n442), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n448), .B1(new_n452), .B2(KEYINPUT32), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(KEYINPUT69), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n445), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT70), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT70), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n445), .A2(new_n453), .A3(new_n458), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n448), .A2(new_n454), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n431), .A2(new_n466), .A3(new_n365), .A4(new_n443), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT71), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n431), .A2(new_n365), .A3(new_n443), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT34), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(G22gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G228gat), .ZN(new_n477));
  INV_X1    g276(.A(G233gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT2), .ZN(new_n480));
  INV_X1    g279(.A(G155gat), .ZN(new_n481));
  INV_X1    g280(.A(G162gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n487));
  INV_X1    g286(.A(G148gat), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(G141gat), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n481), .A2(new_n482), .ZN(new_n493));
  XNOR2_X1  g292(.A(G141gat), .B(G148gat), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n484), .B(new_n493), .C1(new_n494), .C2(KEYINPUT2), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G197gat), .B(G204gat), .ZN(new_n497));
  AND2_X1   g296(.A1(G211gat), .A2(G218gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(KEYINPUT22), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(G211gat), .A2(G218gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n498), .A2(KEYINPUT22), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n503), .B(new_n497), .C1(new_n498), .C2(new_n500), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT29), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n505), .B2(new_n506), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n496), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n502), .A2(new_n504), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT72), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n508), .A3(new_n495), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n512), .A2(KEYINPUT85), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT85), .B1(new_n512), .B2(new_n515), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n479), .B(new_n510), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  OR2_X1    g317(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(G148gat), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n521), .A2(new_n490), .B1(new_n484), .B2(new_n483), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n493), .A2(new_n484), .ZN(new_n523));
  INV_X1    g322(.A(G141gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G148gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n490), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n480), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT83), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(new_n514), .C1(KEYINPUT83), .C2(new_n504), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n528), .B1(new_n530), .B2(new_n508), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n531), .A2(new_n532), .B1(new_n477), .B2(new_n478), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT31), .B(G50gat), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n518), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n518), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n476), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n534), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n533), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n475), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n472), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n460), .A2(new_n464), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n473), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n394), .A2(new_n395), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n371), .A2(new_n373), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT67), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n368), .A2(new_n374), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(new_n379), .ZN(new_n551));
  INV_X1    g350(.A(new_n366), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G190gat), .B2(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n547), .A2(new_n554), .B1(new_n438), .B2(new_n441), .ZN(new_n555));
  NAND2_X1  g354(.A1(G226gat), .A2(G233gat), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT75), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT75), .ZN(new_n558));
  INV_X1    g357(.A(new_n556), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n418), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT74), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n433), .A2(new_n563), .A3(new_n442), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT29), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n561), .B(new_n511), .C1(new_n565), .C2(new_n559), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n559), .A3(new_n564), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n418), .A2(new_n514), .A3(new_n556), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n512), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G8gat), .B(G36gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G64gat), .B(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n566), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT78), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(KEYINPUT78), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G1gat), .B(G29gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT0), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G85gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT3), .B1(new_n522), .B2(new_n527), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n513), .A3(new_n430), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n492), .A2(new_n495), .A3(new_n421), .A4(new_n429), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT4), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n528), .A2(new_n436), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G225gat), .A2(G233gat), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n587), .A2(new_n590), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT5), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI22_X1  g396(.A1(new_n522), .A2(new_n527), .B1(new_n434), .B2(new_n435), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT81), .A3(new_n588), .ZN(new_n599));
  INV_X1    g398(.A(new_n593), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT81), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n496), .A2(new_n601), .A3(new_n430), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n588), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n587), .B2(new_n591), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT5), .B(new_n593), .C1(new_n588), .C2(new_n589), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n585), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n587), .A2(new_n591), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(new_n585), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n596), .A3(new_n603), .A4(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT6), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n597), .A2(new_n607), .A3(new_n585), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT82), .B1(new_n616), .B2(KEYINPUT6), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT82), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n613), .A2(new_n618), .A3(new_n614), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n615), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n575), .B1(new_n566), .B2(new_n569), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n566), .A2(new_n569), .A3(new_n575), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(KEYINPUT30), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n581), .A2(KEYINPUT86), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n363), .B1(new_n546), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n576), .A2(KEYINPUT78), .A3(new_n577), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n623), .B(new_n620), .C1(new_n626), .C2(new_n578), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT86), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n544), .B1(new_n460), .B2(new_n464), .ZN(new_n630));
  AOI211_X1 g429(.A(new_n463), .B(new_n472), .C1(new_n457), .C2(new_n459), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n629), .A2(KEYINPUT35), .A3(new_n543), .A4(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n473), .A2(new_n634), .A3(new_n545), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT36), .B1(new_n630), .B2(new_n631), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n538), .A2(new_n542), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n627), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n623), .B1(new_n626), .B2(new_n578), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n600), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n599), .A2(new_n602), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n642), .B(KEYINPUT39), .C1(new_n600), .C2(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n644), .B(new_n585), .C1(KEYINPUT39), .C2(new_n642), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n647), .A2(new_n648), .A3(new_n616), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n566), .A2(new_n651), .A3(new_n569), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n574), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n566), .B2(new_n569), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT38), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT29), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n433), .A2(new_n563), .A3(new_n442), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n563), .B1(new_n433), .B2(new_n442), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n556), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n511), .B1(new_n660), .B2(new_n561), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n512), .B1(new_n567), .B2(new_n568), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT37), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n574), .A4(new_n652), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n618), .B1(new_n613), .B2(new_n614), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n616), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n616), .A2(KEYINPUT6), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n666), .A2(new_n667), .B1(new_n668), .B2(new_n608), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n655), .A2(new_n665), .A3(new_n669), .A4(new_n576), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n650), .A2(new_n543), .A3(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n625), .B(new_n633), .C1(new_n639), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n362), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n669), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n640), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n640), .ZN(new_n679));
  OAI21_X1  g478(.A(G8gat), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g480(.A(new_n678), .B(new_n681), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g481(.A1(new_n635), .A2(new_n636), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n673), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n632), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n673), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n543), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  AND2_X1   g490(.A1(new_n672), .A2(new_n270), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT12), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n335), .B(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT18), .B1(new_n338), .B2(new_n340), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(KEYINPUT97), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n359), .B(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n298), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(new_n698), .A3(new_n324), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n692), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n210), .A3(new_n669), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n672), .A2(new_n704), .A3(new_n270), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n672), .A2(new_n704), .A3(KEYINPUT44), .A4(new_n270), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n699), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n620), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n710), .B2(new_n679), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n701), .A2(new_n211), .A3(new_n640), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n713), .B(new_n717), .C1(new_n715), .C2(new_n714), .ZN(G1329gat));
  NOR3_X1   g517(.A1(new_n700), .A2(G43gat), .A3(new_n686), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n683), .A3(new_n699), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(G43gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n700), .B2(new_n543), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n543), .A2(new_n723), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n710), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g527(.A1(new_n672), .A2(new_n697), .A3(new_n299), .A4(new_n324), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n669), .B(KEYINPUT108), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n276), .ZN(G1332gat));
  XNOR2_X1  g531(.A(new_n729), .B(KEYINPUT109), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n679), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n733), .B2(new_n684), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n729), .A2(G71gat), .A3(new_n686), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n733), .A2(new_n543), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g544(.A1(new_n360), .A2(new_n698), .A3(new_n325), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n709), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n620), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n360), .A2(new_n698), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n672), .A2(new_n270), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n672), .A2(KEYINPUT51), .A3(new_n270), .A4(new_n749), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n750), .A2(KEYINPUT111), .A3(new_n751), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n620), .A2(G85gat), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n755), .A2(new_n324), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n748), .A2(new_n758), .ZN(G1336gat));
  NOR3_X1   g558(.A1(new_n679), .A2(G92gat), .A3(new_n325), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n707), .A2(new_n640), .A3(new_n708), .A4(new_n746), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n752), .A2(new_n754), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n760), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT112), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n762), .A2(G92gat), .B1(new_n766), .B2(new_n760), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n770), .B(new_n771), .C1(new_n764), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(G1337gat));
  OAI21_X1  g573(.A(G99gat), .B1(new_n747), .B2(new_n684), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n686), .A2(G99gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n755), .A2(new_n324), .A3(new_n756), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n709), .A2(new_n637), .A3(new_n746), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G106gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n543), .A2(new_n325), .A3(G106gat), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n755), .A2(new_n756), .A3(new_n783), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n779), .A2(G106gat), .B1(new_n766), .B2(new_n783), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n782), .A2(new_n784), .B1(new_n785), .B2(new_n781), .ZN(G1339gat));
  NAND3_X1  g585(.A1(new_n299), .A2(new_n697), .A3(new_n325), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n338), .A2(new_n340), .B1(new_n352), .B2(new_n355), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n335), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n324), .B(new_n789), .C1(new_n694), .C2(new_n359), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n314), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n317), .B1(new_n322), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n794), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n319), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n790), .B1(new_n697), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n270), .ZN(new_n801));
  INV_X1    g600(.A(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n789), .B1(new_n359), .B2(new_n694), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n268), .B2(new_n269), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n787), .B1(new_n805), .B2(new_n698), .ZN(new_n806));
  INV_X1    g605(.A(new_n730), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n806), .A2(new_n543), .A3(new_n632), .A4(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n640), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n787), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n800), .A2(new_n801), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n804), .A2(new_n802), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n814), .B2(new_n298), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n546), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT113), .A3(new_n807), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n360), .A2(new_n424), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(new_n669), .A3(new_n679), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n697), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1340gat));
  NOR3_X1   g623(.A1(new_n822), .A2(new_n422), .A3(new_n325), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n324), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n422), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n818), .A2(new_n828), .A3(new_n698), .ZN(new_n829));
  OAI21_X1  g628(.A(G127gat), .B1(new_n822), .B2(new_n298), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1342gat));
  NOR2_X1   g630(.A1(new_n801), .A2(G134gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n817), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT115), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n822), .B2(new_n801), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n815), .A2(new_n543), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n683), .A2(new_n640), .A3(new_n730), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(G141gat), .A3(new_n697), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(KEYINPUT58), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n486), .A2(new_n487), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n683), .A2(new_n620), .A3(new_n640), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n806), .B2(new_n637), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n637), .A2(KEYINPUT57), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n798), .A2(new_n319), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n795), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n792), .A2(KEYINPUT116), .A3(new_n794), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n796), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n360), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n270), .B1(new_n856), .B2(new_n790), .ZN(new_n857));
  INV_X1    g656(.A(new_n813), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n298), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n850), .B1(new_n859), .B2(new_n787), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n848), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n847), .B1(new_n861), .B2(new_n697), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT117), .B(new_n848), .C1(new_n849), .C2(new_n860), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n360), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n844), .B1(new_n867), .B2(new_n847), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(G1344gat));
  NOR3_X1   g669(.A1(new_n843), .A2(G148gat), .A3(new_n325), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT118), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n324), .A3(new_n866), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n488), .A2(KEYINPUT59), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n543), .A2(KEYINPUT57), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n328), .A2(new_n697), .A3(new_n361), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n790), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n801), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n698), .B1(new_n879), .B2(new_n813), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT57), .B1(new_n815), .B2(new_n543), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n848), .A2(new_n324), .ZN(new_n884));
  OAI21_X1  g683(.A(G148gat), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n875), .B2(new_n886), .ZN(G1345gat));
  INV_X1    g686(.A(new_n843), .ZN(new_n888));
  AOI21_X1  g687(.A(G155gat), .B1(new_n888), .B2(new_n698), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n865), .A2(new_n866), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n298), .A2(new_n481), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT119), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n888), .B2(new_n270), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n801), .A2(new_n482), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n890), .B2(new_n895), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n807), .A2(new_n679), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n816), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n387), .A3(new_n697), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n815), .B2(new_n669), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n806), .A2(KEYINPUT120), .A3(new_n620), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n546), .A2(new_n679), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n360), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n899), .B1(new_n906), .B2(new_n387), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n388), .A3(new_n324), .ZN(new_n908));
  OAI21_X1  g707(.A(G176gat), .B1(new_n898), .B2(new_n325), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n898), .B2(new_n298), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n298), .A2(new_n376), .A3(new_n375), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n903), .A2(new_n904), .A3(new_n913), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT60), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n905), .A2(new_n367), .A3(new_n270), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n898), .B2(new_n801), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  XNOR2_X1  g721(.A(KEYINPUT123), .B(G197gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n683), .A2(new_n807), .A3(new_n679), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n881), .A2(new_n882), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(new_n697), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n683), .A2(new_n679), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n637), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n901), .A2(new_n902), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n697), .A2(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n930), .A2(new_n929), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n325), .A2(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n903), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n931), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n925), .B2(new_n325), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(KEYINPUT62), .A3(new_n942), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G1353gat));
  NAND4_X1  g747(.A1(new_n881), .A2(new_n882), .A3(new_n698), .A4(new_n924), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n298), .A2(G211gat), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n950), .A2(new_n951), .B1(new_n931), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n950), .A2(new_n951), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n949), .A2(G211gat), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n954), .B2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n925), .B2(new_n801), .ZN(new_n959));
  INV_X1    g758(.A(new_n931), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n801), .A2(G218gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(G1355gat));
endmodule


