

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G2104), .A2(n537), .ZN(n890) );
  NOR2_X2 U554 ( .A1(G2105), .A2(n538), .ZN(n573) );
  XNOR2_X2 U555 ( .A(KEYINPUT67), .B(n547), .ZN(n594) );
  XOR2_X1 U556 ( .A(KEYINPUT29), .B(KEYINPUT100), .Z(n523) );
  XOR2_X1 U557 ( .A(KEYINPUT66), .B(n539), .Z(n524) );
  OR2_X1 U558 ( .A1(n723), .A2(G301), .ZN(n525) );
  XNOR2_X1 U559 ( .A(n694), .B(KEYINPUT26), .ZN(n698) );
  AND2_X1 U560 ( .A1(n722), .A2(n525), .ZN(n732) );
  NOR2_X1 U561 ( .A1(n732), .A2(n731), .ZN(n742) );
  AND2_X1 U562 ( .A1(G40), .A2(n693), .ZN(n802) );
  NOR2_X1 U563 ( .A1(n538), .A2(n537), .ZN(n891) );
  NOR2_X1 U564 ( .A1(G651), .A2(n651), .ZN(n659) );
  INV_X1 U565 ( .A(G2104), .ZN(n538) );
  NAND2_X1 U566 ( .A1(n573), .A2(G101), .ZN(n526) );
  XOR2_X1 U567 ( .A(n526), .B(KEYINPUT23), .Z(n528) );
  INV_X1 U568 ( .A(G2105), .ZN(n537) );
  NAND2_X1 U569 ( .A1(n890), .A2(G125), .ZN(n527) );
  NAND2_X1 U570 ( .A1(n528), .A2(n527), .ZN(n531) );
  INV_X1 U571 ( .A(n531), .ZN(n530) );
  INV_X1 U572 ( .A(KEYINPUT65), .ZN(n529) );
  NAND2_X1 U573 ( .A1(n530), .A2(n529), .ZN(n533) );
  NAND2_X1 U574 ( .A1(n531), .A2(KEYINPUT65), .ZN(n532) );
  NAND2_X1 U575 ( .A1(n533), .A2(n532), .ZN(n536) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n534), .Z(n894) );
  NAND2_X1 U578 ( .A1(G137), .A2(n894), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U580 ( .A1(n891), .A2(G113), .ZN(n539) );
  NOR2_X1 U581 ( .A1(n540), .A2(n524), .ZN(n541) );
  XNOR2_X1 U582 ( .A(KEYINPUT64), .B(n541), .ZN(n693) );
  BUF_X1 U583 ( .A(n693), .Z(G160) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n651) );
  NAND2_X1 U585 ( .A1(n659), .A2(G52), .ZN(n545) );
  INV_X1 U586 ( .A(G651), .ZN(n546) );
  NOR2_X1 U587 ( .A1(G543), .A2(n546), .ZN(n542) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n542), .Z(n543) );
  XNOR2_X1 U589 ( .A(KEYINPUT68), .B(n543), .ZN(n662) );
  NAND2_X1 U590 ( .A1(G64), .A2(n662), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n545), .A2(n544), .ZN(n552) );
  NOR2_X1 U592 ( .A1(G651), .A2(G543), .ZN(n658) );
  NAND2_X1 U593 ( .A1(G90), .A2(n658), .ZN(n549) );
  OR2_X1 U594 ( .A1(n546), .A2(n651), .ZN(n547) );
  NAND2_X1 U595 ( .A1(G77), .A2(n594), .ZN(n548) );
  NAND2_X1 U596 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U597 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U598 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(G88), .A2(n658), .ZN(n554) );
  NAND2_X1 U604 ( .A1(G75), .A2(n594), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U606 ( .A1(n659), .A2(G50), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G62), .A2(n662), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U609 ( .A1(n558), .A2(n557), .ZN(G166) );
  XNOR2_X1 U610 ( .A(KEYINPUT78), .B(KEYINPUT6), .ZN(n563) );
  NAND2_X1 U611 ( .A1(n659), .A2(G51), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G63), .A2(n662), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT77), .B(n559), .Z(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U615 ( .A(n563), .B(n562), .Z(n570) );
  XNOR2_X1 U616 ( .A(KEYINPUT76), .B(KEYINPUT5), .ZN(n568) );
  NAND2_X1 U617 ( .A1(n658), .A2(G89), .ZN(n564) );
  XNOR2_X1 U618 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G76), .A2(n594), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U621 ( .A(n568), .B(n567), .ZN(n569) );
  NAND2_X1 U622 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U623 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .ZN(n572) );
  XNOR2_X1 U625 ( .A(n572), .B(KEYINPUT79), .ZN(G286) );
  NAND2_X1 U626 ( .A1(G138), .A2(n894), .ZN(n575) );
  NAND2_X1 U627 ( .A1(G102), .A2(n573), .ZN(n574) );
  NAND2_X1 U628 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U629 ( .A1(G126), .A2(n890), .ZN(n577) );
  NAND2_X1 U630 ( .A1(G114), .A2(n891), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U632 ( .A1(n579), .A2(n578), .ZN(G164) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U634 ( .A(n580), .B(KEYINPUT10), .ZN(n581) );
  XNOR2_X1 U635 ( .A(KEYINPUT72), .B(n581), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n839) );
  NAND2_X1 U637 ( .A1(n839), .A2(G567), .ZN(n582) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U639 ( .A1(n662), .A2(G56), .ZN(n583) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U641 ( .A1(n658), .A2(G81), .ZN(n584) );
  XNOR2_X1 U642 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U643 ( .A1(G68), .A2(n594), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U646 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n659), .A2(G43), .ZN(n590) );
  NAND2_X1 U648 ( .A1(n591), .A2(n590), .ZN(n1011) );
  XNOR2_X1 U649 ( .A(G860), .B(KEYINPUT73), .ZN(n615) );
  OR2_X1 U650 ( .A1(n1011), .A2(n615), .ZN(G153) );
  NAND2_X1 U651 ( .A1(G868), .A2(G171), .ZN(n602) );
  NAND2_X1 U652 ( .A1(G66), .A2(n662), .ZN(n599) );
  NAND2_X1 U653 ( .A1(G92), .A2(n658), .ZN(n593) );
  NAND2_X1 U654 ( .A1(G54), .A2(n659), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U656 ( .A1(n594), .A2(G79), .ZN(n595) );
  XOR2_X1 U657 ( .A(KEYINPUT74), .B(n595), .Z(n596) );
  NOR2_X1 U658 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U659 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n600), .Z(n1024) );
  INV_X1 U661 ( .A(n1024), .ZN(n636) );
  INV_X1 U662 ( .A(G868), .ZN(n676) );
  NAND2_X1 U663 ( .A1(n636), .A2(n676), .ZN(n601) );
  NAND2_X1 U664 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U665 ( .A(n603), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G91), .A2(n658), .ZN(n604) );
  XNOR2_X1 U667 ( .A(n604), .B(KEYINPUT70), .ZN(n611) );
  NAND2_X1 U668 ( .A1(n659), .A2(G53), .ZN(n606) );
  NAND2_X1 U669 ( .A1(G65), .A2(n662), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U671 ( .A1(G78), .A2(n594), .ZN(n607) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(n607), .ZN(n608) );
  NOR2_X1 U673 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n611), .A2(n610), .ZN(G299) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n612) );
  XNOR2_X1 U676 ( .A(n612), .B(KEYINPUT80), .ZN(n614) );
  NOR2_X1 U677 ( .A1(n676), .A2(G286), .ZN(n613) );
  NOR2_X1 U678 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n615), .A2(G559), .ZN(n616) );
  NAND2_X1 U680 ( .A1(n616), .A2(n636), .ZN(n617) );
  XNOR2_X1 U681 ( .A(n617), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n1011), .ZN(n620) );
  NAND2_X1 U683 ( .A1(G868), .A2(n636), .ZN(n618) );
  NOR2_X1 U684 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U685 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U686 ( .A1(G123), .A2(n890), .ZN(n621) );
  XNOR2_X1 U687 ( .A(n621), .B(KEYINPUT18), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n573), .A2(G99), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U690 ( .A1(G135), .A2(n894), .ZN(n625) );
  NAND2_X1 U691 ( .A1(G111), .A2(n891), .ZN(n624) );
  NAND2_X1 U692 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U693 ( .A1(n627), .A2(n626), .ZN(n982) );
  XNOR2_X1 U694 ( .A(n982), .B(G2096), .ZN(n629) );
  INV_X1 U695 ( .A(G2100), .ZN(n628) );
  NAND2_X1 U696 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U697 ( .A1(n658), .A2(G93), .ZN(n631) );
  NAND2_X1 U698 ( .A1(G67), .A2(n662), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U700 ( .A1(G80), .A2(n594), .ZN(n633) );
  NAND2_X1 U701 ( .A1(G55), .A2(n659), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n677) );
  NAND2_X1 U704 ( .A1(G559), .A2(n636), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n1011), .B(n637), .ZN(n674) );
  NOR2_X1 U706 ( .A1(G860), .A2(n674), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT81), .B(n638), .Z(n639) );
  XOR2_X1 U708 ( .A(n677), .B(n639), .Z(G145) );
  NAND2_X1 U709 ( .A1(n658), .A2(G86), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(KEYINPUT84), .ZN(n642) );
  NAND2_X1 U711 ( .A1(G61), .A2(n662), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(KEYINPUT85), .ZN(n645) );
  NAND2_X1 U714 ( .A1(G48), .A2(n659), .ZN(n644) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U716 ( .A1(n594), .A2(G73), .ZN(n646) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U719 ( .A(KEYINPUT86), .B(n649), .Z(G305) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT82), .ZN(n654) );
  NAND2_X1 U722 ( .A1(G87), .A2(n651), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT83), .B(n652), .Z(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n662), .A2(n655), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n659), .A2(G49), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G85), .A2(n658), .ZN(n661) );
  NAND2_X1 U729 ( .A1(G47), .A2(n659), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n594), .A2(G72), .ZN(n664) );
  NAND2_X1 U732 ( .A1(G60), .A2(n662), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT69), .ZN(G290) );
  XOR2_X1 U736 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n668) );
  XNOR2_X1 U737 ( .A(G288), .B(n668), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(n677), .ZN(n671) );
  INV_X1 U739 ( .A(G299), .ZN(n714) );
  XNOR2_X1 U740 ( .A(G166), .B(n714), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U742 ( .A(G305), .B(n672), .Z(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(G290), .ZN(n909) );
  XNOR2_X1 U744 ( .A(n909), .B(n674), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n679) );
  NOR2_X1 U746 ( .A1(G868), .A2(n677), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(KEYINPUT88), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U753 ( .A1(G2072), .A2(n684), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U757 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U758 ( .A1(G96), .A2(n687), .ZN(n844) );
  NAND2_X1 U759 ( .A1(n844), .A2(G2106), .ZN(n691) );
  NAND2_X1 U760 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U761 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U762 ( .A1(G108), .A2(n689), .ZN(n845) );
  NAND2_X1 U763 ( .A1(n845), .A2(G567), .ZN(n690) );
  NAND2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n846) );
  NAND2_X1 U765 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U766 ( .A1(n846), .A2(n692), .ZN(n843) );
  NAND2_X1 U767 ( .A1(n843), .A2(G36), .ZN(G176) );
  INV_X1 U768 ( .A(G166), .ZN(G303) );
  INV_X1 U769 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U770 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n838) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n804) );
  NAND2_X1 U772 ( .A1(n804), .A2(n802), .ZN(n745) );
  NAND2_X1 U773 ( .A1(G8), .A2(n745), .ZN(n773) );
  NOR2_X1 U774 ( .A1(G1966), .A2(n773), .ZN(n733) );
  AND2_X2 U775 ( .A1(n804), .A2(n802), .ZN(n719) );
  NAND2_X1 U776 ( .A1(n719), .A2(G1996), .ZN(n694) );
  NAND2_X1 U777 ( .A1(G1341), .A2(n745), .ZN(n696) );
  INV_X1 U778 ( .A(n1011), .ZN(n695) );
  AND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U780 ( .A1(n698), .A2(n697), .ZN(n705) );
  NOR2_X1 U781 ( .A1(n705), .A2(n1024), .ZN(n699) );
  XOR2_X1 U782 ( .A(KEYINPUT98), .B(n699), .Z(n704) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n745), .ZN(n701) );
  NAND2_X1 U784 ( .A1(G2067), .A2(n719), .ZN(n700) );
  NAND2_X1 U785 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U786 ( .A(KEYINPUT99), .B(n702), .Z(n703) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U788 ( .A1(n705), .A2(n1024), .ZN(n706) );
  NAND2_X1 U789 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U790 ( .A1(n719), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U791 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U792 ( .A(G1956), .ZN(n939) );
  NOR2_X1 U793 ( .A1(n719), .A2(n939), .ZN(n709) );
  NOR2_X1 U794 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U795 ( .A1(n714), .A2(n713), .ZN(n711) );
  NAND2_X1 U796 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U797 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U798 ( .A(n715), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U799 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U800 ( .A(n718), .B(n523), .ZN(n722) );
  XOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .Z(n963) );
  NOR2_X1 U802 ( .A1(n963), .A2(n745), .ZN(n721) );
  XOR2_X1 U803 ( .A(G1961), .B(KEYINPUT97), .Z(n935) );
  NOR2_X1 U804 ( .A1(n719), .A2(n935), .ZN(n720) );
  NOR2_X1 U805 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U806 ( .A1(n723), .A2(G301), .ZN(n724) );
  XNOR2_X1 U807 ( .A(n724), .B(KEYINPUT101), .ZN(n729) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n745), .ZN(n734) );
  NOR2_X1 U809 ( .A1(n733), .A2(n734), .ZN(n725) );
  NAND2_X1 U810 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U811 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U812 ( .A1(n727), .A2(G168), .ZN(n728) );
  NOR2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U814 ( .A(n730), .B(KEYINPUT31), .ZN(n731) );
  NOR2_X1 U815 ( .A1(n733), .A2(n742), .ZN(n736) );
  NAND2_X1 U816 ( .A1(G8), .A2(n734), .ZN(n735) );
  NAND2_X1 U817 ( .A1(n736), .A2(n735), .ZN(n739) );
  INV_X1 U818 ( .A(n739), .ZN(n738) );
  INV_X1 U819 ( .A(KEYINPUT102), .ZN(n737) );
  NAND2_X1 U820 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U821 ( .A1(KEYINPUT102), .A2(n739), .ZN(n740) );
  NAND2_X1 U822 ( .A1(n741), .A2(n740), .ZN(n756) );
  INV_X1 U823 ( .A(n742), .ZN(n744) );
  AND2_X1 U824 ( .A1(G286), .A2(G8), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n744), .A2(n743), .ZN(n753) );
  INV_X1 U826 ( .A(G8), .ZN(n751) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n773), .ZN(n747) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U829 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U830 ( .A(KEYINPUT103), .B(n748), .Z(n749) );
  NAND2_X1 U831 ( .A1(n749), .A2(G303), .ZN(n750) );
  OR2_X1 U832 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U833 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U834 ( .A(n754), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U835 ( .A1(n756), .A2(n755), .ZN(n769) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U838 ( .A1(n760), .A2(n757), .ZN(n1017) );
  NAND2_X1 U839 ( .A1(n769), .A2(n1017), .ZN(n758) );
  XNOR2_X1 U840 ( .A(n758), .B(KEYINPUT104), .ZN(n766) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n1016) );
  INV_X1 U842 ( .A(n1016), .ZN(n759) );
  NOR2_X1 U843 ( .A1(n773), .A2(n759), .ZN(n763) );
  NAND2_X1 U844 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U845 ( .A1(n761), .A2(n773), .ZN(n775) );
  INV_X1 U846 ( .A(n775), .ZN(n762) );
  AND2_X1 U847 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U848 ( .A(G305), .B(G1981), .Z(n1031) );
  AND2_X1 U849 ( .A1(n764), .A2(n1031), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n783) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n770), .A2(n773), .ZN(n781) );
  NOR2_X1 U855 ( .A1(G305), .A2(G1981), .ZN(n771) );
  XOR2_X1 U856 ( .A(n771), .B(KEYINPUT24), .Z(n772) );
  OR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n779) );
  INV_X1 U858 ( .A(n1031), .ZN(n777) );
  INV_X1 U859 ( .A(KEYINPUT33), .ZN(n774) );
  OR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  AND2_X1 U863 ( .A1(n781), .A2(n780), .ZN(n782) );
  AND2_X1 U864 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U865 ( .A(n784), .B(KEYINPUT105), .ZN(n823) );
  XNOR2_X1 U866 ( .A(KEYINPUT94), .B(G1991), .ZN(n959) );
  NAND2_X1 U867 ( .A1(G107), .A2(n891), .ZN(n791) );
  NAND2_X1 U868 ( .A1(G95), .A2(n573), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G119), .A2(n890), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n894), .A2(G131), .ZN(n787) );
  XOR2_X1 U872 ( .A(KEYINPUT92), .B(n787), .Z(n788) );
  NOR2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U875 ( .A(n792), .B(KEYINPUT93), .Z(n900) );
  AND2_X1 U876 ( .A1(n959), .A2(n900), .ZN(n801) );
  NAND2_X1 U877 ( .A1(G141), .A2(n894), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G129), .A2(n890), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U880 ( .A1(n573), .A2(G105), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n891), .A2(G117), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n885) );
  AND2_X1 U885 ( .A1(n885), .A2(G1996), .ZN(n800) );
  NOR2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n985) );
  INV_X1 U887 ( .A(n802), .ZN(n803) );
  NOR2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n833) );
  XNOR2_X1 U889 ( .A(KEYINPUT95), .B(n833), .ZN(n805) );
  NOR2_X1 U890 ( .A1(n985), .A2(n805), .ZN(n827) );
  XNOR2_X1 U891 ( .A(KEYINPUT96), .B(n827), .ZN(n819) );
  XOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .Z(n806) );
  XNOR2_X1 U893 ( .A(KEYINPUT89), .B(n806), .ZN(n824) );
  NAND2_X1 U894 ( .A1(G140), .A2(n894), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G104), .A2(n573), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n809), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G128), .A2(n890), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G116), .A2(n891), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT90), .B(n812), .Z(n813) );
  XNOR2_X1 U902 ( .A(KEYINPUT35), .B(n813), .ZN(n814) );
  NOR2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n816), .ZN(n903) );
  NOR2_X1 U905 ( .A1(n824), .A2(n903), .ZN(n993) );
  NAND2_X1 U906 ( .A1(n993), .A2(n833), .ZN(n817) );
  XOR2_X1 U907 ( .A(KEYINPUT91), .B(n817), .Z(n830) );
  INV_X1 U908 ( .A(n830), .ZN(n818) );
  NOR2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n821) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n1015) );
  NAND2_X1 U911 ( .A1(n1015), .A2(n833), .ZN(n820) );
  AND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n836) );
  NAND2_X1 U914 ( .A1(n824), .A2(n903), .ZN(n997) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n885), .ZN(n989) );
  NOR2_X1 U916 ( .A1(n959), .A2(n900), .ZN(n983) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n983), .A2(n825), .ZN(n826) );
  NOR2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U920 ( .A1(n989), .A2(n828), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n997), .A2(n832), .ZN(n834) );
  NAND2_X1 U924 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U926 ( .A(n838), .B(n837), .ZN(G329) );
  NAND2_X1 U927 ( .A1(n839), .A2(G2106), .ZN(n840) );
  XNOR2_X1 U928 ( .A(n840), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U930 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U932 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n846), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n848) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2072), .Z(n850) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U946 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1976), .B(G1981), .Z(n856) );
  XNOR2_X1 U950 ( .A(G1971), .B(G1966), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U952 ( .A(n857), .B(KEYINPUT41), .Z(n859) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U955 ( .A(G2474), .B(G1956), .Z(n861) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1961), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n890), .ZN(n864) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(n864), .Z(n865) );
  XNOR2_X1 U961 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U962 ( .A1(G136), .A2(n894), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U964 ( .A1(G100), .A2(n573), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G112), .A2(n891), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(KEYINPUT110), .B(n872), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n874) );
  XNOR2_X1 U970 ( .A(KEYINPUT114), .B(KEYINPUT113), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U972 ( .A(n875), .B(KEYINPUT48), .Z(n877) );
  XNOR2_X1 U973 ( .A(G164), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n889) );
  XNOR2_X1 U975 ( .A(G162), .B(n982), .ZN(n887) );
  NAND2_X1 U976 ( .A1(G139), .A2(n894), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G103), .A2(n573), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G127), .A2(n890), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G115), .A2(n891), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n999) );
  XOR2_X1 U984 ( .A(n885), .B(n999), .Z(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n905) );
  NAND2_X1 U987 ( .A1(G130), .A2(n890), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U990 ( .A1(G142), .A2(n894), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G106), .A2(n573), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U993 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U998 ( .A(n906), .B(G160), .Z(n907) );
  NOR2_X1 U999 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n1024), .B(n1011), .Z(n908) );
  XOR2_X1 U1001 ( .A(n908), .B(KEYINPUT115), .Z(n911) );
  XNOR2_X1 U1002 ( .A(G171), .B(n909), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1004 ( .A(G286), .B(n912), .Z(n913) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n913), .ZN(G397) );
  XOR2_X1 U1006 ( .A(KEYINPUT107), .B(G2451), .Z(n915) );
  XNOR2_X1 U1007 ( .A(G2446), .B(G2427), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(n922) );
  XOR2_X1 U1009 ( .A(G2438), .B(G2435), .Z(n917) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2430), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1012 ( .A(n918), .B(G2454), .Z(n920) );
  XNOR2_X1 U1013 ( .A(G1341), .B(G1348), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n922), .B(n921), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(n923), .A2(G14), .ZN(n929) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n929), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n924), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G108), .ZN(G238) );
  INV_X1 U1025 ( .A(n929), .ZN(G401) );
  XOR2_X1 U1026 ( .A(G1976), .B(G23), .Z(n931) );
  XOR2_X1 U1027 ( .A(G1971), .B(G22), .Z(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G24), .B(G1986), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT58), .B(n934), .Z(n955) );
  XOR2_X1 U1032 ( .A(n935), .B(G5), .Z(n938) );
  XNOR2_X1 U1033 ( .A(G21), .B(KEYINPUT125), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n936), .B(G1966), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n952) );
  XNOR2_X1 U1036 ( .A(n939), .B(G20), .ZN(n948) );
  XOR2_X1 U1037 ( .A(G1341), .B(G19), .Z(n943) );
  XOR2_X1 U1038 ( .A(KEYINPUT59), .B(G4), .Z(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT123), .B(n940), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(G1348), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT122), .B(G1981), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G6), .B(n944), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n949), .B(KEYINPUT60), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(n950), .B(KEYINPUT124), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT126), .B(n953), .Z(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT61), .B(n956), .Z(n957) );
  NOR2_X1 U1052 ( .A1(G16), .A2(n957), .ZN(n981) );
  INV_X1 U1053 ( .A(KEYINPUT55), .ZN(n1006) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G35), .ZN(n972) );
  XOR2_X1 U1055 ( .A(G2072), .B(G33), .Z(n958) );
  NAND2_X1 U1056 ( .A1(n958), .A2(G28), .ZN(n969) );
  XOR2_X1 U1057 ( .A(KEYINPUT118), .B(n959), .Z(n960) );
  XNOR2_X1 U1058 ( .A(n960), .B(G25), .ZN(n967) );
  XOR2_X1 U1059 ( .A(G2067), .B(G26), .Z(n962) );
  XOR2_X1 U1060 ( .A(G1996), .B(G32), .Z(n961) );
  NAND2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(G27), .B(n963), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT53), .B(n970), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G2084), .B(KEYINPUT54), .Z(n973) );
  XNOR2_X1 U1069 ( .A(G34), .B(n973), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(n1006), .B(n976), .ZN(n978) );
  INV_X1 U1072 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n1010) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G2084), .B(G160), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n990), .B(KEYINPUT51), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(KEYINPUT116), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT117), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1004) );
  XOR2_X1 U1088 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1091 ( .A(KEYINPUT50), .B(n1002), .Z(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(G29), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1039) );
  XNOR2_X1 U1097 ( .A(G301), .B(G1961), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1011), .B(G1341), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1028) );
  XNOR2_X1 U1100 ( .A(G1956), .B(G299), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1023) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  INV_X1 U1103 ( .A(G1971), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(G166), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT121), .B(n1021), .Z(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(G1348), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(n1034) );
  XNOR2_X1 U1111 ( .A(G168), .B(G1966), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT120), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(KEYINPUT57), .B(n1032), .Z(n1033) );
  NOR2_X1 U1115 ( .A1(n1034), .A2(n1033), .ZN(n1037) );
  XNOR2_X1 U1116 ( .A(G16), .B(KEYINPUT119), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(KEYINPUT56), .B(n1035), .ZN(n1036) );
  NOR2_X1 U1118 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1119 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1120 ( .A(n1040), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

