//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AND2_X1   g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n471), .A2(new_n468), .A3(G101), .A4(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n467), .A2(G137), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n474), .B1(new_n465), .B2(new_n466), .ZN(new_n475));
  AND2_X1   g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  XNOR2_X1  g054(.A(new_n467), .B(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n468), .B1(new_n465), .B2(new_n466), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n468), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(G2104), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n468), .C1(new_n495), .C2(new_n496), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT3), .B(G2104), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G138), .A4(new_n468), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n500), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n518), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n515), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n512), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(G543), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT73), .B(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n529), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(G52), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n522), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n519), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n519), .A2(G53), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n512), .A2(new_n521), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n555), .B(new_n557), .C1(new_n514), .C2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G166), .ZN(G303));
  OAI21_X1  g136(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT75), .Z(new_n563));
  AOI22_X1  g138(.A1(new_n556), .A2(G87), .B1(G49), .B2(new_n519), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(G288));
  INV_X1    g140(.A(G61), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n510), .B2(new_n511), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  INV_X1    g143(.A(G73), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(new_n516), .ZN(new_n570));
  AND2_X1   g145(.A1(KEYINPUT5), .A2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT5), .A2(G543), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n568), .B(G61), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n522), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n514), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n519), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n522), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n556), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n526), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G321));
  MUX2_X1   g173(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g174(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g175(.A(KEYINPUT77), .B(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n596), .B1(G860), .B2(new_n601), .ZN(G148));
  NAND2_X1  g177(.A1(new_n596), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g181(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n607));
  NOR3_X1   g182(.A1(new_n463), .A2(new_n464), .A3(G2105), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G2100), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT79), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n480), .A2(G135), .ZN(new_n614));
  INV_X1    g189(.A(G111), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n615), .A2(KEYINPUT80), .A3(G2105), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT80), .B1(new_n615), .B2(G2105), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n616), .A2(new_n619), .B1(new_n485), .B2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G2096), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n611), .A2(G2100), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n613), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(G156));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT81), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n632), .B(new_n636), .Z(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(G14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT83), .B(KEYINPUT17), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n644), .B2(new_n647), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n652), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n660), .A2(new_n665), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(new_n665), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n668));
  AOI211_X1 g243(.A(new_n664), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT85), .Z(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n671), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G23), .ZN(new_n680));
  INV_X1    g255(.A(G288), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT87), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT33), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(G1976), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(G1976), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n679), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n569), .A2(new_n516), .ZN(new_n691));
  OAI21_X1  g266(.A(G61), .B1(new_n571), .B2(new_n572), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(KEYINPUT76), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n514), .B1(new_n693), .B2(new_n573), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(new_n578), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n690), .B1(new_n695), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n689), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n685), .A2(new_n686), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n703));
  NOR2_X1   g278(.A1(G16), .A2(G24), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n586), .B2(G16), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT88), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n480), .A2(G131), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n485), .A2(G119), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n468), .A2(G107), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G25), .B(new_n713), .S(G29), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n708), .B(new_n717), .C1(new_n707), .C2(new_n706), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n702), .A2(new_n703), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n679), .A2(G4), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n596), .B2(new_n679), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1348), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT95), .B(G2078), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G27), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G164), .B2(new_n726), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G168), .A2(new_n679), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n679), .B2(G21), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT91), .B(G1966), .Z(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n548), .B2(G16), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n731), .A2(new_n732), .B1(new_n734), .B2(G1341), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT31), .B(G11), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT93), .B(G28), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT94), .Z(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n621), .B2(new_n726), .ZN(new_n742));
  NOR2_X1   g317(.A1(G171), .A2(new_n679), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G5), .B2(new_n679), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n735), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  INV_X1    g323(.A(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n749), .B2(KEYINPUT24), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT24), .B2(new_n749), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n478), .B2(new_n726), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n734), .A2(G1341), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n748), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n744), .B2(new_n745), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n747), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G35), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G162), .B2(G29), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n726), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n480), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n485), .A2(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n468), .A2(G116), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(G2067), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n726), .A2(G33), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n504), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n468), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n480), .B2(G139), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n773), .B1(new_n778), .B2(new_n726), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2072), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n762), .A2(new_n772), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n729), .A2(new_n756), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n726), .A2(G32), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT26), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n784), .B(new_n786), .C1(G129), .C2(new_n485), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G141), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n726), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT90), .Z(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n793), .A2(new_n794), .B1(new_n761), .B2(new_n760), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n731), .A2(new_n732), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT92), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n679), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT97), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n798), .B(new_n803), .C1(new_n725), .C2(new_n728), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n782), .A2(new_n796), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n721), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n719), .A2(new_n720), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(G311));
  INV_X1    g383(.A(new_n807), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n809), .A2(new_n721), .A3(new_n805), .ZN(G150));
  NAND2_X1  g385(.A1(new_n596), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n514), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n519), .A2(G55), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n522), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n548), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n548), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n812), .B(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n824), .A2(new_n825), .A3(G860), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n814), .B2(new_n817), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT98), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  OR2_X1    g404(.A1(new_n826), .A2(new_n829), .ZN(G145));
  XNOR2_X1  g405(.A(new_n769), .B(new_n789), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n507), .A2(KEYINPUT99), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n503), .A2(new_n506), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n498), .A2(KEYINPUT100), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n494), .A2(new_n836), .A3(new_n497), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n832), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n831), .A2(new_n839), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n778), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n778), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n713), .B(new_n609), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n480), .A2(G142), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G118), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n849), .A2(new_n850), .B1(new_n852), .B2(G2105), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n851), .A2(new_n853), .B1(new_n485), .B2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n847), .B(new_n855), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n846), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n621), .B(new_n487), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n478), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n857), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g437(.A(G288), .B(new_n695), .ZN(new_n863));
  XOR2_X1   g438(.A(G166), .B(new_n586), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT103), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n595), .B(G299), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(KEYINPUT41), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n603), .B(new_n822), .ZN(new_n871));
  MUX2_X1   g446(.A(new_n869), .B(new_n870), .S(new_n871), .Z(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT104), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(KEYINPUT104), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n873), .A2(new_n867), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G868), .B2(new_n818), .ZN(G295));
  OAI21_X1  g453(.A(new_n877), .B1(G868), .B2(new_n818), .ZN(G331));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  OAI21_X1  g456(.A(G286), .B1(G171), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(G171), .A2(new_n881), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n882), .B(new_n883), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n821), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n882), .B(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n822), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n868), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n885), .A2(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n870), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n891), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n892), .A2(new_n865), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n870), .A2(new_n886), .A3(new_n889), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n868), .B2(new_n893), .ZN(new_n898));
  INV_X1    g473(.A(new_n865), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(KEYINPUT109), .A3(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n880), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n894), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n890), .A2(new_n891), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n896), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(new_n880), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT44), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(new_n913), .A3(KEYINPUT43), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n910), .B2(KEYINPUT43), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n912), .B1(new_n917), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n835), .A2(new_n834), .A3(new_n837), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n833), .B1(new_n503), .B2(new_n506), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n473), .A2(new_n477), .A3(G40), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n473), .A2(new_n477), .A3(KEYINPUT110), .A4(G40), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n930), .A2(KEYINPUT111), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(KEYINPUT111), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1996), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n790), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT112), .Z(new_n936));
  AND2_X1   g511(.A1(new_n713), .A2(new_n716), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n716), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G2067), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n769), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n934), .B2(new_n790), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n936), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n586), .A2(new_n707), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n933), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n927), .A3(new_n928), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT45), .B1(new_n838), .B2(new_n919), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n732), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n498), .A2(new_n499), .B1(new_n503), .B2(new_n506), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n955), .B2(new_n501), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n508), .A2(new_n919), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n838), .A2(new_n957), .A3(new_n919), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n927), .A2(new_n748), .A3(new_n928), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n953), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  NOR2_X1   g540(.A1(G168), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT121), .Z(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(G8), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n969), .B(new_n970), .C1(new_n965), .C2(G168), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT122), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n965), .B1(new_n953), .B2(new_n963), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n966), .B1(new_n974), .B2(KEYINPUT122), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n976), .B2(KEYINPUT123), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT123), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n978), .B(new_n970), .C1(new_n973), .C2(new_n975), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n968), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n960), .A2(new_n961), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n927), .A2(new_n928), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT114), .B(G2090), .Z(new_n983));
  NAND4_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n958), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n508), .B2(new_n919), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n929), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n838), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n987));
  AOI21_X1  g562(.A(G1971), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n965), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G166), .A2(new_n965), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n991), .A2(KEYINPUT55), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(KEYINPUT55), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT115), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n994), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n927), .B(new_n928), .C1(new_n959), .C2(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n957), .B1(new_n838), .B2(new_n919), .ZN(new_n1001));
  INV_X1    g576(.A(new_n983), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G8), .B1(new_n1003), .B2(new_n988), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n990), .A2(new_n998), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n838), .A2(new_n919), .A3(new_n927), .A4(new_n928), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n563), .A2(G1976), .A3(new_n564), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(G8), .A4(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1009), .B(G8), .C1(new_n922), .C2(new_n929), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n575), .B2(new_n579), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n694), .A2(G1981), .A3(new_n578), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT116), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1015), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1016), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT49), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(G8), .A3(new_n1008), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1010), .B(new_n1012), .C1(new_n1021), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n922), .A2(new_n929), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n965), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(new_n1024), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(KEYINPUT117), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1005), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n982), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT124), .B(G1961), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n959), .A2(new_n923), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n987), .A2(new_n1039), .A3(new_n982), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(G2078), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n924), .A2(new_n982), .A3(new_n950), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1038), .A2(G2078), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1037), .B(new_n1041), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G171), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT125), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT125), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1045), .A2(new_n1049), .A3(G171), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n925), .A2(new_n1044), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n924), .A2(new_n987), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1037), .A2(new_n1041), .A3(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1045), .A2(G301), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(KEYINPUT54), .C1(new_n1053), .C2(G301), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1034), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  XNOR2_X1  g634(.A(G299), .B(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n986), .A2(new_n987), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1060), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1068), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT61), .B1(new_n1070), .B2(new_n1065), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT58), .B(G1341), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n1040), .A2(G1996), .B1(new_n1029), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n548), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT59), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n1077));
  INV_X1    g652(.A(G1348), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1035), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1029), .A2(KEYINPUT119), .A3(new_n940), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1008), .B2(G2067), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1077), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1084), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n1079), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1087), .A3(new_n596), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n595), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1072), .A2(new_n1076), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n595), .B1(new_n1086), .B2(new_n1079), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1066), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1089), .A2(KEYINPUT120), .A3(new_n595), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1068), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n980), .A2(new_n1058), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n969), .A2(G286), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1005), .A2(new_n1033), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1005), .A2(new_n1033), .A3(KEYINPUT118), .A4(new_n1099), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1026), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(KEYINPUT63), .A3(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n990), .A2(new_n998), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n990), .B2(new_n994), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1031), .A2(new_n1006), .A3(new_n681), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1023), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1108), .A2(new_n1106), .B1(new_n1113), .B2(new_n1030), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1098), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1117), .B(new_n968), .C1(new_n977), .C2(new_n979), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1034), .B1(new_n1050), .B2(new_n1047), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n949), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n936), .A2(new_n938), .A3(new_n943), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n769), .A2(G2067), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n933), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n933), .A2(new_n934), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT46), .ZN(new_n1128));
  INV_X1    g703(.A(new_n941), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n933), .B1(new_n789), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT47), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n933), .A2(new_n946), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT48), .Z(new_n1134));
  OR2_X1    g709(.A1(new_n944), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1126), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT126), .B1(new_n1121), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1098), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n945), .B(new_n948), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1131), .A2(KEYINPUT47), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1131), .A2(KEYINPUT47), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1142), .A2(new_n1143), .B1(new_n944), .B2(new_n1134), .ZN(new_n1144));
  INV_X1    g719(.A(new_n933), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1140), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1137), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g724(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1151));
  XNOR2_X1  g725(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g726(.A1(new_n861), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n917), .A2(new_n1153), .ZN(G308));
  OR2_X1    g728(.A1(new_n915), .A2(new_n916), .ZN(new_n1155));
  OAI211_X1 g729(.A(new_n861), .B(new_n1152), .C1(new_n1155), .C2(new_n914), .ZN(G225));
endmodule


