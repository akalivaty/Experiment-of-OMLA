

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733;

  XNOR2_X1 U367 ( .A(n659), .B(n346), .ZN(G75) );
  XNOR2_X1 U368 ( .A(n660), .B(KEYINPUT53), .ZN(n346) );
  XNOR2_X1 U369 ( .A(n539), .B(KEYINPUT1), .ZN(n580) );
  XNOR2_X1 U370 ( .A(n449), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X2 U371 ( .A(n501), .B(n500), .ZN(n696) );
  XNOR2_X2 U372 ( .A(n477), .B(n476), .ZN(n724) );
  XNOR2_X1 U373 ( .A(n412), .B(KEYINPUT10), .ZN(n723) );
  INV_X1 U374 ( .A(G953), .ZN(n726) );
  XNOR2_X2 U375 ( .A(n545), .B(KEYINPUT40), .ZN(n372) );
  XNOR2_X2 U376 ( .A(n521), .B(n520), .ZN(n687) );
  NOR2_X2 U377 ( .A1(n609), .A2(n509), .ZN(n510) );
  XNOR2_X2 U378 ( .A(n381), .B(n508), .ZN(n609) );
  XNOR2_X2 U379 ( .A(n495), .B(n494), .ZN(n550) );
  NAND2_X1 U380 ( .A1(n594), .A2(n593), .ZN(n600) );
  AND2_X1 U381 ( .A1(n397), .A2(n398), .ZN(n383) );
  NAND2_X1 U382 ( .A1(n359), .A2(n562), .ZN(n611) );
  OR2_X1 U383 ( .A1(n586), .A2(n544), .ZN(n545) );
  OR2_X1 U384 ( .A1(n530), .A2(n371), .ZN(n370) );
  XNOR2_X1 U385 ( .A(n556), .B(KEYINPUT42), .ZN(n608) );
  XNOR2_X1 U386 ( .A(n564), .B(KEYINPUT79), .ZN(n682) );
  XNOR2_X1 U387 ( .A(n559), .B(KEYINPUT111), .ZN(n560) );
  NAND2_X2 U388 ( .A1(n390), .A2(n387), .ZN(n625) );
  XNOR2_X1 U389 ( .A(n402), .B(n401), .ZN(n704) );
  XNOR2_X1 U390 ( .A(n348), .B(n489), .ZN(n401) );
  XNOR2_X1 U391 ( .A(n438), .B(G113), .ZN(n483) );
  XNOR2_X2 U392 ( .A(KEYINPUT3), .B(G116), .ZN(n438) );
  XNOR2_X1 U393 ( .A(G125), .B(G146), .ZN(n443) );
  AND2_X2 U394 ( .A1(n600), .A2(n621), .ZN(n347) );
  XNOR2_X1 U395 ( .A(n403), .B(n723), .ZN(n402) );
  XNOR2_X2 U396 ( .A(n724), .B(G146), .ZN(n501) );
  XNOR2_X1 U397 ( .A(KEYINPUT68), .B(G131), .ZN(n475) );
  OR2_X1 U398 ( .A1(n550), .A2(n623), .ZN(n627) );
  XNOR2_X1 U399 ( .A(G101), .B(KEYINPUT89), .ZN(n441) );
  XOR2_X1 U400 ( .A(G104), .B(G107), .Z(n442) );
  XNOR2_X1 U401 ( .A(n611), .B(KEYINPUT86), .ZN(n574) );
  INV_X1 U402 ( .A(KEYINPUT46), .ZN(n379) );
  NAND2_X1 U403 ( .A1(n696), .A2(G469), .ZN(n355) );
  XNOR2_X1 U404 ( .A(G134), .B(G107), .ZN(n427) );
  XNOR2_X1 U405 ( .A(G113), .B(G143), .ZN(n417) );
  INV_X1 U406 ( .A(G137), .ZN(n473) );
  INV_X1 U407 ( .A(KEYINPUT84), .ZN(n595) );
  INV_X1 U408 ( .A(n638), .ZN(n377) );
  NAND2_X2 U409 ( .A1(n356), .A2(n357), .ZN(n539) );
  OR2_X1 U410 ( .A1(n696), .A2(n361), .ZN(n357) );
  AND2_X1 U411 ( .A1(n355), .A2(n350), .ZN(n356) );
  NAND2_X1 U412 ( .A1(n693), .A2(n362), .ZN(n361) );
  NAND2_X1 U413 ( .A1(n389), .A2(n362), .ZN(n388) );
  INV_X1 U414 ( .A(G140), .ZN(n411) );
  XNOR2_X1 U415 ( .A(n367), .B(n451), .ZN(n613) );
  XNOR2_X1 U416 ( .A(n717), .B(n499), .ZN(n367) );
  XNOR2_X1 U417 ( .A(n448), .B(n447), .ZN(n450) );
  BUF_X1 U418 ( .A(n580), .Z(n363) );
  XNOR2_X1 U419 ( .A(n373), .B(n543), .ZN(n586) );
  XNOR2_X1 U420 ( .A(n456), .B(n457), .ZN(n369) );
  INV_X1 U421 ( .A(KEYINPUT6), .ZN(n393) );
  XNOR2_X1 U422 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U423 ( .A(n472), .B(n471), .ZN(n530) );
  XNOR2_X1 U424 ( .A(n470), .B(KEYINPUT64), .ZN(n471) );
  AND2_X1 U425 ( .A1(n682), .A2(n565), .ZN(n566) );
  NAND2_X1 U426 ( .A1(n639), .A2(n638), .ZN(n378) );
  XNOR2_X1 U427 ( .A(G119), .B(G101), .ZN(n479) );
  XNOR2_X1 U428 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U429 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n446) );
  NAND2_X1 U430 ( .A1(G237), .A2(G234), .ZN(n458) );
  XNOR2_X1 U431 ( .A(n368), .B(n440), .ZN(n717) );
  XNOR2_X1 U432 ( .A(n483), .B(KEYINPUT16), .ZN(n368) );
  XOR2_X1 U433 ( .A(KEYINPUT74), .B(G122), .Z(n439) );
  XNOR2_X1 U434 ( .A(G119), .B(G110), .ZN(n490) );
  XNOR2_X1 U435 ( .A(n404), .B(G137), .ZN(n403) );
  XNOR2_X1 U436 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U437 ( .A(n395), .B(n394), .ZN(n487) );
  INV_X1 U438 ( .A(KEYINPUT8), .ZN(n394) );
  NAND2_X1 U439 ( .A1(n726), .A2(G234), .ZN(n395) );
  XNOR2_X1 U440 ( .A(G116), .B(G122), .ZN(n426) );
  XOR2_X1 U441 ( .A(G104), .B(G122), .Z(n419) );
  INV_X1 U442 ( .A(KEYINPUT77), .ZN(n598) );
  NAND2_X1 U443 ( .A1(n709), .A2(n597), .ZN(n599) );
  NOR2_X1 U444 ( .A1(n641), .A2(n377), .ZN(n376) );
  AND2_X1 U445 ( .A1(n374), .A2(n352), .ZN(n571) );
  INV_X1 U446 ( .A(n627), .ZN(n522) );
  NAND2_X1 U447 ( .A1(n369), .A2(n465), .ZN(n468) );
  AND2_X1 U448 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U449 ( .A1(n486), .A2(G902), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n601), .B(KEYINPUT62), .ZN(n602) );
  INV_X1 U451 ( .A(n728), .ZN(n375) );
  XNOR2_X1 U452 ( .A(G140), .B(G110), .ZN(n497) );
  XNOR2_X1 U453 ( .A(n613), .B(n612), .ZN(n614) );
  AND2_X1 U454 ( .A1(n604), .A2(G953), .ZN(n706) );
  XNOR2_X1 U455 ( .A(n360), .B(n561), .ZN(n359) );
  NAND2_X1 U456 ( .A1(n560), .A2(n385), .ZN(n360) );
  NAND2_X1 U457 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U458 ( .A1(n396), .A2(n400), .ZN(n382) );
  NAND2_X1 U459 ( .A1(n351), .A2(n562), .ZN(n371) );
  XNOR2_X1 U460 ( .A(n519), .B(KEYINPUT31), .ZN(n520) );
  AND2_X1 U461 ( .A1(n513), .A2(n512), .ZN(n684) );
  XNOR2_X1 U462 ( .A(G128), .B(n490), .ZN(n348) );
  XOR2_X1 U463 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n349) );
  NAND2_X1 U464 ( .A1(G469), .A2(G902), .ZN(n350) );
  AND2_X1 U465 ( .A1(n365), .A2(n550), .ZN(n351) );
  AND2_X1 U466 ( .A1(n539), .A2(n540), .ZN(n352) );
  INV_X1 U467 ( .A(n557), .ZN(n365) );
  XNOR2_X1 U468 ( .A(n625), .B(n393), .ZN(n557) );
  AND2_X1 U469 ( .A1(n587), .A2(KEYINPUT2), .ZN(n353) );
  XOR2_X1 U470 ( .A(KEYINPUT112), .B(KEYINPUT30), .Z(n354) );
  INV_X1 U471 ( .A(G902), .ZN(n362) );
  NAND2_X1 U472 ( .A1(n588), .A2(n587), .ZN(n358) );
  NAND2_X1 U473 ( .A1(n588), .A2(n353), .ZN(n596) );
  XNOR2_X1 U474 ( .A(n358), .B(KEYINPUT83), .ZN(n589) );
  XNOR2_X1 U475 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U476 ( .A1(n580), .A2(n522), .ZN(n366) );
  AND2_X1 U477 ( .A1(n406), .A2(n568), .ZN(n385) );
  NAND2_X1 U478 ( .A1(n364), .A2(n557), .ZN(n506) );
  XNOR2_X1 U479 ( .A(n516), .B(KEYINPUT110), .ZN(n364) );
  XNOR2_X2 U480 ( .A(n366), .B(KEYINPUT75), .ZN(n516) );
  NAND2_X1 U481 ( .A1(n563), .A2(n369), .ZN(n564) );
  XNOR2_X2 U482 ( .A(n370), .B(KEYINPUT32), .ZN(n733) );
  NAND2_X1 U483 ( .A1(n372), .A2(n608), .ZN(n380) );
  XNOR2_X1 U484 ( .A(n372), .B(G131), .ZN(G33) );
  NAND2_X1 U485 ( .A1(n571), .A2(n639), .ZN(n373) );
  XNOR2_X1 U486 ( .A(n541), .B(n354), .ZN(n374) );
  XNOR2_X1 U487 ( .A(n589), .B(n375), .ZN(n727) );
  NAND2_X1 U488 ( .A1(n639), .A2(n376), .ZN(n547) );
  NOR2_X1 U489 ( .A1(n637), .A2(n378), .ZN(n643) );
  XNOR2_X1 U490 ( .A(n380), .B(n379), .ZN(n575) );
  INV_X1 U491 ( .A(n539), .ZN(n524) );
  XNOR2_X2 U492 ( .A(n384), .B(G143), .ZN(n449) );
  XNOR2_X2 U493 ( .A(G128), .B(KEYINPUT80), .ZN(n384) );
  NAND2_X1 U494 ( .A1(n560), .A2(n406), .ZN(n581) );
  INV_X1 U495 ( .A(n568), .ZN(n386) );
  OR2_X1 U496 ( .A1(n601), .A2(n388), .ZN(n387) );
  INV_X1 U497 ( .A(n486), .ZN(n389) );
  NAND2_X1 U498 ( .A1(n601), .A2(n486), .ZN(n392) );
  INV_X1 U499 ( .A(n625), .ZN(n514) );
  INV_X1 U500 ( .A(n636), .ZN(n396) );
  XNOR2_X2 U501 ( .A(n506), .B(n505), .ZN(n636) );
  NAND2_X1 U502 ( .A1(n636), .A2(n507), .ZN(n397) );
  AND2_X1 U503 ( .A1(n399), .A2(n567), .ZN(n398) );
  NAND2_X1 U504 ( .A1(n515), .A2(n507), .ZN(n399) );
  NOR2_X1 U505 ( .A1(n515), .A2(n507), .ZN(n400) );
  AND2_X2 U506 ( .A1(n709), .A2(n589), .ZN(n619) );
  XOR2_X1 U507 ( .A(n349), .B(n488), .Z(n404) );
  AND2_X1 U508 ( .A1(G214), .A2(n478), .ZN(n405) );
  AND2_X1 U509 ( .A1(n684), .A2(n638), .ZN(n406) );
  AND2_X1 U510 ( .A1(n573), .A2(n574), .ZN(n407) );
  XOR2_X1 U511 ( .A(KEYINPUT109), .B(n532), .Z(n408) );
  BUF_X1 U512 ( .A(n636), .Z(n651) );
  XNOR2_X1 U513 ( .A(n443), .B(n411), .ZN(n412) );
  XNOR2_X1 U514 ( .A(n415), .B(n405), .ZN(n416) );
  XNOR2_X1 U515 ( .A(n439), .B(n490), .ZN(n440) );
  XNOR2_X1 U516 ( .A(n723), .B(n416), .ZN(n422) );
  XNOR2_X1 U517 ( .A(n423), .B(n662), .ZN(n424) );
  XNOR2_X1 U518 ( .A(n425), .B(n424), .ZN(n511) );
  XNOR2_X1 U519 ( .A(KEYINPUT15), .B(G902), .ZN(n591) );
  NAND2_X1 U520 ( .A1(G234), .A2(n591), .ZN(n409) );
  XNOR2_X1 U521 ( .A(KEYINPUT20), .B(n409), .ZN(n491) );
  NAND2_X1 U522 ( .A1(n491), .A2(G221), .ZN(n410) );
  XNOR2_X1 U523 ( .A(n410), .B(KEYINPUT21), .ZN(n623) );
  XOR2_X1 U524 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n414) );
  XNOR2_X1 U525 ( .A(KEYINPUT103), .B(KEYINPUT11), .ZN(n413) );
  XNOR2_X1 U526 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U527 ( .A1(G953), .A2(G237), .ZN(n478) );
  XOR2_X1 U528 ( .A(n417), .B(KEYINPUT102), .Z(n418) );
  XNOR2_X1 U529 ( .A(n475), .B(n418), .ZN(n420) );
  XNOR2_X1 U530 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U531 ( .A(n422), .B(n421), .ZN(n663) );
  NOR2_X1 U532 ( .A1(G902), .A2(n663), .ZN(n425) );
  XNOR2_X1 U533 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n423) );
  INV_X1 U534 ( .A(G475), .ZN(n662) );
  XNOR2_X1 U535 ( .A(n426), .B(KEYINPUT7), .ZN(n430) );
  XOR2_X1 U536 ( .A(KEYINPUT9), .B(KEYINPUT106), .Z(n428) );
  XNOR2_X1 U537 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U538 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U539 ( .A1(G217), .A2(n487), .ZN(n431) );
  XNOR2_X1 U540 ( .A(n432), .B(n431), .ZN(n434) );
  INV_X1 U541 ( .A(n449), .ZN(n433) );
  XNOR2_X1 U542 ( .A(n434), .B(n433), .ZN(n700) );
  NAND2_X1 U543 ( .A1(n700), .A2(n362), .ZN(n436) );
  XNOR2_X1 U544 ( .A(KEYINPUT107), .B(G478), .ZN(n435) );
  XNOR2_X1 U545 ( .A(n436), .B(n435), .ZN(n512) );
  NAND2_X1 U546 ( .A1(n511), .A2(n512), .ZN(n641) );
  NOR2_X1 U547 ( .A1(n623), .A2(n641), .ZN(n437) );
  XNOR2_X1 U548 ( .A(KEYINPUT108), .B(n437), .ZN(n469) );
  XOR2_X1 U549 ( .A(KEYINPUT19), .B(KEYINPUT65), .Z(n457) );
  XNOR2_X1 U550 ( .A(n442), .B(n441), .ZN(n716) );
  XNOR2_X1 U551 ( .A(n716), .B(KEYINPUT70), .ZN(n499) );
  INV_X1 U552 ( .A(n443), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n444), .B(KEYINPUT18), .ZN(n448) );
  NAND2_X1 U554 ( .A1(G224), .A2(n726), .ZN(n445) );
  XNOR2_X1 U555 ( .A(n477), .B(n450), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n613), .A2(n591), .ZN(n454) );
  OR2_X1 U557 ( .A1(G902), .A2(G237), .ZN(n452) );
  XNOR2_X1 U558 ( .A(KEYINPUT76), .B(n452), .ZN(n455) );
  AND2_X1 U559 ( .A1(n455), .A2(G210), .ZN(n453) );
  XNOR2_X2 U560 ( .A(n454), .B(n453), .ZN(n568) );
  NAND2_X1 U561 ( .A1(n455), .A2(G214), .ZN(n638) );
  NAND2_X1 U562 ( .A1(n568), .A2(n638), .ZN(n456) );
  XNOR2_X1 U563 ( .A(n458), .B(KEYINPUT14), .ZN(n461) );
  NAND2_X1 U564 ( .A1(G952), .A2(n461), .ZN(n649) );
  NOR2_X1 U565 ( .A1(G953), .A2(n649), .ZN(n459) );
  XOR2_X1 U566 ( .A(KEYINPUT91), .B(n459), .Z(n537) );
  NOR2_X1 U567 ( .A1(G898), .A2(n726), .ZN(n460) );
  XOR2_X1 U568 ( .A(KEYINPUT92), .B(n460), .Z(n719) );
  NAND2_X1 U569 ( .A1(n461), .A2(G902), .ZN(n462) );
  XOR2_X1 U570 ( .A(KEYINPUT93), .B(n462), .Z(n535) );
  NOR2_X1 U571 ( .A1(n719), .A2(n535), .ZN(n463) );
  NOR2_X1 U572 ( .A1(n537), .A2(n463), .ZN(n464) );
  XOR2_X1 U573 ( .A(KEYINPUT94), .B(n464), .Z(n465) );
  INV_X1 U574 ( .A(KEYINPUT66), .ZN(n466) );
  XNOR2_X1 U575 ( .A(n466), .B(KEYINPUT0), .ZN(n467) );
  XNOR2_X2 U576 ( .A(n468), .B(n467), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n469), .A2(n523), .ZN(n472) );
  XOR2_X1 U578 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n470) );
  XNOR2_X1 U579 ( .A(n473), .B(G134), .ZN(n474) );
  XNOR2_X1 U580 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U581 ( .A1(n478), .A2(G210), .ZN(n480) );
  XNOR2_X1 U582 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U583 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U586 ( .A(n501), .B(n485), .ZN(n601) );
  XNOR2_X1 U587 ( .A(KEYINPUT98), .B(G472), .ZN(n486) );
  NAND2_X1 U588 ( .A1(G221), .A2(n487), .ZN(n489) );
  NOR2_X1 U589 ( .A1(n704), .A2(G902), .ZN(n495) );
  NAND2_X1 U590 ( .A1(n491), .A2(G217), .ZN(n493) );
  INV_X1 U591 ( .A(KEYINPUT25), .ZN(n492) );
  NAND2_X1 U592 ( .A1(n726), .A2(G227), .ZN(n496) );
  XNOR2_X1 U593 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U594 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U595 ( .A(G469), .ZN(n693) );
  XNOR2_X1 U596 ( .A(n363), .B(KEYINPUT88), .ZN(n562) );
  INV_X1 U597 ( .A(n363), .ZN(n628) );
  AND2_X1 U598 ( .A1(n550), .A2(n514), .ZN(n502) );
  NAND2_X1 U599 ( .A1(n628), .A2(n502), .ZN(n503) );
  NOR2_X1 U600 ( .A1(n530), .A2(n503), .ZN(n676) );
  INV_X1 U601 ( .A(n676), .ZN(n504) );
  NAND2_X1 U602 ( .A1(n733), .A2(n504), .ZN(n509) );
  XNOR2_X1 U603 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n505) );
  INV_X1 U604 ( .A(n523), .ZN(n515) );
  XNOR2_X1 U605 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n507) );
  NOR2_X1 U606 ( .A1(n511), .A2(n512), .ZN(n567) );
  XNOR2_X1 U607 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n510), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U609 ( .A(n511), .B(KEYINPUT105), .ZN(n513) );
  OR2_X1 U610 ( .A1(n513), .A2(n512), .ZN(n585) );
  INV_X1 U611 ( .A(n585), .ZN(n686) );
  NOR2_X1 U612 ( .A1(n684), .A2(n686), .ZN(n637) );
  NOR2_X1 U613 ( .A1(n515), .A2(n514), .ZN(n518) );
  BUF_X1 U614 ( .A(n516), .Z(n517) );
  NAND2_X1 U615 ( .A1(n518), .A2(n517), .ZN(n521) );
  XOR2_X1 U616 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n519) );
  NAND2_X1 U617 ( .A1(n523), .A2(n522), .ZN(n526) );
  OR2_X1 U618 ( .A1(n625), .A2(n524), .ZN(n525) );
  NOR2_X1 U619 ( .A1(n526), .A2(n525), .ZN(n671) );
  NOR2_X1 U620 ( .A1(n687), .A2(n671), .ZN(n527) );
  NOR2_X1 U621 ( .A1(n637), .A2(n527), .ZN(n531) );
  NOR2_X1 U622 ( .A1(n557), .A2(n550), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n528), .A2(n628), .ZN(n529) );
  NOR2_X1 U624 ( .A1(n530), .A2(n529), .ZN(n669) );
  NOR2_X1 U625 ( .A1(n531), .A2(n669), .ZN(n532) );
  NAND2_X1 U626 ( .A1(n533), .A2(n408), .ZN(n534) );
  XNOR2_X2 U627 ( .A(n534), .B(KEYINPUT45), .ZN(n709) );
  OR2_X1 U628 ( .A1(n726), .A2(n535), .ZN(n536) );
  NOR2_X1 U629 ( .A1(G900), .A2(n536), .ZN(n538) );
  NOR2_X1 U630 ( .A1(n538), .A2(n537), .ZN(n548) );
  NOR2_X1 U631 ( .A1(n627), .A2(n548), .ZN(n540) );
  NAND2_X1 U632 ( .A1(n625), .A2(n638), .ZN(n541) );
  INV_X1 U633 ( .A(KEYINPUT38), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n568), .B(n542), .ZN(n639) );
  INV_X1 U635 ( .A(KEYINPUT39), .ZN(n543) );
  INV_X1 U636 ( .A(n684), .ZN(n544) );
  INV_X1 U637 ( .A(KEYINPUT41), .ZN(n546) );
  XNOR2_X1 U638 ( .A(n547), .B(n546), .ZN(n650) );
  NOR2_X1 U639 ( .A1(n548), .A2(n623), .ZN(n549) );
  AND2_X1 U640 ( .A1(n550), .A2(n549), .ZN(n558) );
  NAND2_X1 U641 ( .A1(n558), .A2(n625), .ZN(n552) );
  INV_X1 U642 ( .A(KEYINPUT28), .ZN(n551) );
  XNOR2_X1 U643 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U644 ( .A(n524), .B(KEYINPUT113), .ZN(n553) );
  AND2_X1 U645 ( .A1(n554), .A2(n553), .ZN(n563) );
  INV_X1 U646 ( .A(n563), .ZN(n555) );
  OR2_X1 U647 ( .A1(n650), .A2(n555), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U649 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n561) );
  NOR2_X1 U650 ( .A1(n637), .A2(KEYINPUT67), .ZN(n565) );
  XNOR2_X1 U651 ( .A(n566), .B(KEYINPUT47), .ZN(n572) );
  INV_X1 U652 ( .A(n567), .ZN(n569) );
  NOR2_X1 U653 ( .A1(n569), .A2(n386), .ZN(n570) );
  NAND2_X1 U654 ( .A1(n571), .A2(n570), .ZN(n680) );
  AND2_X1 U655 ( .A1(n572), .A2(n680), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n575), .A2(n407), .ZN(n579) );
  XNOR2_X1 U657 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n577) );
  INV_X1 U658 ( .A(KEYINPUT69), .ZN(n576) );
  XNOR2_X1 U659 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U660 ( .A(n579), .B(n578), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n581), .A2(n363), .ZN(n583) );
  INV_X1 U662 ( .A(KEYINPUT43), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n584), .A2(n386), .ZN(n691) );
  OR2_X1 U665 ( .A1(n586), .A2(n585), .ZN(n689) );
  AND2_X1 U666 ( .A1(n691), .A2(n689), .ZN(n587) );
  INV_X1 U667 ( .A(n591), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n619), .A2(n590), .ZN(n594) );
  XOR2_X1 U669 ( .A(KEYINPUT82), .B(n591), .Z(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(KEYINPUT2), .ZN(n593) );
  XNOR2_X2 U671 ( .A(n599), .B(n598), .ZN(n621) );
  NAND2_X1 U672 ( .A1(n600), .A2(n621), .ZN(n692) );
  NAND2_X1 U673 ( .A1(n347), .A2(G472), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(n602), .ZN(n605) );
  INV_X1 U675 ( .A(G952), .ZN(n604) );
  NOR2_X2 U676 ( .A1(n605), .A2(n706), .ZN(n607) );
  INV_X1 U677 ( .A(KEYINPUT63), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n607), .B(n606), .ZN(G57) );
  XNOR2_X1 U679 ( .A(n608), .B(G137), .ZN(G39) );
  XOR2_X1 U680 ( .A(n609), .B(G122), .Z(G24) );
  XOR2_X1 U681 ( .A(G125), .B(KEYINPUT37), .Z(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(G27) );
  NAND2_X1 U683 ( .A1(n347), .A2(G210), .ZN(n615) );
  XNOR2_X1 U684 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X2 U686 ( .A1(n616), .A2(n706), .ZN(n618) );
  XNOR2_X1 U687 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(G51) );
  NOR2_X1 U689 ( .A1(n619), .A2(KEYINPUT2), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT81), .ZN(n622) );
  AND2_X1 U691 ( .A1(n621), .A2(n622), .ZN(n658) );
  NAND2_X1 U692 ( .A1(n517), .A2(n625), .ZN(n633) );
  NAND2_X1 U693 ( .A1(n550), .A2(n623), .ZN(n624) );
  XNOR2_X1 U694 ( .A(KEYINPUT49), .B(n624), .ZN(n626) );
  NOR2_X1 U695 ( .A1(n626), .A2(n625), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(KEYINPUT50), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U699 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n634), .B(KEYINPUT51), .ZN(n635) );
  NOR2_X1 U701 ( .A1(n635), .A2(n650), .ZN(n646) );
  NOR2_X1 U702 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U703 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U704 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U705 ( .A1(n651), .A2(n644), .ZN(n645) );
  NOR2_X1 U706 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U707 ( .A(n647), .B(KEYINPUT52), .ZN(n648) );
  NOR2_X1 U708 ( .A1(n649), .A2(n648), .ZN(n655) );
  OR2_X1 U709 ( .A1(n651), .A2(n650), .ZN(n653) );
  INV_X1 U710 ( .A(KEYINPUT118), .ZN(n652) );
  XNOR2_X1 U711 ( .A(n653), .B(n652), .ZN(n654) );
  OR2_X1 U712 ( .A1(n655), .A2(n654), .ZN(n656) );
  OR2_X1 U713 ( .A1(G953), .A2(n656), .ZN(n657) );
  NOR2_X1 U714 ( .A1(n658), .A2(n657), .ZN(n659) );
  INV_X1 U715 ( .A(KEYINPUT119), .ZN(n660) );
  NOR2_X1 U716 ( .A1(n692), .A2(n662), .ZN(n665) );
  XNOR2_X1 U717 ( .A(n663), .B(KEYINPUT59), .ZN(n664) );
  XNOR2_X1 U718 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U719 ( .A1(n666), .A2(n706), .ZN(n668) );
  XNOR2_X1 U720 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n667) );
  XNOR2_X1 U721 ( .A(n668), .B(n667), .ZN(G60) );
  XOR2_X1 U722 ( .A(G101), .B(n669), .Z(G3) );
  NAND2_X1 U723 ( .A1(n671), .A2(n684), .ZN(n670) );
  XNOR2_X1 U724 ( .A(n670), .B(G104), .ZN(G6) );
  XNOR2_X1 U725 ( .A(G107), .B(KEYINPUT27), .ZN(n675) );
  XOR2_X1 U726 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n673) );
  NAND2_X1 U727 ( .A1(n671), .A2(n686), .ZN(n672) );
  XNOR2_X1 U728 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U729 ( .A(n675), .B(n674), .ZN(G9) );
  XNOR2_X1 U730 ( .A(G110), .B(n676), .ZN(n677) );
  XNOR2_X1 U731 ( .A(n677), .B(KEYINPUT115), .ZN(G12) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n679) );
  NAND2_X1 U733 ( .A1(n682), .A2(n686), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n679), .B(n678), .ZN(G30) );
  XNOR2_X1 U735 ( .A(n680), .B(G143), .ZN(n681) );
  XNOR2_X1 U736 ( .A(KEYINPUT116), .B(n681), .ZN(G45) );
  NAND2_X1 U737 ( .A1(n682), .A2(n684), .ZN(n683) );
  XNOR2_X1 U738 ( .A(n683), .B(G146), .ZN(G48) );
  NAND2_X1 U739 ( .A1(n687), .A2(n684), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n685), .B(G113), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n688), .B(G116), .ZN(G18) );
  XOR2_X1 U743 ( .A(G134), .B(n689), .Z(n690) );
  XNOR2_X1 U744 ( .A(n690), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U745 ( .A(G140), .B(n691), .ZN(G42) );
  NOR2_X1 U746 ( .A1(n692), .A2(n693), .ZN(n698) );
  XNOR2_X1 U747 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n694) );
  XOR2_X1 U748 ( .A(n694), .B(KEYINPUT57), .Z(n695) );
  XNOR2_X1 U749 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U751 ( .A1(n706), .A2(n699), .ZN(G54) );
  NAND2_X1 U752 ( .A1(n347), .A2(G478), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n700), .B(KEYINPUT123), .ZN(n701) );
  XNOR2_X1 U754 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U755 ( .A1(n706), .A2(n703), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n347), .A2(G217), .ZN(n705) );
  XNOR2_X1 U757 ( .A(n705), .B(n704), .ZN(n707) );
  NOR2_X2 U758 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n708), .B(KEYINPUT124), .ZN(G66) );
  BUF_X1 U760 ( .A(n709), .Z(n710) );
  NAND2_X1 U761 ( .A1(n710), .A2(n726), .ZN(n715) );
  XOR2_X1 U762 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n712) );
  NAND2_X1 U763 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n713), .A2(G898), .ZN(n714) );
  NAND2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n722) );
  XNOR2_X1 U767 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(KEYINPUT126), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U770 ( .A(n722), .B(n721), .Z(G69) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT127), .ZN(n725) );
  XNOR2_X1 U772 ( .A(n724), .B(n725), .ZN(n728) );
  NAND2_X1 U773 ( .A1(n727), .A2(n726), .ZN(n732) );
  XNOR2_X1 U774 ( .A(G227), .B(n728), .ZN(n729) );
  NAND2_X1 U775 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U776 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U777 ( .A1(n732), .A2(n731), .ZN(G72) );
  XNOR2_X1 U778 ( .A(n733), .B(G119), .ZN(G21) );
endmodule

