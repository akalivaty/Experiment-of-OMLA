//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  AND2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n211), .B1(new_n212), .B2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n214), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n208), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n203), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n218), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n205), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n231), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n207), .A2(new_n232), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n232), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n257), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n214), .A2(new_n232), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n257), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n205), .B1(new_n268), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(new_n269), .B1(new_n205), .B2(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT9), .Z(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n286), .B1(new_n208), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n279), .B(new_n283), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n291), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT10), .B1(new_n272), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n272), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n291), .A2(new_n293), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT67), .Z(new_n300));
  OAI21_X1  g0100(.A(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n271), .B1(new_n291), .B2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n278), .B1(new_n281), .B2(new_n220), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n284), .A2(G226), .A3(new_n285), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n309), .B(new_n310), .C1(new_n287), .C2(new_n238), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n308), .B1(new_n311), .B2(new_n290), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(KEYINPUT13), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n314), .A2(new_n303), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(KEYINPUT69), .A3(KEYINPUT13), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT69), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n312), .B2(new_n315), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n312), .A2(KEYINPUT68), .A3(new_n315), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT68), .B1(new_n312), .B2(new_n315), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n319), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .A3(G169), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT14), .B1(new_n324), .B2(G169), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n318), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n266), .A2(new_n202), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n268), .A2(G20), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n267), .A2(G68), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n263), .A2(new_n205), .B1(new_n232), .B2(G68), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n260), .A2(new_n208), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n257), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g0138(.A(new_n338), .B(KEYINPUT11), .Z(new_n339));
  NOR3_X1   g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n328), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n314), .A2(new_n344), .A3(new_n316), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n324), .A2(G200), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n257), .ZN(new_n349));
  INV_X1    g0149(.A(new_n259), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT15), .B(G87), .Z(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n232), .A3(G33), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n267), .A2(G77), .A3(new_n331), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n214), .A2(G1), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G20), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(G77), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n287), .A2(new_n220), .B1(new_n226), .B2(new_n284), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G33), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n364), .A2(new_n238), .A3(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n290), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n279), .B1(G244), .B2(new_n282), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n359), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G179), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(G200), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n359), .C1(new_n344), .C2(new_n368), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n348), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n307), .A2(new_n343), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n349), .A2(new_n357), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n350), .A2(new_n331), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(KEYINPUT75), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(KEYINPUT75), .B2(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n259), .A2(new_n266), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n201), .A2(new_n202), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n204), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n262), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT71), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n390), .A3(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n361), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n232), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n392), .B2(new_n232), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT16), .B(new_n387), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n257), .ZN(new_n398));
  AOI21_X1  g0198(.A(G20), .B1(new_n361), .B2(new_n363), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT72), .B1(new_n399), .B2(KEYINPUT7), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n393), .C1(new_n284), .C2(G20), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT71), .B(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n363), .B1(new_n404), .B2(G33), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n393), .A2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(G68), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n400), .A2(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT73), .B1(new_n411), .B2(new_n202), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n412), .A3(new_n387), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n398), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n384), .B1(new_n415), .B2(KEYINPUT74), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n202), .B1(new_n403), .B2(new_n407), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n387), .B1(new_n417), .B2(new_n409), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n411), .A2(KEYINPUT73), .A3(new_n202), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n398), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n288), .A2(new_n285), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G226), .B2(new_n285), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n392), .A2(new_n426), .B1(new_n273), .B2(new_n221), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n290), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT77), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n279), .B1(G232), .B2(new_n282), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n344), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n293), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n416), .A2(new_n424), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g0235(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(KEYINPUT78), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n416), .A2(new_n424), .A3(new_n434), .A4(new_n441), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n438), .B1(new_n437), .B2(new_n442), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n430), .A2(new_n303), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n429), .A2(new_n445), .B1(new_n369), .B2(new_n432), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n420), .A2(KEYINPUT74), .A3(new_n421), .ZN(new_n447));
  INV_X1    g0247(.A(new_n384), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n415), .A2(KEYINPUT74), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT18), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n416), .A2(new_n424), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n446), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n443), .A2(new_n444), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n375), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n268), .A2(G33), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n267), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT25), .B1(new_n266), .B2(new_n226), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n461), .A2(new_n226), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n221), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n391), .A2(new_n232), .A3(new_n361), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n232), .A2(G87), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n364), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n232), .B2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n273), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n472), .A2(new_n473), .B1(new_n475), .B2(new_n232), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n468), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT86), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n257), .B1(new_n478), .B2(KEYINPUT24), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n477), .A2(KEYINPUT86), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT24), .A3(new_n478), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n465), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT88), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n276), .A2(G1), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G264), .A3(new_n275), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n290), .B1(new_n486), .B2(new_n485), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT87), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(G264), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n222), .A2(new_n285), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(G257), .B2(new_n285), .ZN(new_n494));
  INV_X1    g0294(.A(G294), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n392), .A2(new_n494), .B1(new_n273), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n489), .A2(new_n492), .B1(new_n496), .B2(new_n290), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n275), .A2(G274), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n487), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n484), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(new_n484), .A3(new_n500), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(G169), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n497), .A2(G179), .A3(new_n500), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n483), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n503), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n344), .B1(new_n507), .B2(new_n501), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n497), .A2(new_n500), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n293), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n506), .B1(new_n483), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n513));
  OR3_X1    g0313(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n474), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT84), .B1(new_n461), .B2(new_n474), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G283), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n517), .B(new_n232), .C1(G33), .C2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n257), .C1(new_n232), .C2(G116), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT20), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n232), .A2(G116), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n522), .A2(new_n523), .B1(new_n356), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G169), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n499), .B1(new_n490), .B2(G270), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n391), .A2(new_n361), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G257), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n227), .B2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n364), .A2(G303), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n275), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n530), .A3(new_n535), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n513), .B1(new_n527), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n369), .B1(new_n516), .B2(new_n525), .ZN(new_n541));
  INV_X1    g0341(.A(new_n513), .ZN(new_n542));
  INV_X1    g0342(.A(new_n538), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n543), .A2(new_n536), .A3(new_n275), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n541), .B(new_n542), .C1(new_n544), .C2(new_n529), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n539), .A2(G179), .A3(new_n526), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n540), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n516), .B(new_n525), .C1(new_n539), .C2(new_n293), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n544), .A2(new_n344), .A3(new_n529), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  INV_X1    g0352(.A(new_n486), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT80), .B1(new_n498), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n275), .A2(new_n555), .A3(G274), .A4(new_n486), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n486), .A2(new_n222), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n554), .A2(new_n556), .B1(new_n275), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G238), .A2(G1698), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n225), .B2(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n531), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n475), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n275), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n552), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n290), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT81), .A3(new_n558), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n568), .A3(new_n303), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n531), .A2(new_n232), .A3(G68), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n221), .B1(new_n310), .B2(new_n232), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n260), .A2(KEYINPUT19), .A3(new_n518), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n352), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n257), .B1(new_n266), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n352), .B(KEYINPUT82), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n461), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n565), .A2(new_n568), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n569), .B(new_n580), .C1(new_n581), .C2(G169), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n565), .A2(new_n568), .A3(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n267), .A2(G87), .A3(new_n460), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n585), .C1(new_n581), .C2(new_n293), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n225), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT4), .B1(new_n531), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n517), .C1(new_n222), .C2(new_n287), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n290), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n490), .A2(G257), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n500), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n369), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n518), .A3(G107), .ZN(new_n596));
  XNOR2_X1  g0396(.A(G97), .B(G107), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n598), .A2(new_n232), .B1(new_n208), .B2(new_n263), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n408), .B2(G107), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(new_n349), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n266), .A2(new_n518), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n461), .B2(new_n518), .ZN(new_n603));
  OAI221_X1 g0403(.A(new_n594), .B1(G179), .B2(new_n593), .C1(new_n601), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n600), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n603), .B1(new_n605), .B2(new_n257), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n593), .A2(G200), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n344), .C2(new_n593), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n582), .A2(new_n586), .A3(new_n604), .A4(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n459), .A2(new_n512), .A3(new_n551), .A4(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n444), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n612));
  INV_X1    g0412(.A(new_n348), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n342), .B1(new_n613), .B2(new_n371), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n456), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n305), .B1(new_n617), .B2(new_n301), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n547), .A2(KEYINPUT89), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n540), .A2(new_n624), .A3(new_n545), .A4(new_n546), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n506), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n608), .A2(new_n604), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n511), .A2(new_n483), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n559), .A2(new_n564), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n569), .B(new_n580), .C1(G169), .C2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n559), .B2(new_n564), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n585), .A2(new_n583), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n628), .A2(new_n629), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n506), .B1(new_n623), .B2(new_n625), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n636), .A3(new_n631), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT90), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n594), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n593), .A2(G179), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n642), .A2(new_n606), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n582), .A3(new_n586), .A4(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n633), .A2(new_n635), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n604), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n645), .B(KEYINPUT91), .C1(new_n647), .C2(KEYINPUT26), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(KEYINPUT91), .ZN(new_n649));
  INV_X1    g0449(.A(new_n633), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n638), .A2(new_n641), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n459), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n622), .A2(new_n653), .ZN(G369));
  NAND2_X1  g0454(.A1(new_n356), .A2(new_n232), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT93), .ZN(new_n657));
  OAI21_X1  g0457(.A(G213), .B1(new_n655), .B2(KEYINPUT27), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n526), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT94), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n551), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n626), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n662), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n512), .B1(new_n483), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n627), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n547), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n662), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n674), .A2(new_n512), .B1(new_n506), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n216), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n571), .A2(new_n221), .A3(new_n474), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n678), .A2(new_n268), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n235), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT28), .Z(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n652), .B2(new_n669), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n640), .B1(new_n673), .B2(new_n627), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT26), .B1(new_n646), .B2(new_n604), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n644), .A2(new_n582), .A3(new_n586), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n686), .B(new_n633), .C1(KEYINPUT26), .C2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n669), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n609), .A2(new_n512), .A3(new_n551), .A4(new_n669), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT31), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n565), .A2(new_n568), .A3(new_n497), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT95), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n565), .A2(new_n568), .A3(KEYINPUT95), .A4(new_n497), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n591), .A2(new_n592), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n539), .A2(G179), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n695), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n698), .B2(new_n699), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT30), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n632), .A2(G179), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n706), .A2(new_n509), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n537), .A2(new_n538), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n528), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n707), .A2(KEYINPUT96), .A3(new_n709), .A4(new_n593), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n509), .A3(new_n706), .A4(new_n593), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT96), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n703), .A2(new_n705), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n662), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n694), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n662), .A2(KEYINPUT31), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n703), .A2(new_n711), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n705), .ZN(new_n719));
  OAI21_X1  g0519(.A(G330), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n692), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n682), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n214), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n268), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n678), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n231), .B1(G20), .B2(new_n369), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n232), .A2(G179), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT99), .B(G159), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT32), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n232), .A2(new_n303), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n731), .A2(new_n344), .A3(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n741), .A2(G68), .B1(new_n743), .B2(G107), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n344), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n232), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G97), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n221), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n744), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n737), .A2(KEYINPUT32), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n740), .A2(new_n344), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n753), .B1(new_n205), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n739), .A2(new_n732), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n739), .A2(G190), .A3(new_n293), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n284), .B1(new_n757), .B2(new_n208), .C1(new_n201), .C2(new_n758), .ZN(new_n759));
  OR4_X1    g0559(.A1(new_n738), .A2(new_n752), .A3(new_n756), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G322), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n364), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n762), .B(new_n764), .C1(G329), .C2(new_n734), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n754), .A2(G326), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G294), .A2(new_n747), .B1(new_n741), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n749), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G303), .B1(new_n743), .B2(G283), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n730), .B1(new_n760), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n729), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n254), .A2(new_n276), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n531), .A2(new_n677), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n276), .B2(new_n235), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n781), .B2(new_n780), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n677), .A2(new_n364), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G355), .B1(new_n474), .B2(new_n677), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n728), .B(new_n772), .C1(new_n776), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n775), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n666), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT100), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n666), .A2(G330), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n791), .A2(new_n667), .A3(new_n728), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n652), .A2(new_n669), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n373), .B1(new_n669), .B2(new_n359), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n371), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n371), .A2(new_n662), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n652), .A2(new_n669), .A3(new_n800), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n727), .B1(new_n804), .B2(new_n720), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n720), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n730), .A2(new_n774), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n727), .B1(G77), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n758), .ZN(new_n809));
  INV_X1    g0609(.A(new_n757), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n809), .A2(G143), .B1(new_n810), .B2(new_n736), .ZN(new_n811));
  INV_X1    g0611(.A(new_n741), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n261), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G137), .B2(new_n754), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n743), .A2(G68), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n205), .B2(new_n749), .C1(new_n201), .C2(new_n746), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n392), .B(new_n818), .C1(G132), .C2(new_n734), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n812), .B1(new_n755), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G107), .B2(new_n769), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n758), .A2(new_n495), .B1(new_n733), .B2(new_n763), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n284), .B(new_n825), .C1(G116), .C2(new_n810), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n743), .A2(G87), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n748), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n820), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n808), .B1(new_n829), .B2(new_n729), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n800), .B2(new_n774), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n806), .A2(new_n831), .ZN(G384));
  INV_X1    g0632(.A(new_n598), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT35), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT35), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n834), .A2(G116), .A3(new_n233), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT36), .Z(new_n837));
  OR3_X1    g0637(.A1(new_n234), .A2(new_n208), .A3(new_n385), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n268), .B(G13), .C1(new_n838), .C2(new_n250), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n324), .A2(G169), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT14), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n317), .B1(new_n843), .B2(new_n325), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT102), .B1(new_n844), .B2(new_n340), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT102), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n328), .A2(new_n846), .A3(new_n341), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n669), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n453), .A2(new_n659), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(new_n451), .A4(new_n435), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n387), .B1(new_n395), .B2(new_n396), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n854), .A2(new_n414), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n381), .B(new_n379), .C1(new_n855), .C2(new_n398), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n446), .B2(new_n659), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n435), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n659), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT38), .B(new_n860), .C1(new_n457), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT106), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n611), .A2(new_n616), .A3(new_n612), .ZN(new_n865));
  INV_X1    g0665(.A(new_n861), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n867), .A2(KEYINPUT106), .A3(KEYINPUT38), .A4(new_n860), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n851), .A2(new_n451), .A3(new_n435), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n853), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n437), .A2(new_n442), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n873), .A2(new_n452), .A3(new_n455), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n874), .B2(new_n851), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n864), .A2(new_n868), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(KEYINPUT107), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT107), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n864), .A2(new_n868), .A3(new_n880), .A4(new_n877), .ZN(new_n881));
  INV_X1    g0681(.A(new_n862), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n867), .B2(new_n860), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n850), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n799), .B(KEYINPUT101), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n803), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n340), .A2(new_n669), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n328), .B2(new_n613), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n613), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n845), .A2(new_n847), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n845), .A2(new_n847), .A3(new_n892), .A4(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT104), .ZN(new_n900));
  INV_X1    g0700(.A(new_n883), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n899), .A2(new_n900), .B1(new_n901), .B2(new_n862), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n888), .A2(KEYINPUT104), .A3(new_n898), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n902), .A2(new_n903), .B1(new_n456), .B2(new_n660), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n886), .A2(new_n904), .ZN(new_n905));
  OR3_X1    g0705(.A1(new_n684), .A2(new_n458), .A3(new_n691), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n622), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n710), .B(new_n713), .C1(new_n704), .C2(KEYINPUT30), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n704), .A2(KEYINPUT30), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT31), .B(new_n662), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT108), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n714), .A2(KEYINPUT108), .A3(KEYINPUT31), .A4(new_n662), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n913), .A2(new_n914), .B1(new_n694), .B2(new_n715), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n897), .A2(new_n915), .A3(new_n801), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n883), .B2(new_n882), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n875), .A2(new_n876), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n864), .A2(new_n868), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n915), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n459), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(G330), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n908), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n268), .B2(new_n724), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n908), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n840), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n674), .A2(new_n512), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n671), .B2(new_n674), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT111), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n667), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n667), .A2(new_n935), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n722), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n630), .B1(new_n606), .B2(new_n669), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n644), .A2(new_n662), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n675), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT45), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n675), .A2(new_n943), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n672), .A2(KEYINPUT110), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n721), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n953));
  XNOR2_X1  g0753(.A(new_n678), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n725), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n943), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n933), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n604), .B1(new_n941), .B2(new_n627), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n958), .A2(KEYINPUT42), .B1(new_n669), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n585), .A2(new_n669), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n646), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n650), .A2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n959), .A2(new_n961), .B1(KEYINPUT43), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n966), .B(new_n967), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n672), .A2(new_n956), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n955), .A2(new_n970), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n776), .B1(new_n216), .B2(new_n577), .C1(new_n779), .C2(new_n244), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n727), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n758), .A2(new_n261), .B1(new_n757), .B2(new_n205), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n364), .B(new_n974), .C1(G137), .C2(new_n734), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n747), .A2(G68), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n741), .A2(new_n736), .B1(new_n769), .B2(G58), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n754), .A2(G143), .B1(new_n743), .B2(G77), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n755), .A2(new_n763), .B1(new_n226), .B2(new_n746), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G294), .B2(new_n741), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n758), .A2(new_n822), .B1(new_n757), .B2(new_n821), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G317), .B2(new_n734), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n531), .B1(G97), .B2(new_n743), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n749), .A2(new_n474), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n979), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT47), .Z(new_n989));
  OAI221_X1 g0789(.A(new_n973), .B1(new_n730), .B2(new_n989), .C1(new_n965), .C2(new_n788), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n971), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT112), .Z(G387));
  NAND2_X1  g0792(.A1(new_n938), .A2(new_n721), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n940), .A2(new_n678), .A3(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n809), .A2(G317), .B1(new_n810), .B2(G303), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n755), .B2(new_n761), .C1(new_n763), .C2(new_n812), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT113), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT48), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n747), .A2(G283), .B1(new_n769), .B2(G294), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n531), .B1(G326), .B2(new_n734), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n474), .B2(new_n742), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT114), .Z(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n749), .A2(new_n208), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G159), .B2(new_n754), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n259), .B2(new_n812), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n579), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n747), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n758), .A2(new_n205), .B1(new_n733), .B2(new_n261), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G68), .B2(new_n810), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n392), .B1(G97), .B2(new_n743), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1004), .A2(new_n1009), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT115), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n730), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n671), .A2(new_n788), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n241), .A2(new_n276), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1024), .A2(new_n778), .B1(new_n679), .B2(new_n784), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n350), .B2(new_n205), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n259), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n276), .B1(new_n202), .B2(new_n208), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n679), .A4(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1025), .A2(new_n1030), .B1(G107), .B2(new_n216), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n728), .B1(new_n1031), .B2(new_n776), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1022), .A2(new_n1023), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n939), .B2(new_n726), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n994), .A2(new_n1034), .ZN(G393));
  OAI21_X1  g0835(.A(new_n678), .B1(new_n940), .B2(new_n950), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n948), .B(new_n672), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n722), .B2(new_n939), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT117), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1037), .A2(new_n726), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n776), .B1(new_n518), .B2(new_n216), .C1(new_n779), .C2(new_n248), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n727), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n746), .A2(new_n208), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n827), .B1(new_n202), .B2(new_n749), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G50), .C2(new_n741), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n350), .A2(new_n810), .B1(new_n734), .B2(G143), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G150), .A2(new_n754), .B1(new_n809), .B2(G159), .ZN(new_n1048));
  XOR2_X1   g0848(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1046), .A2(new_n531), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G317), .A2(new_n754), .B1(new_n809), .B2(G311), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n812), .A2(new_n822), .B1(new_n474), .B2(new_n746), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n364), .B1(new_n733), .B2(new_n761), .C1(new_n495), .C2(new_n757), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n226), .A2(new_n742), .B1(new_n749), .B2(new_n821), .ZN(new_n1056));
  OR3_X1    g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1051), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1043), .B1(new_n1058), .B2(new_n729), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n943), .B2(new_n788), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1041), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1040), .A2(new_n1062), .ZN(G390));
  NAND2_X1  g0863(.A1(new_n878), .A2(KEYINPUT107), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n899), .A2(new_n849), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1064), .A2(new_n884), .A3(new_n881), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n799), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n689), .B2(new_n798), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n850), .B1(new_n898), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n921), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n897), .A2(new_n801), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(G330), .A3(new_n924), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(G330), .B(new_n800), .C1(new_n716), .C2(new_n719), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1066), .B(new_n1070), .C1(new_n897), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n924), .A2(G330), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n906), .B1(new_n458), .B2(new_n1079), .C1(new_n620), .C2(new_n621), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(new_n897), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1076), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1068), .B1(new_n1083), .B2(new_n898), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n897), .B1(new_n1079), .B2(new_n801), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1082), .A2(new_n888), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1078), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1075), .A2(new_n1077), .A3(new_n1087), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n678), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1064), .A2(new_n773), .A3(new_n884), .A4(new_n881), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n727), .B1(new_n350), .B2(new_n807), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n749), .A2(new_n261), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT53), .ZN(new_n1094));
  INV_X1    g0894(.A(G132), .ZN(new_n1095));
  INV_X1    g0895(.A(G125), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n758), .A2(new_n1095), .B1(new_n733), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n284), .B1(new_n757), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n754), .A2(G128), .B1(new_n743), .B2(G50), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G159), .A2(new_n747), .B1(new_n741), .B2(G137), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1094), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT118), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT118), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1044), .B1(G283), .B2(new_n754), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n226), .B2(new_n812), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n758), .A2(new_n474), .B1(new_n733), .B2(new_n495), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n284), .B(new_n1108), .C1(G97), .C2(new_n810), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n751), .A3(new_n817), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1104), .B(new_n1105), .C1(new_n1107), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1092), .B1(new_n1111), .B2(new_n729), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1078), .A2(new_n726), .B1(new_n1091), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1090), .A2(new_n1113), .ZN(G378));
  INV_X1    g0914(.A(new_n1080), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1089), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n919), .A2(new_n922), .A3(new_n1117), .A4(G330), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n905), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n271), .A2(new_n659), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n307), .B(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1122), .B(new_n1123), .Z(new_n1124));
  NAND3_X1  g0924(.A1(new_n919), .A2(new_n922), .A3(G330), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(KEYINPUT121), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n886), .A2(new_n1118), .A3(new_n904), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1120), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1126), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n886), .A2(new_n1118), .A3(new_n904), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1118), .B1(new_n886), .B2(new_n904), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1116), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT122), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1116), .A2(new_n1132), .A3(KEYINPUT57), .A4(new_n1128), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1138), .A2(new_n678), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1133), .A2(KEYINPUT122), .A3(new_n1134), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1132), .A2(new_n1128), .A3(new_n726), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n727), .B1(G50), .B2(new_n807), .ZN(new_n1143));
  AOI211_X1 g0943(.A(G33), .B(G41), .C1(new_n734), .C2(G124), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n742), .B2(new_n735), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n741), .A2(G132), .B1(new_n810), .B2(G137), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT120), .Z(new_n1147));
  NOR2_X1   g0947(.A1(new_n746), .A2(new_n261), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n758), .A2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n755), .A2(new_n1096), .B1(new_n749), .B2(new_n1098), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1145), .B1(new_n1153), .B2(KEYINPUT59), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(KEYINPUT59), .B2(new_n1153), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n531), .A2(G41), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G50), .B(new_n1156), .C1(new_n273), .C2(new_n274), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1013), .A2(new_n810), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n809), .A2(G107), .B1(new_n734), .B2(G283), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n976), .A3(new_n1156), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n742), .A2(new_n201), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n518), .A2(new_n812), .B1(new_n755), .B2(new_n474), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1160), .A2(new_n1010), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1157), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1155), .B(new_n1165), .C1(new_n1164), .C2(new_n1163), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1143), .B1(new_n1166), .B2(new_n729), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1124), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n774), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1142), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1141), .A2(new_n1171), .ZN(G375));
  INV_X1    g0972(.A(new_n1086), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n897), .A2(new_n773), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n727), .B1(G68), .B2(new_n807), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n741), .A2(G116), .B1(new_n810), .B2(G107), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT123), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n755), .A2(new_n495), .B1(new_n742), .B2(new_n208), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G97), .B2(new_n769), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n364), .B1(new_n733), .B2(new_n822), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G283), .B2(new_n809), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n1179), .A3(new_n1014), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G159), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n201), .A2(new_n742), .B1(new_n749), .B2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n531), .B1(new_n1149), .B2(new_n733), .C1(new_n261), .C2(new_n757), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G50), .C2(new_n747), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT124), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n809), .A2(G137), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n755), .B2(new_n1095), .C1(new_n812), .C2(new_n1098), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1175), .B1(new_n1190), .B2(new_n729), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1173), .A2(new_n726), .B1(new_n1174), .B2(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1087), .A2(new_n954), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1115), .A2(new_n1173), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(G381));
  NAND3_X1  g0995(.A1(new_n994), .A2(new_n793), .A3(new_n1034), .ZN(new_n1196));
  OR4_X1    g0996(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1196), .ZN(new_n1197));
  OR4_X1    g0997(.A1(G387), .A2(new_n1197), .A3(G375), .A4(G378), .ZN(G407));
  AOI21_X1  g0998(.A(KEYINPUT122), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1138), .A2(new_n678), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1170), .B1(new_n1201), .B2(new_n1140), .ZN(new_n1202));
  INV_X1    g1002(.A(G378), .ZN(new_n1203));
  INV_X1    g1003(.A(G213), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(G343), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(G407), .A2(G213), .A3(new_n1206), .ZN(G409));
  NAND3_X1  g1007(.A1(new_n1141), .A2(G378), .A3(new_n1171), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1133), .A2(new_n954), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1171), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1205), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1205), .A2(G2897), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1080), .A2(new_n1086), .A3(KEYINPUT60), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1215), .A2(new_n678), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT60), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1087), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1218), .B2(new_n1194), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G384), .B1(new_n1219), .B2(new_n1192), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(G384), .A3(new_n1192), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1214), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1222), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1224), .A2(new_n1220), .A3(new_n1213), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT125), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1213), .B1(new_n1224), .B2(new_n1220), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1221), .A2(new_n1222), .A3(new_n1214), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT126), .B1(new_n1212), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G378), .B1(new_n1171), .B2(new_n1209), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1202), .B2(G378), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1233), .B(new_n1234), .C1(new_n1236), .C2(new_n1205), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1224), .A2(new_n1220), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1212), .A2(KEYINPUT63), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G393), .A2(G396), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1196), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT127), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(KEYINPUT127), .A3(new_n1196), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G390), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT112), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(G390), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n971), .A3(new_n990), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1247), .B(new_n991), .C1(G390), .C2(new_n1248), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1205), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1239), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1253), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1238), .A2(new_n1240), .A3(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1251), .B1(new_n1212), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1212), .B2(new_n1239), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1260), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1259), .B1(new_n1265), .B2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1203), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1208), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1270), .A2(new_n1239), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1239), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1266), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(new_n1267), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G402));
endmodule


