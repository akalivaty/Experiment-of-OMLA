//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n208), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n202), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n221), .B(new_n226), .C1(KEYINPUT1), .C2(new_n216), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n218), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G58), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G97), .B(G107), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  OAI21_X1  g0043(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n244));
  INV_X1    g0044(.A(G150), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT67), .A2(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT8), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n206), .A2(G33), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n244), .B1(new_n245), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n224), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n254), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n205), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  MUX2_X1   g0059(.A(new_n256), .B(new_n259), .S(G50), .Z(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT9), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n265), .B1(new_n266), .B2(new_n263), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  OAI211_X1 g0076(.A(G1), .B(G13), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT66), .B1(new_n273), .B2(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n281), .B1(new_n286), .B2(G226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n274), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n262), .B(new_n289), .C1(new_n290), .C2(new_n288), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n274), .A2(new_n295), .A3(new_n287), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n261), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n259), .A2(new_n249), .ZN(new_n299));
  INV_X1    g0099(.A(new_n256), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n249), .ZN(new_n301));
  INV_X1    g0101(.A(G58), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G20), .B1(new_n304), .B2(new_n201), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n246), .A2(G159), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n263), .B2(G20), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n303), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n308), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT16), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n263), .A2(new_n309), .A3(G20), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n267), .A2(KEYINPUT73), .A3(new_n268), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n311), .B2(new_n312), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n324), .A3(new_n206), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n325), .B2(new_n309), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT16), .B(new_n308), .C1(new_n326), .C2(new_n303), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n254), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n301), .B1(new_n320), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n271), .A2(new_n264), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(G226), .B2(new_n264), .C1(new_n311), .C2(new_n312), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n273), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n277), .A2(G232), .A3(new_n284), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n280), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT75), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n277), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT75), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n339), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n293), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n339), .A2(new_n336), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n295), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n329), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT18), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n338), .B2(new_n341), .ZN(new_n350));
  INV_X1    g0150(.A(new_n343), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(G190), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT16), .ZN(new_n353));
  INV_X1    g0153(.A(new_n319), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n317), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n254), .A3(new_n327), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n356), .A3(new_n301), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT17), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n329), .A2(new_n346), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n301), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n327), .A2(new_n254), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(KEYINPUT17), .A3(new_n352), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n348), .A2(new_n359), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G13), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(G1), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT68), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(G77), .ZN(new_n373));
  INV_X1    g0173(.A(new_n372), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n254), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n375), .A2(G77), .A3(new_n258), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT8), .B(G58), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n246), .B1(G20), .B2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n251), .B2(new_n380), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n373), .B(new_n376), .C1(new_n254), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n263), .A2(G232), .A3(new_n264), .ZN(new_n383));
  INV_X1    g0183(.A(G107), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n383), .B1(new_n384), .B2(new_n263), .C1(new_n270), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n273), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n281), .B1(new_n286), .B2(G244), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n382), .B1(new_n293), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n295), .A3(new_n388), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(G200), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n382), .B(new_n393), .C1(new_n290), .C2(new_n389), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n298), .A2(new_n366), .A3(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n264), .A2(G232), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n263), .B(new_n397), .C1(G226), .C2(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n277), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n273), .A2(new_n279), .A3(KEYINPUT66), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n283), .B1(new_n277), .B2(new_n284), .ZN(new_n403));
  OAI21_X1  g0203(.A(G238), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT69), .B1(new_n404), .B2(new_n280), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n385), .B1(new_n282), .B2(new_n285), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT69), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n406), .A2(new_n407), .A3(new_n281), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n401), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT71), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT13), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n407), .B1(new_n406), .B2(new_n281), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n404), .A2(KEYINPUT69), .A3(new_n280), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n400), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT71), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g0216(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n411), .A2(new_n416), .A3(G190), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n303), .A2(G20), .ZN(new_n420));
  INV_X1    g0220(.A(G50), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n251), .B2(new_n266), .C1(new_n247), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n254), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT11), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n375), .A2(G68), .A3(new_n258), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n368), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n427), .A2(KEYINPUT12), .A3(new_n420), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n374), .A2(new_n303), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(KEYINPUT12), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n414), .A2(new_n417), .ZN(new_n432));
  INV_X1    g0232(.A(new_n417), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n433), .B(new_n400), .C1(new_n412), .C2(new_n413), .ZN(new_n434));
  OAI21_X1  g0234(.A(G200), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n419), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(G169), .C1(new_n432), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT72), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n409), .A2(new_n433), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n418), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT72), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n437), .A4(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(G169), .B1(new_n432), .B2(new_n434), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n411), .A2(new_n416), .A3(G179), .A4(new_n418), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n439), .A2(new_n443), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n431), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n436), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n396), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G41), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n205), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n205), .A4(G45), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n273), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G270), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n263), .A2(G264), .A3(G1698), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n263), .A2(G257), .A3(new_n264), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n313), .A2(G303), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n273), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n276), .A2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n205), .A2(G45), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n454), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n452), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n467), .A2(new_n457), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G274), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n273), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n459), .A2(new_n464), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n374), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n205), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n372), .A2(G116), .A3(new_n257), .A4(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n253), .A2(new_n224), .B1(G20), .B2(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n206), .C1(G33), .C2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n478), .A2(KEYINPUT20), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT20), .B1(new_n478), .B2(new_n481), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n475), .B(new_n477), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n473), .A2(G169), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT21), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(KEYINPUT81), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n459), .A2(new_n464), .A3(new_n472), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G179), .A3(new_n484), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n484), .B1(new_n473), .B2(G200), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n290), .B2(new_n473), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n487), .A2(new_n489), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n264), .C1(new_n311), .C2(new_n312), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT76), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n269), .A2(G250), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n479), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n495), .B2(new_n496), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n273), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(G257), .A2(new_n458), .B1(new_n469), .B2(new_n471), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n480), .A3(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n508), .A2(new_n206), .B1(new_n266), .B2(new_n247), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n384), .B1(new_n310), .B2(new_n314), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n254), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n256), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n257), .A2(new_n256), .A3(new_n476), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n480), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n504), .A2(new_n293), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n502), .A2(new_n503), .A3(new_n295), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n504), .A2(G200), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n507), .A2(new_n505), .ZN(new_n522));
  INV_X1    g0322(.A(new_n506), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(G20), .B1(G77), .B2(new_n246), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n310), .A2(new_n314), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n515), .B1(new_n528), .B2(new_n254), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n521), .B(new_n529), .C1(new_n290), .C2(new_n504), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n520), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n206), .B(G68), .C1(new_n311), .C2(new_n312), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n251), .B2(new_n480), .ZN(new_n534));
  OR2_X1    g0334(.A1(KEYINPUT79), .A2(G87), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  NAND2_X1  g0336(.A1(KEYINPUT79), .A2(G87), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n540), .A2(new_n206), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n532), .B(new_n534), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n254), .B1(new_n374), .B2(new_n380), .ZN(new_n543));
  INV_X1    g0343(.A(new_n514), .ZN(new_n544));
  INV_X1    g0344(.A(new_n380), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT80), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n537), .ZN(new_n548));
  NOR2_X1   g0348(.A1(KEYINPUT79), .A2(G87), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n541), .B1(new_n536), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n532), .A2(new_n534), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n254), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n374), .A2(new_n380), .ZN(new_n554));
  AND4_X1   g0354(.A1(KEYINPUT80), .A2(new_n553), .A3(new_n546), .A4(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G238), .B(new_n264), .C1(new_n311), .C2(new_n312), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT78), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT78), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n263), .A2(new_n558), .A3(G238), .A4(new_n264), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n263), .A2(G244), .A3(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n273), .ZN(new_n563));
  INV_X1    g0363(.A(G250), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n466), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n205), .A2(new_n470), .A3(G45), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n277), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n293), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n567), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n295), .B(new_n569), .C1(new_n562), .C2(new_n273), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n547), .A2(new_n555), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n562), .B2(new_n273), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G190), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n544), .A2(G87), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n553), .A2(new_n574), .A3(new_n554), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n575), .C1(new_n349), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n494), .A2(new_n531), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT86), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n467), .A2(new_n457), .A3(new_n468), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(G264), .A3(new_n277), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT84), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT84), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n458), .A2(new_n583), .A3(G264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n586));
  OAI211_X1 g0386(.A(G250), .B(new_n264), .C1(new_n311), .C2(new_n312), .ZN(new_n587));
  INV_X1    g0387(.A(G294), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n587), .C1(new_n275), .C2(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n471), .A2(new_n469), .B1(new_n589), .B2(new_n273), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(G179), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n583), .B1(new_n458), .B2(G264), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n583), .A2(new_n580), .A3(G264), .A4(new_n277), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n590), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n593), .B1(new_n585), .B2(new_n590), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n599), .B2(G169), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n384), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT25), .B1(new_n300), .B2(new_n384), .ZN(new_n603));
  XOR2_X1   g0403(.A(new_n602), .B(new_n603), .Z(new_n604));
  NAND2_X1  g0404(.A1(new_n544), .A2(G107), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n263), .A2(new_n206), .A3(G87), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT22), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT23), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n384), .A3(G20), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT82), .ZN(new_n612));
  OAI221_X1 g0412(.A(new_n610), .B1(G20), .B2(new_n560), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n612), .B2(new_n611), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n615), .B(KEYINPUT24), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n606), .B1(new_n616), .B2(new_n254), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n579), .B1(new_n600), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n585), .A2(new_n590), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT85), .ZN(new_n620));
  AOI21_X1  g0420(.A(G190), .B1(new_n620), .B2(new_n596), .ZN(new_n621));
  AOI21_X1  g0421(.A(G200), .B1(new_n585), .B2(new_n590), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n617), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(G169), .A3(new_n596), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n591), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n626), .A3(KEYINPUT86), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n578), .A2(new_n618), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n450), .A2(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n297), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n364), .A2(KEYINPUT18), .A3(new_n345), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n360), .B1(new_n329), .B2(new_n346), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n436), .A2(new_n392), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n448), .B2(new_n447), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n357), .A2(new_n358), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT17), .B1(new_n364), .B2(new_n352), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n633), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT88), .ZN(new_n641));
  INV_X1    g0441(.A(new_n292), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n640), .B2(KEYINPUT88), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n630), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT87), .B1(new_n568), .B2(new_n570), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n563), .A2(G179), .A3(new_n567), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n646), .B(new_n647), .C1(new_n293), .C2(new_n572), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n553), .A2(new_n546), .A3(new_n554), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT80), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n543), .A2(KEYINPUT80), .A3(new_n546), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n645), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n571), .A2(new_n576), .A3(new_n519), .A4(new_n517), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n655), .B1(KEYINPUT26), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(new_n576), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AOI21_X1  g0460(.A(G169), .B1(new_n502), .B2(new_n503), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n518), .A2(new_n661), .A3(new_n529), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n531), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n623), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n624), .B2(new_n626), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n657), .B(new_n663), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n644), .B1(new_n450), .B2(new_n669), .ZN(G369));
  OR3_X1    g0470(.A1(new_n427), .A2(KEYINPUT27), .A3(G20), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT27), .B1(new_n427), .B2(G20), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n624), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n618), .A2(new_n627), .A3(new_n623), .A4(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n600), .A2(new_n617), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n675), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n666), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n484), .A2(new_n675), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n493), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n681), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n681), .A2(new_n675), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(new_n618), .A3(new_n623), .A4(new_n627), .ZN(new_n688));
  INV_X1    g0488(.A(new_n675), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n219), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n539), .A2(new_n474), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n696), .A2(new_n697), .B1(new_n222), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n668), .A2(new_n689), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT90), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT90), .ZN(new_n703));
  AOI211_X1 g0503(.A(new_n703), .B(KEYINPUT29), .C1(new_n668), .C2(new_n689), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n618), .A2(new_n627), .A3(new_n681), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n665), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n618), .A2(new_n627), .A3(KEYINPUT93), .A4(new_n681), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n654), .A2(new_n662), .A3(KEYINPUT26), .A4(new_n576), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT92), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n656), .A2(new_n715), .A3(new_n660), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n656), .B2(new_n660), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n713), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n655), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n675), .B1(new_n711), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n705), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n504), .A2(new_n295), .A3(new_n473), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n589), .A2(new_n273), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n585), .A2(new_n725), .A3(new_n572), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n727), .A3(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n490), .A2(G179), .A3(new_n502), .A4(new_n503), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n490), .A2(G179), .A3(new_n572), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n619), .A3(new_n504), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n675), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(new_n733), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT89), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(new_n733), .A3(KEYINPUT89), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n728), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n675), .A2(KEYINPUT31), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n628), .B2(new_n675), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n699), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n685), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n367), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n205), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n694), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n684), .ZN(new_n754));
  INV_X1    g0554(.A(new_n752), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n224), .B1(G20), .B2(new_n293), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n322), .A2(new_n324), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n693), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n278), .B2(new_n223), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT96), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n239), .A2(new_n278), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT95), .Z(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(KEYINPUT96), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n313), .B(new_n693), .C1(KEYINPUT94), .C2(G355), .ZN(new_n771));
  OR2_X1    g0571(.A1(G355), .A2(KEYINPUT94), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(new_n474), .B2(new_n693), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n761), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n206), .A2(G179), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n263), .B1(new_n778), .B2(G329), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n206), .A2(new_n295), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n776), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n349), .A2(G190), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n206), .A3(new_n295), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n779), .B1(new_n780), .B2(new_n782), .C1(new_n783), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n781), .A2(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G190), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n775), .A2(new_n290), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n789), .A2(new_n790), .B1(new_n792), .B2(G283), .ZN(new_n793));
  INV_X1    g0593(.A(G303), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n788), .A2(new_n290), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n793), .B1(new_n794), .B2(new_n795), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(G20), .B1(new_n784), .B2(G179), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT97), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n787), .B(new_n799), .C1(G294), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n777), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n792), .A2(G107), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(new_n421), .C2(new_n798), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n804), .A2(new_n480), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n263), .B1(new_n266), .B2(new_n782), .C1(new_n786), .C2(new_n302), .ZN(new_n813));
  INV_X1    g0613(.A(new_n789), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n814), .A2(new_n303), .B1(new_n550), .B2(new_n795), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n755), .B(new_n774), .C1(new_n759), .C2(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n758), .B(KEYINPUT98), .Z(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n684), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n754), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  OAI21_X1  g0622(.A(new_n394), .B1(new_n382), .B2(new_n689), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n392), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n390), .A2(new_n391), .A3(new_n689), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n700), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n826), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(new_n668), .A3(new_n689), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n752), .B1(new_n830), .B2(new_n744), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n744), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n759), .A2(new_n756), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n755), .B1(new_n266), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n759), .ZN(new_n835));
  INV_X1    g0635(.A(new_n762), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G132), .B2(new_n778), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n421), .B2(new_n795), .C1(new_n303), .C2(new_n791), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G58), .B2(new_n805), .ZN(new_n839));
  INV_X1    g0639(.A(new_n782), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(G159), .B1(new_n785), .B2(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n798), .B2(new_n842), .C1(new_n245), .C2(new_n814), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT34), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n313), .B1(new_n795), .B2(new_n384), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n792), .A2(G87), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n798), .B2(new_n794), .C1(new_n848), .C2(new_n814), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n840), .A2(G116), .B1(new_n785), .B2(G294), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n780), .B2(new_n777), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n812), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n839), .A2(new_n844), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n834), .B1(new_n835), .B2(new_n853), .C1(new_n828), .C2(new_n757), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n832), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  OR2_X1    g0656(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n225), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  OR3_X1    g0660(.A1(new_n222), .A2(new_n266), .A3(new_n304), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n421), .A2(G68), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT100), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n205), .B(G13), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n673), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n633), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n448), .B(new_n675), .C1(new_n447), .C2(new_n436), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n431), .A2(new_n689), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n870), .B(new_n436), .C1(new_n447), .C2(new_n448), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n825), .B2(new_n829), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n308), .B1(new_n326), .B2(new_n303), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n353), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n254), .A3(new_n327), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n301), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n866), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n638), .B2(new_n633), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n352), .A2(new_n356), .A3(new_n301), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n345), .A2(new_n673), .B1(new_n877), .B2(new_n301), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n329), .A2(new_n866), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n347), .A2(new_n884), .A3(new_n357), .A4(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n874), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n886), .ZN(new_n889));
  INV_X1    g0689(.A(new_n366), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT38), .B(new_n889), .C1(new_n890), .C2(new_n879), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n867), .B1(new_n873), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n447), .A2(new_n448), .A3(new_n689), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n347), .A2(new_n884), .A3(new_n357), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(new_n885), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n884), .B1(new_n638), .B2(new_n633), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n874), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT101), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n891), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(new_n891), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT101), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n888), .B2(new_n891), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n895), .B(new_n902), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n893), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n450), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n705), .A3(new_n722), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n644), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n907), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n447), .A2(new_n448), .ZN(new_n912));
  INV_X1    g0712(.A(new_n436), .ZN(new_n913));
  INV_X1    g0713(.A(new_n870), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n868), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n735), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n628), .B2(new_n675), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n828), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT102), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n916), .A2(KEYINPUT102), .A3(new_n828), .A4(new_n919), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n899), .B2(new_n891), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n888), .A2(new_n891), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n908), .A2(new_n919), .ZN(new_n930));
  OAI21_X1  g0730(.A(G330), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n911), .A2(new_n932), .B1(new_n205), .B2(new_n749), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n911), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n865), .B1(new_n933), .B2(new_n934), .ZN(G367));
  OAI221_X1 g0735(.A(new_n760), .B1(new_n219), .B2(new_n380), .C1(new_n764), .C2(new_n235), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n936), .A2(new_n752), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n689), .A2(new_n575), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n655), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n658), .B2(new_n938), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n263), .B1(new_n421), .B2(new_n782), .C1(new_n786), .C2(new_n245), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n792), .A2(G77), .ZN(new_n942));
  INV_X1    g0742(.A(G143), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n798), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n941), .B(new_n944), .C1(G159), .C2(new_n789), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n795), .A2(new_n302), .B1(new_n777), .B2(new_n842), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n805), .A2(G68), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n945), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n762), .B1(new_n797), .B2(G311), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n789), .A2(G294), .B1(new_n792), .B2(G97), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n804), .C2(new_n384), .ZN(new_n953));
  XNOR2_X1  g0753(.A(KEYINPUT107), .B(G317), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n778), .A2(new_n954), .B1(new_n785), .B2(G303), .ZN(new_n955));
  INV_X1    g0755(.A(new_n795), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(KEYINPUT46), .A3(G116), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT46), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n795), .B2(new_n474), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n840), .A2(G283), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n955), .A2(new_n957), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n950), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  OAI221_X1 g0763(.A(new_n937), .B1(new_n819), .B2(new_n940), .C1(new_n963), .C2(new_n835), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n664), .B1(new_n529), .B2(new_n689), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n662), .A2(new_n675), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n691), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n691), .A2(new_n967), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n686), .ZN(new_n974));
  INV_X1    g0774(.A(new_n686), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n677), .A2(new_n679), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n688), .B1(new_n978), .B2(new_n687), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n748), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n723), .A2(new_n744), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT104), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n723), .A2(KEYINPUT104), .A3(new_n744), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n977), .B1(new_n985), .B2(KEYINPUT105), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT105), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n745), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n694), .B(KEYINPUT41), .Z(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT106), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT106), .ZN(new_n992));
  INV_X1    g0792(.A(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(new_n988), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n987), .B1(new_n983), .B2(new_n984), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n994), .A2(new_n995), .A3(new_n977), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n992), .B(new_n993), .C1(new_n996), .C2(new_n745), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n751), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n967), .A2(new_n688), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT42), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n965), .B1(new_n618), .B2(new_n627), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n689), .B1(new_n1001), .B2(new_n662), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n940), .B(KEYINPUT43), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n1003), .A2(KEYINPUT103), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT103), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n975), .A2(new_n967), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1009), .B(new_n1010), .Z(new_n1011));
  OAI21_X1  g0811(.A(new_n964), .B1(new_n998), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT109), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT109), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1015), .A2(new_n1018), .ZN(G387));
  INV_X1    g0819(.A(new_n980), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n695), .B1(new_n745), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n985), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n763), .B1(new_n232), .B2(new_n278), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n697), .A2(new_n219), .A3(new_n263), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n377), .A2(G50), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT110), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G45), .B(new_n697), .C1(G68), .C2(G77), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1025), .A2(new_n1031), .B1(new_n384), .B2(new_n693), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n752), .B1(new_n1032), .B2(new_n761), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n840), .A2(G303), .B1(new_n785), .B2(new_n954), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n798), .B2(new_n783), .C1(new_n780), .C2(new_n814), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n805), .A2(G283), .B1(G294), .B2(new_n956), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT49), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n836), .B1(new_n474), .B2(new_n791), .C1(new_n796), .C2(new_n777), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n814), .A2(new_n250), .B1(new_n266), .B2(new_n795), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G159), .B2(new_n797), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n805), .A2(new_n545), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n786), .A2(new_n421), .B1(new_n777), .B2(new_n245), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G68), .B2(new_n840), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n836), .B1(G97), .B2(new_n792), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1033), .B1(new_n1054), .B2(new_n759), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n978), .B2(new_n819), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1020), .B2(new_n750), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1022), .A2(new_n1058), .ZN(G393));
  NAND2_X1  g0859(.A1(new_n977), .A2(KEYINPUT112), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT112), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n974), .A2(new_n1061), .A3(new_n976), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n751), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n967), .A2(new_n758), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n797), .A2(G317), .B1(G311), .B2(new_n785), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT113), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n805), .A2(G116), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n313), .B1(new_n777), .B2(new_n783), .C1(new_n588), .C2(new_n782), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n810), .B1(new_n814), .B2(new_n794), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G283), .C2(new_n956), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n847), .B1(new_n303), .B2(new_n795), .C1(new_n814), .C2(new_n421), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n782), .A2(new_n377), .B1(new_n777), .B2(new_n943), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1074), .A2(new_n836), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n798), .A2(new_n245), .B1(new_n807), .B2(new_n786), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT51), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n805), .A2(G77), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n835), .B1(new_n1073), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n764), .A2(new_n242), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n761), .B(new_n1084), .C1(G97), .C2(new_n693), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1083), .A2(new_n755), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1064), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n695), .B1(new_n985), .B2(new_n977), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1063), .B(new_n1087), .C1(new_n996), .C2(new_n1089), .ZN(G390));
  OAI21_X1  g0890(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n829), .A2(new_n825), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n894), .B1(new_n1092), .B2(new_n872), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n711), .A2(new_n720), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n689), .A3(new_n824), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n872), .B1(new_n1096), .B2(new_n825), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT114), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n895), .B1(new_n899), .B2(new_n891), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n824), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n675), .B(new_n1102), .C1(new_n711), .C2(new_n720), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n825), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n916), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT114), .B1(new_n1105), .B2(new_n1099), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1094), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n919), .A2(G330), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n872), .A2(new_n1108), .A3(new_n826), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n916), .A2(new_n743), .A3(G330), .A4(new_n828), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1104), .B1(new_n721), .B2(new_n824), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n872), .B1(new_n1108), .B2(new_n826), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT115), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1117), .A2(new_n1121), .A3(new_n1111), .A4(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1109), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n872), .B1(new_n744), .B2(new_n826), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1092), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n450), .A2(new_n1108), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n644), .A2(new_n909), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1116), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1115), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1098), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n1099), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1107), .A2(new_n1109), .B1(new_n1137), .B2(new_n1113), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1120), .A2(new_n1122), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(new_n1131), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1140), .B2(new_n1116), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1141), .A3(new_n694), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT117), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1114), .A2(new_n751), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1124), .B1(new_n1137), .B2(new_n1094), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n750), .B1(new_n1137), .B2(new_n1113), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1110), .A2(KEYINPUT117), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1091), .A2(new_n756), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n786), .A2(new_n474), .B1(new_n782), .B2(new_n480), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n263), .B(new_n1151), .C1(G294), .C2(new_n778), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n789), .A2(G107), .B1(new_n792), .B2(G68), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n797), .A2(G283), .B1(new_n956), .B2(G87), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1152), .A2(new_n1080), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n840), .A2(new_n1157), .B1(new_n778), .B2(G125), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n245), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT53), .B1(new_n795), .B2(new_n245), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n313), .B1(new_n785), .B2(G132), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n797), .A2(G128), .B1(new_n792), .B2(G50), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n842), .B2(new_n814), .C1(new_n804), .C2(new_n807), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1155), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT118), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n835), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n755), .B1(new_n250), .B2(new_n833), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1150), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT119), .B1(new_n1149), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT119), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1170), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1142), .B1(new_n1171), .B2(new_n1174), .ZN(G378));
  INV_X1    g0975(.A(G330), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n826), .B1(new_n915), .B2(new_n868), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n892), .A3(new_n919), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1178), .B2(new_n924), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n261), .A2(new_n866), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT55), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n292), .A2(new_n297), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n292), .B2(new_n297), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1181), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1187), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n926), .A2(new_n1179), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n926), .B2(new_n1179), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n907), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n923), .A2(new_n925), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT102), .B1(new_n1177), .B2(new_n919), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n928), .B(G330), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1191), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n893), .A2(new_n906), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n926), .A2(new_n1179), .A3(new_n1192), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1195), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n751), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n833), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n752), .B1(new_n1205), .B2(G50), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G33), .A2(G41), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT120), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n421), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n276), .B2(new_n836), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n840), .A2(new_n545), .B1(new_n785), .B2(G107), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n848), .B2(new_n777), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1212), .A2(G41), .A3(new_n762), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n956), .A2(G77), .B1(new_n792), .B2(G58), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n789), .A2(G97), .B1(new_n797), .B2(G116), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1213), .A2(new_n948), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n786), .A2(new_n1219), .B1(new_n782), .B2(new_n842), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G132), .B2(new_n789), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n797), .A2(G125), .B1(new_n956), .B2(new_n1157), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n245), .C2(new_n804), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1208), .B1(G124), .B2(new_n778), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n807), .C2(new_n791), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1218), .B1(new_n1217), .B2(new_n1216), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1206), .B1(new_n1228), .B2(new_n759), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1191), .B2(new_n757), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1204), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1131), .B1(new_n1138), .B2(new_n1129), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1195), .A2(new_n1202), .A3(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT122), .A4(new_n1201), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(KEYINPUT57), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n694), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1135), .A2(new_n1136), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1129), .B(new_n1114), .C1(new_n1238), .C2(new_n1124), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1132), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1203), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1231), .B1(new_n1237), .B2(new_n1241), .ZN(G375));
  INV_X1    g1042(.A(new_n1140), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1139), .A2(new_n1131), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n993), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n872), .A2(new_n756), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n795), .A2(new_n480), .B1(new_n777), .B2(new_n794), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT123), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1049), .A2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n942), .B1(new_n798), .B2(new_n588), .C1(new_n474), .C2(new_n814), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n313), .B1(new_n384), .B2(new_n782), .C1(new_n786), .C2(new_n848), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n804), .A2(new_n421), .B1(new_n245), .B2(new_n782), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT124), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n797), .A2(G132), .B1(new_n792), .B2(G58), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n807), .B2(new_n795), .C1(new_n814), .C2(new_n1156), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n786), .A2(new_n842), .B1(new_n777), .B2(new_n1219), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n836), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1254), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n752), .B1(G68), .B2(new_n1205), .C1(new_n1261), .C2(new_n835), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT125), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1246), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1139), .B2(new_n750), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1245), .A2(new_n1266), .ZN(G381));
  AND3_X1   g1067(.A1(new_n1134), .A2(new_n1141), .A3(new_n694), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1144), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT117), .B1(new_n1110), .B2(new_n1147), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1170), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1172), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1170), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1268), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1063), .A2(new_n1087), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n986), .A2(new_n988), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1088), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(G375), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1015), .B2(new_n1018), .ZN(G407));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  AOI211_X1 g1082(.A(G375), .B(new_n1279), .C1(new_n1014), .C2(new_n1017), .ZN(new_n1283));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n1274), .A3(new_n674), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(G213), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(G407), .A2(KEYINPUT126), .A3(G213), .A4(new_n1285), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G409));
  NAND3_X1  g1089(.A1(new_n1234), .A2(new_n751), .A3(new_n1235), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1290), .A2(new_n1230), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1240), .A2(new_n993), .A3(new_n1203), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1293), .B(new_n1142), .C1(new_n1171), .C2(new_n1174), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1274), .B2(G375), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n674), .A2(G213), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(new_n694), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT60), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1244), .B1(new_n1140), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1301), .B2(new_n1266), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n855), .B(new_n1265), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1295), .A2(new_n1296), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1266), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n855), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1301), .A2(G384), .A3(new_n1266), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1313), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n821), .B1(new_n1022), .B2(new_n1058), .ZN(new_n1319));
  AOI211_X1 g1119(.A(G396), .B(new_n1057), .C1(new_n985), .C2(new_n1021), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G390), .A2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT109), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1277), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1012), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1325), .B(new_n964), .C1(new_n998), .C2(new_n1011), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1318), .A2(new_n1329), .A3(KEYINPUT61), .ZN(new_n1330));
  OR2_X1    g1130(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1305), .A2(KEYINPUT127), .A3(new_n1306), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1309), .A2(new_n1330), .A3(new_n1331), .A4(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1305), .A2(KEYINPUT62), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1317), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1295), .A2(new_n1304), .A3(new_n1339), .A4(new_n1296), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1334), .A2(new_n1337), .A3(new_n1338), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1329), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1333), .A2(new_n1342), .ZN(G405));
  XNOR2_X1  g1143(.A(G378), .B(G375), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1304), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1347));
  OR3_X1    g1147(.A1(new_n1346), .A2(new_n1347), .A3(new_n1329), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1329), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(G402));
endmodule


