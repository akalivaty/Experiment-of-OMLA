//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n190));
  OR2_X1    g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT2), .B(G113), .Z(new_n192));
  XOR2_X1   g006(.A(new_n191), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G134), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n195), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(new_n196), .ZN(new_n206));
  INV_X1    g020(.A(new_n197), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT67), .A3(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n211), .A2(new_n202), .A3(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n203), .A2(new_n205), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n217), .A3(new_n211), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n200), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G143), .B2(new_n220), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n224), .B(KEYINPUT68), .C1(new_n227), .C2(new_n226), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n221), .A2(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n225), .A3(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n210), .A2(new_n219), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT0), .B(G128), .Z(new_n238));
  OAI211_X1 g052(.A(new_n237), .B(KEYINPUT64), .C1(new_n232), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n213), .A2(new_n216), .A3(new_n218), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n242), .B2(new_n219), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n237), .B1(new_n232), .B2(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n245), .A2(KEYINPUT64), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n235), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n194), .B1(new_n247), .B2(KEYINPUT30), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n206), .A2(new_n217), .A3(new_n211), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n217), .B1(new_n206), .B2(new_n211), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n200), .B1(new_n251), .B2(new_n216), .ZN(new_n252));
  INV_X1    g066(.A(new_n219), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n210), .A2(new_n219), .A3(new_n234), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n210), .A2(new_n219), .A3(new_n234), .A4(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT30), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n242), .A2(new_n219), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n262), .A2(new_n244), .B1(new_n255), .B2(KEYINPUT70), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n263), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n258), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n248), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  AND4_X1   g079(.A1(new_n193), .A2(new_n254), .A3(new_n256), .A4(new_n258), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n267), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n271), .B(new_n272), .Z(new_n273));
  NOR3_X1   g087(.A1(new_n265), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n273), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n262), .A2(new_n246), .A3(new_n239), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n193), .B1(new_n276), .B2(new_n255), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT28), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n235), .B1(new_n244), .B2(new_n262), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT28), .B1(new_n279), .B2(new_n193), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n275), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n188), .B1(new_n274), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n194), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n263), .A2(new_n193), .A3(new_n258), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n280), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n275), .A2(new_n188), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n187), .B1(new_n283), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n287), .A2(new_n273), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n261), .A2(new_n264), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n276), .A2(new_n255), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT30), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n193), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n278), .A2(new_n281), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n275), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT31), .B1(new_n265), .B2(new_n296), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n293), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n297), .A2(new_n300), .ZN(new_n309));
  INV_X1    g123(.A(new_n296), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n275), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n305), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n294), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n292), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  OR3_X1    g134(.A1(new_n320), .A2(KEYINPUT16), .A3(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n220), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(G146), .A3(new_n321), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G110), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n227), .A2(G119), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n331), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT24), .B(G110), .ZN(new_n335));
  OAI221_X1 g149(.A(new_n325), .B1(new_n326), .B2(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n318), .A2(new_n220), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n326), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n335), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n196), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G902), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(KEYINPUT76), .Z(new_n352));
  OAI211_X1 g166(.A(new_n350), .B(new_n351), .C1(new_n345), .C2(new_n352), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n353), .B(KEYINPUT25), .Z(new_n354));
  INV_X1    g168(.A(G217), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(G234), .B2(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n350), .B1(new_n345), .B2(new_n352), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n357), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n317), .A2(KEYINPUT77), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G122), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT84), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G107), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n367), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n371), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(G101), .C1(new_n372), .C2(new_n376), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n381), .A2(new_n194), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n189), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n330), .A2(G116), .ZN(new_n387));
  OAI21_X1  g201(.A(G113), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n192), .A2(new_n189), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  INV_X1    g206(.A(new_n369), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n374), .B(KEYINPUT79), .ZN(new_n395));
  OAI21_X1  g209(.A(G101), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n380), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n380), .A2(new_n392), .A3(new_n396), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n366), .B1(new_n384), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n391), .ZN(new_n402));
  INV_X1    g216(.A(new_n399), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n397), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n381), .A2(new_n194), .A3(new_n383), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n365), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n234), .A2(new_n320), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n320), .B2(new_n245), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n269), .A2(G224), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n412), .B(new_n366), .C1(new_n384), .C2(new_n400), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n409), .B1(KEYINPUT7), .B2(new_n410), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n365), .B(KEYINPUT8), .Z(new_n416));
  AND2_X1   g230(.A1(new_n380), .A2(new_n396), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT85), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n390), .B1(new_n419), .B2(new_n388), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n416), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n380), .A2(new_n396), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n402), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n415), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n410), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n406), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n414), .A2(new_n351), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G210), .B1(G237), .B2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT86), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G214), .B1(G237), .B2(G902), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n414), .A2(new_n351), .A3(new_n429), .A4(new_n426), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n269), .A2(G952), .ZN(new_n435));
  INV_X1    g249(.A(G234), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(new_n268), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n351), .B(new_n269), .C1(G234), .C2(G237), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT21), .B(G898), .Z(new_n440));
  OAI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n417), .A2(new_n234), .ZN(new_n444));
  INV_X1    g258(.A(new_n233), .ZN(new_n445));
  INV_X1    g259(.A(new_n226), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n227), .B1(new_n446), .B2(KEYINPUT80), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(KEYINPUT80), .B2(new_n446), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n448), .B2(new_n224), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n422), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n262), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT12), .ZN(new_n452));
  OAI211_X1 g266(.A(KEYINPUT10), .B(new_n234), .C1(new_n403), .C2(new_n397), .ZN(new_n453));
  INV_X1    g267(.A(new_n262), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n381), .A2(new_n244), .A3(new_n383), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n449), .B2(new_n422), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G140), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n269), .A2(G227), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n459), .B(new_n460), .Z(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n262), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n465), .B2(new_n458), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n443), .B(new_n351), .C1(new_n463), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n443), .A2(new_n351), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n461), .ZN(new_n470));
  INV_X1    g284(.A(new_n458), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n452), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n458), .A3(new_n461), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n467), .B(new_n469), .C1(new_n474), .C2(new_n443), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT9), .B(G234), .Z(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G221), .B1(new_n477), .B2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G475), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT90), .B(G104), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n318), .B(KEYINPUT19), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n220), .ZN(new_n486));
  INV_X1    g300(.A(new_n338), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT89), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n222), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G131), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(G143), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n200), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n339), .A2(new_n497), .A3(new_n486), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n318), .A2(new_n220), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT87), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n340), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n340), .B2(new_n500), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n493), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT18), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n495), .B(KEYINPUT88), .C1(KEYINPUT18), .C2(new_n492), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n494), .B(new_n508), .C1(new_n509), .C2(new_n200), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n484), .B1(new_n499), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n325), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n505), .A2(KEYINPUT17), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n514), .C1(KEYINPUT17), .C2(new_n496), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n511), .A3(new_n484), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n480), .B(new_n351), .C1(new_n512), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n519));
  AND4_X1   g333(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n337), .A2(new_n338), .B1(new_n220), .B2(new_n485), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n521), .A2(new_n497), .B1(new_n493), .B2(new_n495), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n522), .B2(new_n490), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n523), .B2(new_n484), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n480), .A4(new_n351), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n526), .A3(KEYINPUT20), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n484), .B1(new_n515), .B2(new_n511), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n351), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT92), .B(G475), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n518), .A2(KEYINPUT91), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n477), .A2(new_n355), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n227), .B2(G143), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n222), .A2(KEYINPUT94), .A3(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT13), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n227), .A2(G143), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n541), .B2(new_n542), .ZN(new_n546));
  OAI21_X1  g360(.A(G134), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n541), .A2(new_n545), .A3(new_n215), .ZN(new_n548));
  INV_X1    g362(.A(G116), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT93), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n549), .A2(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n369), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n393), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n547), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n551), .A2(KEYINPUT14), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n552), .B1(new_n551), .B2(KEYINPUT14), .ZN(new_n559));
  OAI21_X1  g373(.A(G107), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n548), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n215), .B1(new_n541), .B2(new_n545), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n560), .B(new_n555), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n537), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n557), .A2(new_n563), .A3(new_n537), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n536), .B1(new_n568), .B2(G902), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n567), .B(new_n351), .C1(KEYINPUT15), .C2(new_n535), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(KEYINPUT96), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT96), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR4_X1   g387(.A1(new_n442), .A2(new_n479), .A3(new_n534), .A4(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n316), .B2(new_n361), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n363), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  AOI21_X1  g392(.A(new_n187), .B1(new_n313), .B2(new_n351), .ZN(new_n579));
  NOR4_X1   g393(.A1(new_n479), .A2(new_n361), .A3(new_n306), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n565), .A2(KEYINPUT97), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n567), .A2(new_n581), .A3(KEYINPUT33), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n565), .B(new_n566), .C1(KEYINPUT97), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(G478), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n567), .A2(new_n535), .A3(new_n351), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n535), .A2(new_n351), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n534), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n442), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT34), .B(G104), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  INV_X1    g408(.A(new_n573), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n442), .A2(new_n534), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n580), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT98), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT35), .B(G107), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  NOR2_X1   g414(.A1(new_n579), .A2(new_n306), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n352), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n345), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n345), .A2(new_n602), .A3(new_n352), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n359), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT99), .Z(new_n608));
  NAND2_X1  g422(.A1(new_n357), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n574), .A2(new_n601), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G110), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n610), .B(new_n612), .ZN(G12));
  INV_X1    g427(.A(new_n434), .ZN(new_n614));
  INV_X1    g428(.A(new_n609), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n316), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n479), .ZN(new_n617));
  INV_X1    g431(.A(new_n437), .ZN(new_n618));
  INV_X1    g432(.A(G900), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n438), .B2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n595), .A2(new_n534), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  INV_X1    g437(.A(new_n534), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n595), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n620), .B(KEYINPUT39), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n617), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n625), .B1(new_n628), .B2(KEYINPUT40), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n431), .A2(new_n433), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT38), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n629), .A2(new_n609), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n308), .A2(new_n315), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n265), .A2(new_n266), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n275), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n286), .A2(new_n287), .A3(new_n275), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n351), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n628), .A2(KEYINPUT40), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n632), .A2(new_n432), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G143), .ZN(G45));
  INV_X1    g456(.A(new_n620), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n589), .A2(new_n534), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n616), .A2(new_n617), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G146), .ZN(G48));
  NOR2_X1   g460(.A1(new_n316), .A2(new_n361), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n351), .B1(new_n463), .B2(new_n466), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G469), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n478), .A3(new_n467), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n647), .A2(new_n591), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  NAND3_X1  g467(.A1(new_n647), .A2(new_n596), .A3(new_n650), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G116), .ZN(G18));
  NOR2_X1   g469(.A1(new_n316), .A2(new_n615), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n442), .A2(new_n534), .A3(new_n573), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n650), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT101), .B(G119), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G21));
  OAI21_X1  g474(.A(new_n275), .B1(new_n288), .B2(new_n280), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n305), .A2(new_n311), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n294), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(KEYINPUT102), .A3(new_n294), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n579), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n362), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT103), .B1(new_n595), .B2(new_n624), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n573), .A2(new_n671), .A3(new_n534), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n442), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n650), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G122), .ZN(G24));
  NAND2_X1  g489(.A1(new_n313), .A2(new_n351), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n662), .A2(KEYINPUT102), .A3(new_n294), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n662), .B2(new_n294), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n677), .B(new_n609), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n665), .A2(new_n666), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n677), .A4(new_n609), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n644), .A2(new_n650), .A3(new_n434), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT105), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n681), .A2(new_n684), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n689));
  INV_X1    g503(.A(new_n686), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  NAND2_X1  g507(.A1(new_n314), .A2(new_n293), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n292), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n314), .B2(new_n293), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n306), .A2(new_n699), .A3(KEYINPUT32), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n362), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n630), .A2(new_n432), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n630), .A2(KEYINPUT106), .A3(new_n432), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n617), .A2(new_n705), .A3(new_n644), .A4(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT42), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n479), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n647), .A3(new_n711), .A4(new_n644), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n200), .ZN(G33));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n647), .A3(new_n621), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G134), .ZN(G36));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n717), .B1(new_n474), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n443), .B1(new_n474), .B2(new_n718), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n472), .A2(KEYINPUT109), .A3(KEYINPUT45), .A4(new_n473), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n469), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n467), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT46), .B1(new_n722), .B2(new_n469), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n478), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n726), .A2(new_n626), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n534), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT43), .B1(new_n534), .B2(new_n729), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n601), .A3(new_n615), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n709), .B1(new_n735), .B2(KEYINPUT44), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n728), .B(new_n736), .C1(KEYINPUT44), .C2(new_n735), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(KEYINPUT47), .B(new_n478), .C1(new_n724), .C2(new_n725), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n709), .A2(new_n590), .A3(new_n620), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n316), .A3(new_n361), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  NAND2_X1  g559(.A1(new_n649), .A2(new_n467), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT49), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n478), .A2(new_n631), .A3(new_n730), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n639), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n361), .B1(new_n746), .B2(KEYINPUT49), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n432), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n752));
  INV_X1    g566(.A(new_n478), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n709), .A2(new_n753), .A3(new_n746), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n361), .A2(new_n437), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n534), .A3(new_n589), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n754), .A2(new_n618), .A3(new_n733), .A4(new_n732), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(new_n685), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n732), .A2(new_n618), .A3(new_n733), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n668), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n432), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n631), .A4(new_n650), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n758), .B(new_n760), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n649), .A2(new_n753), .A3(new_n467), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n740), .A2(new_n741), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n668), .A2(new_n761), .A3(new_n709), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n752), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n768), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n757), .B1(new_n775), .B2(new_n766), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n740), .A2(KEYINPUT115), .A3(new_n741), .A4(new_n770), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n776), .A2(new_n780), .A3(KEYINPUT51), .A4(new_n760), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n774), .A2(new_n781), .A3(new_n435), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n756), .A2(new_n590), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n759), .B1(KEYINPUT116), .B2(KEYINPUT48), .ZN(new_n784));
  INV_X1    g598(.A(new_n702), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n786), .B(new_n787), .Z(new_n788));
  NAND3_X1  g602(.A1(new_n762), .A2(new_n434), .A3(new_n650), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n782), .A2(new_n783), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n616), .B(new_n617), .C1(new_n621), .C2(new_n644), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n614), .B1(new_n670), .B2(new_n672), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n620), .A2(KEYINPUT111), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n620), .A2(KEYINPUT111), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n479), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n615), .A3(new_n639), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n692), .A2(new_n791), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n799));
  AOI211_X1 g613(.A(KEYINPUT105), .B(new_n686), .C1(new_n681), .C2(new_n684), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n792), .B(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n569), .A2(new_n570), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n534), .A2(new_n803), .A3(new_n620), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n705), .A2(new_n706), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n705), .A2(KEYINPUT110), .A3(new_n706), .A4(new_n804), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n656), .A3(new_n617), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n803), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n590), .B1(new_n534), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n580), .A2(new_n434), .A3(new_n441), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n577), .A2(new_n809), .A3(new_n610), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n715), .B1(new_n685), .B2(new_n707), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n674), .A2(new_n651), .A3(new_n654), .A4(new_n658), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n713), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n798), .A2(new_n802), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n820));
  OAI211_X1 g634(.A(new_n819), .B(KEYINPUT54), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n801), .B(new_n791), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n817), .B2(KEYINPUT113), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n713), .B2(new_n816), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n822), .A2(new_n815), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  INV_X1    g642(.A(new_n820), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n818), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n821), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n790), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(G952), .A2(G953), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n751), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(KEYINPUT117), .B(new_n751), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(G75));
  AOI21_X1  g656(.A(new_n351), .B1(new_n827), .B2(new_n830), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(new_n429), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n407), .A2(new_n413), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(new_n411), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT55), .Z(new_n848));
  AND2_X1   g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n845), .A2(new_n848), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n269), .A2(G952), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G51));
  NAND2_X1  g666(.A1(new_n827), .A2(new_n830), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n831), .ZN(new_n855));
  XOR2_X1   g669(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n468), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n468), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(new_n466), .B2(new_n463), .ZN(new_n859));
  INV_X1    g673(.A(new_n722), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n843), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n851), .B1(new_n859), .B2(new_n861), .ZN(G54));
  NAND4_X1  g676(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n863));
  INV_X1    g677(.A(new_n524), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n851), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n863), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n863), .B2(new_n864), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n866), .B(KEYINPUT120), .C1(new_n869), .C2(new_n868), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(G60));
  XNOR2_X1  g688(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n588), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n582), .A2(new_n584), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT121), .Z(new_n878));
  AOI211_X1 g692(.A(new_n876), .B(new_n878), .C1(new_n854), .C2(new_n831), .ZN(new_n879));
  INV_X1    g693(.A(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n833), .A2(new_n835), .A3(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n851), .B(new_n879), .C1(new_n881), .C2(new_n878), .ZN(G63));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n883));
  NAND2_X1  g697(.A1(G217), .A2(G902), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT60), .Z(new_n885));
  NAND3_X1  g699(.A1(new_n853), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n853), .B2(new_n885), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n606), .B(new_n605), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n851), .ZN(new_n890));
  INV_X1    g704(.A(new_n888), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n358), .A3(new_n886), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n889), .A2(new_n892), .A3(KEYINPUT61), .A4(new_n890), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(G66));
  NAND2_X1  g711(.A1(new_n440), .A2(G224), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(G953), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n577), .A2(new_n610), .A3(new_n812), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n816), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n901), .B2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n846), .B1(G898), .B2(new_n269), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(G69));
  OAI21_X1  g718(.A(new_n297), .B1(KEYINPUT30), .B2(new_n247), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(new_n485), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n363), .A2(new_n576), .A3(new_n627), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n710), .A2(new_n811), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n692), .A2(new_n792), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(KEYINPUT62), .A3(new_n641), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n641), .A2(new_n692), .A3(new_n792), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n737), .A2(new_n744), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT124), .B(new_n907), .C1(new_n918), .C2(G953), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  AOI21_X1  g735(.A(G953), .B1(new_n916), .B2(new_n917), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n906), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(G227), .A2(G900), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(G953), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(G900), .A2(G953), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n728), .A2(new_n785), .A3(new_n793), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n708), .A2(new_n712), .A3(new_n715), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n917), .A2(new_n911), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n906), .B(new_n927), .C1(new_n930), .C2(G953), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n919), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n926), .B(new_n932), .ZN(G72));
  XNOR2_X1  g747(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n187), .A2(new_n351), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(new_n936));
  INV_X1    g750(.A(new_n901), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n274), .B(KEYINPUT127), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n851), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n936), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n918), .B2(new_n901), .ZN(new_n942));
  INV_X1    g756(.A(new_n635), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n819), .B1(new_n818), .B2(new_n820), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n945), .A2(new_n274), .A3(new_n635), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n936), .B2(new_n946), .ZN(G57));
endmodule


