//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G250), .B1(G257), .B2(G264), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n215), .A2(KEYINPUT0), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n222), .B(new_n230), .C1(KEYINPUT0), .C2(new_n215), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G116), .Z(new_n240));
  NAND2_X1  g0040(.A1(G97), .A2(G107), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n209), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n240), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n201), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n251), .A2(new_n253), .A3(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n253), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n254), .A2(G223), .B1(G77), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G222), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n251), .B(new_n253), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n262), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n265), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n267), .B1(new_n270), .B2(G226), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n216), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n205), .A2(G20), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT8), .B(G58), .Z(new_n278));
  NAND2_X1  g0078(.A1(new_n217), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n217), .A2(new_n250), .A3(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G20), .B2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n278), .A2(new_n280), .B1(new_n284), .B2(G150), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n276), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n201), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n276), .B1(G1), .B2(new_n217), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n201), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n273), .A2(G190), .B1(KEYINPUT9), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n272), .A2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n293), .A2(new_n300), .A3(new_n294), .A4(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n254), .A2(G238), .B1(G107), .B2(new_n255), .ZN(new_n303));
  INV_X1    g0103(.A(G232), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n260), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n262), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n267), .B1(new_n270), .B2(G244), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT68), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT15), .B(G87), .Z(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n278), .A2(new_n284), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n276), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G77), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n288), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n290), .B2(new_n316), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n308), .B2(G200), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n292), .B1(new_n272), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G179), .B2(new_n272), .ZN(new_n324));
  INV_X1    g0124(.A(new_n308), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n319), .B1(new_n325), .B2(G169), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AND4_X1   g0130(.A1(new_n302), .A2(new_n321), .A3(new_n324), .A4(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  INV_X1    g0133(.A(G226), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n260), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT3), .B(G33), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT66), .B(G1698), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT69), .A4(G226), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n251), .A2(new_n253), .A3(G232), .A4(G1698), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n335), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n262), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n268), .A2(G238), .A3(new_n265), .ZN(new_n343));
  INV_X1    g0143(.A(new_n267), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n332), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  AOI211_X1 g0147(.A(KEYINPUT13), .B(new_n345), .C1(new_n341), .C2(new_n262), .ZN(new_n348));
  OAI21_X1  g0148(.A(G200), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n340), .A2(new_n339), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n336), .A2(new_n337), .A3(G226), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n333), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n268), .B1(new_n352), .B2(new_n338), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT13), .B1(new_n353), .B2(new_n345), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n342), .A2(new_n332), .A3(new_n346), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G190), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n287), .B2(G68), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT12), .Z(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n203), .B2(new_n290), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n281), .A2(new_n283), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n201), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n279), .A2(new_n316), .B1(new_n217), .B2(G68), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n275), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(KEYINPUT11), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(KEYINPUT11), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n360), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n349), .A2(new_n356), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT71), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n349), .A2(new_n356), .A3(new_n370), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n367), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n354), .A2(G179), .A3(new_n355), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n322), .B1(new_n354), .B2(new_n355), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n373), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n331), .A2(new_n372), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n255), .B2(new_n217), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n383), .B(G20), .C1(new_n251), .C2(new_n253), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G159), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n281), .B2(new_n283), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n217), .B1(new_n220), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT72), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n220), .A2(new_n388), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G20), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n361), .C2(new_n386), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n390), .A4(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n383), .B1(new_n336), .B2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n203), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n392), .B1(new_n361), .B2(new_n386), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n275), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n395), .A2(new_n401), .A3(KEYINPUT74), .A4(new_n275), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n278), .A2(new_n288), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n278), .B2(new_n290), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n344), .B1(new_n269), .B2(new_n304), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n251), .A2(new_n253), .A3(G226), .A4(G1698), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  INV_X1    g0213(.A(G223), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(new_n413), .C1(new_n260), .C2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT75), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n268), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n336), .A2(new_n337), .A3(G223), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n418), .A2(KEYINPUT75), .A3(new_n412), .A4(new_n413), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n411), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G179), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n322), .B2(new_n420), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n410), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n408), .B1(new_n404), .B2(new_n405), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n415), .A2(new_n416), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n419), .A3(new_n262), .ZN(new_n427));
  INV_X1    g0227(.A(new_n411), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n322), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(G179), .B2(new_n420), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT76), .B(G190), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n427), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G200), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n427), .B2(new_n428), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n424), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n432), .B1(new_n424), .B2(new_n437), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n423), .A2(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n381), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g0243(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n444));
  OAI21_X1  g0244(.A(G244), .B1(KEYINPUT79), .B2(KEYINPUT4), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n260), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(new_n445), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n336), .A2(new_n337), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(G1698), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n446), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n262), .ZN(new_n453));
  INV_X1    g0253(.A(G41), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n264), .B(G45), .C1(new_n454), .C2(KEYINPUT5), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT80), .B1(new_n454), .B2(KEYINPUT5), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(G274), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT80), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(G41), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n463), .A2(new_n459), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT81), .B1(new_n467), .B2(new_n266), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n262), .B1(new_n457), .B2(new_n459), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n460), .A2(new_n468), .B1(new_n469), .B2(G257), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n453), .A2(new_n470), .A3(G190), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n382), .B2(new_n384), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n208), .A2(G97), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n209), .A3(new_n241), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(G20), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n284), .A2(KEYINPUT77), .A3(G77), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT77), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n361), .B2(new_n316), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n472), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n275), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n287), .A2(G97), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n264), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n287), .A2(new_n486), .A3(new_n216), .A4(new_n274), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(new_n207), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n471), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n435), .B1(new_n453), .B2(new_n470), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n443), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n482), .B2(new_n275), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(KEYINPUT82), .A3(new_n494), .A4(new_n471), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n287), .A2(KEYINPUT25), .A3(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT25), .B1(new_n287), .B2(G107), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n498), .C1(new_n208), .C2(new_n487), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT86), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n487), .A2(new_n208), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT86), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n498), .A4(new_n497), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n217), .A3(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT23), .B1(new_n208), .B2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n506), .A2(new_n507), .B1(G20), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n251), .A2(new_n253), .A3(new_n217), .A4(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT22), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n336), .A2(new_n512), .A3(new_n217), .A4(G87), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n275), .B1(new_n514), .B2(KEYINPUT24), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(new_n509), .C1(new_n511), .C2(new_n513), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n504), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n468), .A2(new_n460), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n469), .A2(G264), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n251), .A2(new_n253), .A3(G257), .A4(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G294), .ZN(new_n523));
  INV_X1    g0323(.A(G250), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n260), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n262), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT87), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT87), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n528), .A3(new_n262), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n521), .A2(new_n527), .A3(new_n309), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n435), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n518), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n465), .B2(G274), .ZN(new_n535));
  NOR4_X1   g0335(.A1(new_n464), .A2(new_n266), .A3(KEYINPUT83), .A4(G1), .ZN(new_n536));
  OAI21_X1  g0336(.A(G250), .B1(new_n464), .B2(G1), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n535), .A2(new_n536), .B1(new_n262), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n336), .A2(G244), .A3(G1698), .ZN(new_n539));
  INV_X1    g0339(.A(G238), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(new_n508), .C1(new_n540), .C2(new_n260), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n262), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n312), .A2(new_n287), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n487), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n336), .A2(new_n217), .A3(G68), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n217), .B1(new_n339), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G87), .B2(new_n209), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n279), .B2(new_n207), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n544), .B(new_n546), .C1(new_n552), .C2(new_n275), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n543), .B(new_n553), .C1(new_n435), .C2(new_n542), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n275), .ZN(new_n555));
  INV_X1    g0355(.A(new_n544), .ZN(new_n556));
  INV_X1    g0356(.A(new_n312), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n487), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n541), .A2(new_n262), .ZN(new_n559));
  INV_X1    g0359(.A(new_n538), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n328), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(new_n561), .C1(G169), .C2(new_n542), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n533), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n483), .A2(new_n489), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n453), .A2(new_n470), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n322), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n453), .A2(new_n470), .A3(new_n328), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n496), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n527), .A2(new_n519), .A3(new_n529), .A4(new_n520), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G169), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT88), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT88), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n574), .A3(G169), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n531), .A2(new_n328), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n518), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n254), .A2(G264), .B1(G303), .B2(new_n255), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT85), .A4(G257), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT85), .ZN(new_n582));
  INV_X1    g0382(.A(G257), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n260), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n262), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n469), .A2(G270), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n519), .A2(new_n587), .A3(KEYINPUT84), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT84), .B1(new_n519), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n450), .B(new_n217), .C1(G33), .C2(new_n207), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n591), .B(new_n275), .C1(new_n217), .C2(G116), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT20), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n288), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n487), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n322), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n590), .A2(new_n598), .A3(KEYINPUT21), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT21), .B1(new_n590), .B2(new_n598), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n519), .A2(new_n587), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n519), .A2(new_n587), .A3(KEYINPUT84), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(new_n262), .B2(new_n585), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n433), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(new_n597), .C1(new_n435), .C2(new_n607), .ZN(new_n609));
  INV_X1    g0409(.A(new_n597), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(G179), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n579), .A2(new_n602), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n442), .A2(new_n570), .A3(new_n612), .ZN(G372));
  NAND2_X1  g0413(.A1(new_n590), .A2(new_n598), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n611), .A3(new_n599), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT89), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n616), .A2(KEYINPUT89), .A3(new_n611), .A4(new_n599), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n579), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n496), .A2(new_n564), .A3(new_n569), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n563), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT26), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n563), .A2(new_n569), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n562), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT90), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT26), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n563), .B2(new_n569), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(new_n562), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n441), .B1(new_n623), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT91), .Z(new_n638));
  NAND3_X1  g0438(.A1(new_n372), .A2(new_n329), .A3(new_n327), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n380), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n406), .A2(new_n409), .A3(new_n437), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n424), .A2(new_n432), .A3(new_n437), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n425), .B1(new_n424), .B2(new_n430), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n410), .A2(KEYINPUT18), .A3(new_n422), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n640), .A2(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n302), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n324), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n638), .A2(new_n649), .ZN(G369));
  INV_X1    g0450(.A(new_n518), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n576), .B1(new_n572), .B2(KEYINPUT88), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n575), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n217), .A2(G13), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n264), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT92), .B1(new_n518), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  INV_X1    g0462(.A(new_n660), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n651), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  OR4_X1    g0464(.A1(new_n533), .A2(new_n653), .A3(new_n661), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n617), .A2(new_n663), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n653), .B2(new_n663), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n663), .A2(new_n597), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n619), .A2(new_n620), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n617), .B1(new_n597), .B2(new_n663), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n609), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n665), .B1(new_n579), .B2(new_n663), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT93), .ZN(G399));
  NOR2_X1   g0478(.A1(new_n213), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n221), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g0483(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n684));
  XNOR2_X1  g0484(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n636), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n621), .A2(new_n622), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n660), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n562), .B(KEYINPUT96), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n617), .A2(new_n653), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n633), .B(new_n691), .C1(new_n692), .C2(new_n570), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n663), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(new_n689), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n542), .A2(new_n526), .A3(new_n520), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n566), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n607), .A2(new_n699), .A3(G179), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n607), .A2(new_n699), .A3(KEYINPUT30), .A4(G179), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n542), .A2(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n590), .A2(new_n566), .A3(new_n531), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n660), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n612), .A2(new_n570), .A3(new_n660), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n706), .B2(new_n660), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n708), .B(G330), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n708), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n622), .A2(new_n692), .A3(new_n609), .A4(new_n663), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n710), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT95), .A3(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n697), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n685), .B1(new_n722), .B2(G1), .ZN(G364));
  NAND3_X1  g0523(.A1(new_n328), .A2(new_n435), .A3(G190), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G97), .ZN(new_n726));
  NOR4_X1   g0526(.A1(new_n217), .A2(new_n309), .A3(new_n435), .A4(G179), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n336), .B(new_n726), .C1(new_n728), .C2(new_n545), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n309), .A2(G20), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT102), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n732), .A2(G179), .A3(new_n435), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n208), .ZN(new_n735));
  NAND2_X1  g0535(.A1(G20), .A2(G179), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT100), .Z(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G200), .A3(new_n433), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n729), .B(new_n735), .C1(G50), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n309), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n435), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n740), .B1(new_n203), .B2(new_n743), .C1(new_n316), .C2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n732), .A2(G179), .A3(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G159), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT32), .Z(new_n749));
  NAND3_X1  g0549(.A1(new_n737), .A2(new_n435), .A3(new_n433), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT101), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n202), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G322), .B1(new_n733), .B2(G283), .ZN(new_n755));
  INV_X1    g0555(.A(G329), .ZN(new_n756));
  INV_X1    g0556(.A(new_n747), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n725), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n255), .B1(new_n759), .B2(new_n760), .C1(new_n728), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(G326), .B2(new_n739), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  OAI221_X1 g0565(.A(new_n763), .B1(new_n764), .B2(new_n745), .C1(new_n743), .C2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n746), .A2(new_n753), .B1(new_n758), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n216), .B1(G20), .B2(new_n322), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n264), .B1(new_n654), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n679), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n213), .A2(new_n594), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n248), .A2(new_n464), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n213), .A2(new_n336), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G45), .B2(new_n221), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n213), .A2(new_n255), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(G355), .B(KEYINPUT98), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n774), .B1(new_n775), .B2(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n768), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n773), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n769), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n672), .B2(new_n785), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n674), .A2(new_n772), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n672), .A2(new_n673), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NOR2_X1   g0595(.A1(new_n330), .A2(new_n660), .ZN(new_n796));
  INV_X1    g0596(.A(new_n319), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n321), .B1(new_n797), .B2(new_n663), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(new_n798), .B2(new_n330), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n784), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n742), .A2(G283), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n733), .A2(G87), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n336), .B1(new_n727), .B2(G107), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n801), .A2(new_n726), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n739), .A2(G303), .B1(new_n747), .B2(G311), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n760), .B2(new_n750), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(G116), .C2(new_n744), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n744), .A2(G159), .B1(new_n739), .B2(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G150), .ZN(new_n809));
  INV_X1    g0609(.A(G143), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n743), .C1(new_n752), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT34), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n336), .B1(new_n728), .B2(new_n201), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G58), .B2(new_n725), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n733), .A2(G68), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n814), .B(new_n815), .C1(new_n816), .C2(new_n757), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT103), .Z(new_n818));
  AOI21_X1  g0618(.A(new_n807), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n768), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n784), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n819), .A2(new_n820), .B1(G77), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n772), .B1(new_n800), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n799), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n715), .B2(new_n720), .ZN(new_n825));
  INV_X1    g0625(.A(new_n688), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n714), .A2(new_n719), .A3(new_n799), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n773), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n826), .B1(new_n825), .B2(new_n827), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT104), .ZN(G384));
  NAND2_X1  g0632(.A1(new_n476), .A2(new_n477), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT35), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n594), .B(new_n219), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT36), .Z(new_n837));
  NAND4_X1  g0637(.A1(new_n220), .A2(G50), .A3(G77), .A4(new_n388), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n264), .B(G13), .C1(new_n838), .C2(new_n244), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n372), .A2(new_n380), .A3(KEYINPUT106), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n367), .A2(new_n663), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n842), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n372), .A2(new_n380), .A3(KEYINPUT106), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n718), .A2(new_n799), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT108), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n410), .A2(new_n422), .ZN(new_n849));
  INV_X1    g0649(.A(new_n658), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n410), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n641), .ZN(new_n853));
  INV_X1    g0653(.A(new_n396), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n385), .A2(new_n394), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n390), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n395), .A2(new_n275), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n409), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n422), .B2(new_n850), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n641), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n645), .A2(new_n646), .B1(new_n642), .B2(new_n643), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n850), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(KEYINPUT38), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n424), .A2(new_n658), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n641), .B1(new_n424), .B2(new_n430), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n867), .B2(new_n866), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n440), .A2(new_n866), .B1(new_n868), .B2(new_n853), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n869), .B2(KEYINPUT38), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT40), .A4(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n853), .A2(new_n861), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n646), .A2(new_n645), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n864), .B1(new_n873), .B2(new_n644), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n440), .A2(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n868), .A2(new_n853), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n718), .A2(new_n846), .A3(KEYINPUT40), .A4(new_n799), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT108), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  INV_X1    g0683(.A(new_n864), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n440), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n885), .B2(new_n862), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n718), .A2(new_n846), .A3(new_n799), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n871), .A2(new_n882), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT109), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n441), .A2(new_n718), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n673), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n891), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n442), .B1(new_n690), .B2(new_n695), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n649), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  NOR2_X1   g0698(.A1(new_n380), .A2(new_n660), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n865), .B(new_n900), .C1(new_n869), .C2(KEYINPUT38), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n875), .B1(new_n872), .B2(new_n874), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n900), .B1(new_n903), .B2(new_n865), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n899), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n663), .B(new_n799), .C1(new_n623), .C2(new_n636), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n796), .B(KEYINPUT105), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n865), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n846), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n873), .A2(new_n850), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n905), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n898), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n264), .B2(new_n654), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n898), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n840), .B1(new_n917), .B2(new_n918), .ZN(G367));
  OAI22_X1  g0719(.A1(new_n750), .A2(new_n809), .B1(new_n203), .B2(new_n759), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT114), .Z(new_n921));
  OAI221_X1 g0721(.A(new_n336), .B1(new_n738), .B2(new_n810), .C1(new_n734), .C2(new_n316), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n201), .A2(new_n745), .B1(new_n743), .B2(new_n386), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(KEYINPUT115), .B(G137), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n747), .A2(new_n925), .B1(G58), .B2(new_n727), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT116), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n727), .A2(G116), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT46), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n208), .B2(new_n759), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(G311), .B2(new_n739), .ZN(new_n931));
  AOI22_X1  g0731(.A1(G283), .A2(new_n744), .B1(new_n742), .B2(G294), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n761), .C2(new_n752), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n733), .A2(G97), .ZN(new_n934));
  INV_X1    g0734(.A(G317), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n255), .C1(new_n757), .C2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT113), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n924), .A2(new_n927), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT47), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n820), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n663), .A2(new_n553), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n624), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n562), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n785), .ZN(new_n947));
  INV_X1    g0747(.A(new_n776), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n238), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n786), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n213), .B2(new_n312), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n773), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n941), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n496), .B(new_n569), .C1(new_n494), .C2(new_n663), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT110), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n625), .A2(new_n660), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n668), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT45), .Z(new_n959));
  NOR2_X1   g0759(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n668), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n668), .B2(new_n957), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n676), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n959), .A2(new_n964), .A3(new_n676), .ZN(new_n967));
  INV_X1    g0767(.A(new_n667), .ZN(new_n968));
  INV_X1    g0768(.A(new_n666), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n675), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n674), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n966), .A2(new_n722), .A3(new_n967), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n722), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n974));
  XNOR2_X1  g0774(.A(new_n679), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n771), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n957), .A2(new_n667), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n569), .B1(new_n955), .B2(new_n579), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n977), .A2(KEYINPUT42), .B1(new_n979), .B2(new_n663), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n946), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n978), .A2(new_n980), .A3(new_n982), .A4(new_n946), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n957), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n676), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n987), .B(new_n989), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n953), .B1(new_n976), .B2(new_n990), .ZN(G387));
  OAI21_X1  g0791(.A(new_n776), .B1(new_n235), .B2(new_n464), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n681), .B2(new_n780), .ZN(new_n993));
  INV_X1    g0793(.A(new_n278), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n994), .A2(KEYINPUT50), .A3(G50), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT50), .B1(new_n994), .B2(G50), .ZN(new_n996));
  AOI21_X1  g0796(.A(G45), .B1(G68), .B2(G77), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n995), .A2(new_n681), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n993), .A2(new_n998), .B1(new_n208), .B2(new_n213), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n772), .B1(new_n999), .B2(new_n950), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n255), .B1(new_n727), .B2(G77), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n934), .B(new_n1001), .C1(new_n757), .C2(new_n809), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT117), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n312), .A2(new_n725), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n738), .B2(new_n386), .C1(new_n201), .C2(new_n750), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n203), .A2(new_n745), .B1(new_n743), .B2(new_n994), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n336), .B1(new_n747), .B2(G326), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n744), .A2(G303), .B1(new_n739), .B2(G322), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n764), .B2(new_n743), .C1(new_n752), .C2(new_n935), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT48), .Z(new_n1011));
  INV_X1    g0811(.A(G283), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n728), .A2(new_n760), .B1(new_n759), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1008), .B1(new_n594), .B2(new_n734), .C1(new_n1014), .C2(KEYINPUT49), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1014), .A2(KEYINPUT49), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1000), .B1(new_n1017), .B2(new_n768), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n665), .B(new_n785), .C1(new_n579), .C2(new_n663), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n971), .A2(new_n771), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n722), .A2(new_n971), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n679), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n722), .A2(new_n971), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G393));
  INV_X1    g0824(.A(new_n967), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n1025), .B2(new_n965), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n972), .A2(new_n1026), .A3(new_n679), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n966), .A2(new_n771), .A3(new_n967), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n988), .A2(new_n785), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n255), .B1(new_n759), .B2(new_n594), .C1(new_n728), .C2(new_n1012), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1030), .B(new_n735), .C1(G322), .C2(new_n747), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G294), .A2(new_n744), .B1(new_n742), .B2(G303), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n764), .A2(new_n750), .B1(new_n738), .B2(new_n935), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT52), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n725), .A2(G77), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n743), .B2(new_n201), .C1(new_n994), .C2(new_n745), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT118), .Z(new_n1038));
  OAI22_X1  g0838(.A1(new_n809), .A2(new_n738), .B1(new_n750), .B2(new_n386), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n747), .A2(G143), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n255), .B1(new_n727), .B2(G68), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1040), .A2(new_n802), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n768), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n786), .B1(new_n207), .B2(new_n212), .C1(new_n243), .C2(new_n948), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1029), .A2(new_n772), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1027), .A2(new_n1028), .A3(new_n1047), .ZN(G390));
  AOI21_X1  g0848(.A(new_n907), .B1(new_n694), .B2(new_n799), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n846), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n870), .B1(new_n380), .B2(new_n660), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n899), .B1(new_n909), .B2(new_n846), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n901), .B1(new_n887), .B2(new_n900), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n712), .A2(new_n1050), .A3(new_n824), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1050), .A2(new_n824), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n714), .A3(new_n719), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1051), .B(new_n1058), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n771), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n772), .B1(new_n821), .B2(new_n278), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n757), .A2(new_n760), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n815), .A2(new_n1036), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n336), .B1(new_n727), .B2(G87), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1062), .B(new_n1063), .C1(KEYINPUT121), .C2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n738), .A2(new_n1012), .B1(new_n1064), .B2(KEYINPUT121), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G116), .B2(new_n754), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G97), .A2(new_n744), .B1(new_n742), .B2(G107), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G128), .A2(new_n739), .B1(new_n754), .B2(G132), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT120), .Z(new_n1071));
  XOR2_X1   g0871(.A(KEYINPUT54), .B(G143), .Z(new_n1072));
  AOI22_X1  g0872(.A1(new_n742), .A2(new_n925), .B1(new_n744), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(KEYINPUT119), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n728), .A2(new_n809), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT53), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1075), .A2(new_n1076), .B1(new_n386), .B2(new_n759), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n255), .B(new_n1077), .C1(new_n1076), .C2(new_n1075), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1073), .A2(KEYINPUT119), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G50), .A2(new_n733), .B1(new_n747), .B2(G125), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1069), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1061), .B1(new_n1082), .B2(new_n768), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1053), .B2(new_n784), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1060), .A2(KEYINPUT122), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT122), .B1(new_n1060), .B2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1050), .B1(new_n712), .B2(new_n824), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1058), .A2(new_n1049), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1055), .B1(new_n827), .B2(new_n1050), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n909), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n892), .A2(new_n673), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n896), .A2(new_n1092), .A3(new_n649), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1056), .A2(new_n1059), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1056), .A2(new_n1091), .A3(new_n1093), .A4(new_n1059), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n679), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1085), .A2(new_n1086), .B1(new_n1094), .B2(new_n1096), .ZN(G378));
  INV_X1    g0897(.A(KEYINPUT125), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n890), .A2(new_n914), .A3(G330), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n871), .A2(new_n882), .A3(new_n889), .A4(G330), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n912), .B1(new_n1053), .B2(new_n899), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n911), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n302), .A2(new_n324), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n292), .A2(new_n658), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1099), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1110), .A2(new_n1111), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1098), .B1(new_n1112), .B2(KEYINPUT57), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n680), .B1(new_n1112), .B2(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1095), .A2(new_n1093), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1111), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1108), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT57), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(KEYINPUT125), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1113), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n771), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n772), .B1(new_n821), .B2(G50), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n336), .A2(G41), .ZN(new_n1124));
  AOI211_X1 g0924(.A(G50), .B(new_n1124), .C1(new_n250), .C2(new_n454), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n759), .B2(new_n203), .C1(new_n728), .C2(new_n316), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n757), .A2(new_n1012), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(G97), .C2(new_n742), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n734), .A2(new_n202), .B1(new_n594), .B2(new_n738), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G107), .B2(new_n754), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(new_n557), .C2(new_n745), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT58), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1125), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G132), .A2(new_n742), .B1(new_n744), .B2(G137), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT123), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n727), .A2(new_n1072), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT124), .Z(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G150), .B2(new_n725), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G125), .A2(new_n739), .B1(new_n754), .B2(G128), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1134), .B1(new_n386), .B2(new_n734), .C1(new_n1141), .C2(KEYINPUT59), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1133), .B1(new_n1132), .B2(new_n1131), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1123), .B1(new_n1144), .B2(new_n768), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1109), .B2(new_n784), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1122), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1121), .A2(new_n1147), .ZN(G375));
  NAND2_X1  g0948(.A1(new_n1091), .A2(new_n771), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n772), .B1(new_n821), .B2(G68), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1012), .A2(new_n750), .B1(new_n738), .B2(new_n760), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G303), .B2(new_n747), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n744), .A2(G107), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n742), .A2(G116), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n255), .B(new_n1004), .C1(new_n728), .C2(new_n207), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G77), .B2(new_n733), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n751), .A2(new_n925), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n336), .B1(new_n759), .B2(new_n201), .C1(new_n728), .C2(new_n386), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G58), .B2(new_n733), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n739), .A2(G132), .B1(new_n747), .B2(G128), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G150), .A2(new_n744), .B1(new_n742), .B2(new_n1072), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1150), .B1(new_n1164), .B2(new_n768), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n846), .B2(new_n784), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1149), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT126), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n975), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(G381));
  INV_X1    g0972(.A(G375), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1096), .A2(new_n1094), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1060), .A2(new_n1084), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  OR4_X1    g0977(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1178));
  OR4_X1    g0978(.A1(G387), .A2(new_n1177), .A3(G381), .A4(new_n1178), .ZN(G407));
  OAI211_X1 g0979(.A(G407), .B(G213), .C1(G343), .C2(new_n1177), .ZN(G409));
  NAND3_X1  g0980(.A1(new_n1121), .A2(G378), .A3(new_n1147), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1112), .A2(new_n975), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1147), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1176), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(G213), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(G343), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n831), .B(KEYINPUT104), .Z(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1169), .A2(new_n1191), .ZN(new_n1192));
  OR3_X1    g0992(.A1(new_n1091), .A2(new_n1093), .A3(new_n1191), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n679), .A3(new_n1170), .A4(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1190), .A2(new_n1168), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1190), .B1(new_n1168), .B2(new_n1194), .ZN(new_n1197));
  INV_X1    g0997(.A(G2897), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1196), .A2(new_n1197), .B1(new_n1198), .B2(new_n1188), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1168), .A2(new_n1194), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(G384), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1201), .A2(G2897), .A3(new_n1187), .A4(new_n1195), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT61), .B1(new_n1189), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT63), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1189), .B2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(G393), .B(new_n794), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1027), .A2(new_n1028), .A3(new_n1047), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1025), .A2(new_n965), .A3(new_n1021), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n722), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n975), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n990), .B1(new_n1213), .B2(new_n770), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n953), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1210), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(G390), .B(new_n953), .C1(new_n976), .C2(new_n990), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT127), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1209), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(KEYINPUT127), .B(new_n1208), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1187), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1206), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT63), .A3(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1204), .A2(new_n1207), .A3(new_n1222), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT62), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1223), .A2(new_n1227), .A3(new_n1224), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1227), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1228), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1226), .B1(new_n1233), .B2(new_n1222), .ZN(G405));
  INV_X1    g1034(.A(new_n1176), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1181), .B1(new_n1173), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1206), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1224), .B(new_n1181), .C1(new_n1173), .C2(new_n1235), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(new_n1222), .ZN(G402));
endmodule


