//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(KEYINPUT16), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n187), .B(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n198), .B2(G128), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT77), .A3(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT76), .B1(new_n199), .B2(KEYINPUT23), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n205), .A2(new_n206), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n212), .A2(G110), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n199), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT24), .B(G110), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n197), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n191), .A2(new_n192), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n193), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(G110), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n214), .A2(new_n215), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT79), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n218), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n228), .ZN(new_n230));
  INV_X1    g044(.A(new_n223), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n217), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT74), .B(G902), .Z(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G234), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n236), .B(KEYINPUT75), .Z(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G902), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT81), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(new_n240), .B(KEYINPUT82), .Z(new_n241));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n229), .A2(new_n235), .A3(new_n232), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT25), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n237), .B1(new_n243), .B2(KEYINPUT25), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n243), .A2(KEYINPUT25), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(KEYINPUT80), .A3(new_n244), .A4(new_n237), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G472), .A2(G902), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT31), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n192), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n256), .A2(KEYINPUT1), .A3(new_n203), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT65), .B(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT1), .B1(new_n254), .B2(G146), .ZN(new_n260));
  AOI221_X4 g074(.A(KEYINPUT66), .B1(new_n253), .B2(new_n255), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n208), .B2(new_n207), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n258), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n258), .C1(new_n261), .C2(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G137), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G134), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n270), .A2(new_n271), .ZN(new_n276));
  OAI21_X1  g090(.A(G131), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(KEYINPUT11), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT11), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n273), .A3(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n266), .A2(new_n268), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT2), .B(G113), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(G116), .B(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n198), .A2(G116), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n198), .A2(G116), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(KEYINPUT0), .A2(G128), .ZN(new_n300));
  OR2_X1    g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n256), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G143), .B(G146), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT0), .A3(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n281), .A2(new_n270), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n307), .B2(new_n283), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n286), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G210), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G101), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT70), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n319), .B(new_n316), .C1(new_n286), .C2(new_n309), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n299), .ZN(new_n322));
  INV_X1    g136(.A(new_n308), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n286), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT30), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  INV_X1    g140(.A(new_n264), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n263), .A2(new_n262), .A3(new_n256), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n257), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n323), .B(new_n326), .C1(new_n329), .C2(new_n284), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n322), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n252), .B1(new_n321), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n286), .B2(new_n323), .ZN(new_n333));
  INV_X1    g147(.A(new_n330), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n299), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n335), .B(KEYINPUT31), .C1(new_n318), .C2(new_n320), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n324), .A2(KEYINPUT71), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n299), .B1(new_n324), .B2(KEYINPUT71), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT28), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n329), .A2(new_n284), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n299), .B1(new_n342), .B2(new_n308), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n310), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n316), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n337), .A2(KEYINPUT72), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT72), .B1(new_n337), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n251), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT73), .B(new_n251), .C1(new_n346), .C2(new_n347), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G472), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n335), .A2(new_n310), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n316), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n340), .A2(new_n344), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n355), .B(new_n357), .C1(new_n358), .C2(new_n316), .ZN(new_n359));
  INV_X1    g173(.A(new_n235), .ZN(new_n360));
  INV_X1    g174(.A(new_n324), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n310), .B1(new_n361), .B2(new_n322), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(KEYINPUT28), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(new_n340), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n316), .A2(new_n355), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n354), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n251), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n337), .A2(new_n345), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n337), .A2(KEYINPUT72), .A3(new_n345), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(KEYINPUT32), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n250), .B1(new_n353), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G104), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n379), .B(new_n380), .C1(new_n382), .C2(KEYINPUT84), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT84), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT83), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(KEYINPUT83), .A3(G104), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n383), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n382), .B2(new_n392), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(KEYINPUT86), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n391), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n384), .A2(KEYINPUT84), .A3(G107), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT3), .B(new_n388), .C1(new_n399), .C2(KEYINPUT83), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n400), .B2(new_n383), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n397), .B1(new_n401), .B2(new_n394), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(new_n329), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n401), .A2(new_n394), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n203), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n258), .B1(new_n303), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n307), .A2(new_n283), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT12), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(KEYINPUT12), .A3(new_n409), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT12), .B1(new_n408), .B2(new_n409), .ZN(new_n416));
  INV_X1    g230(.A(new_n409), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n411), .B(new_n417), .C1(new_n403), .C2(new_n407), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT88), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n266), .A2(new_n268), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT86), .B1(new_n393), .B2(new_n395), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n401), .A2(new_n397), .A3(new_n394), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT87), .B1(new_n396), .B2(new_n402), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT10), .B(new_n420), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n400), .A2(new_n383), .B1(new_n384), .B2(G107), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n393), .B(KEYINPUT4), .C1(new_n391), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n390), .A2(new_n392), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT85), .B(KEYINPUT4), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(G101), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n428), .A2(new_n304), .A3(new_n302), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n407), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n426), .A2(new_n436), .A3(new_n417), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  INV_X1    g252(.A(G227), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G953), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n415), .A2(new_n419), .A3(new_n437), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n417), .B1(new_n426), .B2(new_n436), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n266), .A2(KEYINPUT10), .A3(new_n268), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n423), .B1(new_n421), .B2(new_n422), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n402), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n433), .A2(new_n435), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n448), .A2(new_n409), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n441), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n360), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G469), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n416), .A2(new_n418), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n441), .B1(new_n450), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n442), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(new_n444), .ZN(new_n462));
  INV_X1    g276(.A(G902), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G469), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n378), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT90), .Z(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G113), .B1(new_n291), .B2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n289), .A2(KEYINPUT5), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(new_n288), .B2(new_n289), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n446), .B2(new_n447), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n428), .A2(new_n299), .A3(new_n432), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n474), .B1(new_n424), .B2(new_n425), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n477), .A3(new_n469), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT6), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n470), .C1(new_n476), .C2(new_n478), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n305), .A2(G125), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n265), .B2(G125), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n224), .A2(G224), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n486), .B(new_n487), .Z(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n485), .A2(KEYINPUT92), .B1(KEYINPUT7), .B2(new_n487), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n486), .B(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n421), .A2(new_n422), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n472), .A2(KEYINPUT91), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n473), .B1(new_n472), .B2(KEYINPUT91), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n290), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n492), .A2(new_n495), .B1(new_n404), .B2(new_n474), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n469), .B(KEYINPUT8), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n498), .B2(new_n481), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n489), .A2(new_n499), .A3(new_n501), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n468), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n466), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n384), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT19), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n195), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n509), .B2(new_n187), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n193), .B1(new_n511), .B2(G146), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT96), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n312), .A2(G214), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n254), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n312), .B(G214), .C1(KEYINPUT93), .C2(G143), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT95), .A3(new_n282), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n518), .B2(G131), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n520), .B(new_n522), .C1(new_n282), .C2(new_n519), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n193), .C1(new_n511), .C2(G146), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT94), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n187), .A2(new_n192), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n196), .A2(new_n530), .B1(new_n527), .B2(new_n518), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n508), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n220), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(KEYINPUT17), .A3(G131), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n534), .B(new_n535), .C1(new_n523), .C2(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n532), .ZN(new_n537));
  INV_X1    g351(.A(new_n508), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G475), .A2(G902), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n541), .B(KEYINPUT97), .Z(new_n542));
  OAI21_X1  g356(.A(KEYINPUT20), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  INV_X1    g358(.A(new_n542), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n544), .B(new_n545), .C1(new_n533), .C2(new_n539), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n508), .B1(new_n536), .B2(new_n532), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n463), .B1(new_n539), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n543), .A2(new_n546), .B1(G475), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n209), .A2(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n254), .A2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n269), .ZN(new_n553));
  XOR2_X1   g367(.A(G116), .B(G122), .Z(new_n554));
  INV_X1    g368(.A(G122), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G116), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n381), .B1(new_n556), .B2(KEYINPUT14), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n554), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n551), .B(KEYINPUT13), .Z(new_n559));
  INV_X1    g373(.A(new_n550), .ZN(new_n560));
  OAI21_X1  g374(.A(G134), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n554), .B(G107), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n552), .A2(G134), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n553), .A2(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n376), .A2(new_n234), .A3(G953), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n360), .ZN(new_n568));
  INV_X1    g382(.A(G478), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n568), .A2(new_n570), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n549), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT98), .B(G952), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  NAND2_X1  g390(.A1(G234), .A2(G237), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n360), .A2(G953), .A3(new_n577), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT21), .B(G898), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n375), .A2(new_n506), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AND2_X1   g400(.A1(new_n350), .A2(new_n352), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n235), .B1(new_n346), .B2(new_n347), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  INV_X1    g403(.A(new_n250), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n443), .A2(new_n451), .ZN(new_n591));
  AND4_X1   g405(.A1(KEYINPUT89), .A2(new_n591), .A3(new_n453), .A4(new_n235), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT89), .B1(new_n452), .B2(new_n453), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n465), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n590), .A2(new_n594), .A3(new_n377), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n589), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT99), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n504), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n501), .B1(new_n489), .B2(new_n499), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n500), .A2(KEYINPUT100), .A3(new_n502), .ZN(new_n602));
  INV_X1    g416(.A(new_n468), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n583), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n543), .A2(new_n546), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n548), .A2(G475), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n568), .A2(G478), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n567), .B(KEYINPUT33), .Z(new_n612));
  NOR2_X1   g426(.A1(new_n360), .A2(new_n569), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n597), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n573), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n549), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n607), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n597), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NAND2_X1  g440(.A1(new_n218), .A2(new_n223), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n239), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n247), .A2(new_n249), .A3(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n574), .A2(new_n631), .A3(new_n583), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n506), .A2(new_n587), .A3(new_n589), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(new_n631), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n594), .A2(new_n377), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n353), .B2(new_n374), .ZN(new_n638));
  INV_X1    g452(.A(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n581), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n578), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n622), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n605), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XNOR2_X1  g460(.A(new_n641), .B(KEYINPUT39), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n466), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT40), .Z(new_n649));
  OAI21_X1  g463(.A(new_n335), .B1(new_n318), .B2(new_n320), .ZN(new_n650));
  INV_X1    g464(.A(new_n362), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n317), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n354), .B1(new_n652), .B2(new_n463), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n373), .B2(KEYINPUT32), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n353), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n503), .A2(new_n504), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n610), .A2(new_n621), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(new_n468), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n649), .A2(new_n631), .A3(new_n655), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NAND2_X1  g476(.A1(new_n353), .A2(new_n374), .ZN(new_n663));
  INV_X1    g477(.A(new_n637), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n549), .A2(new_n614), .A3(new_n642), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n468), .B1(new_n599), .B2(new_n600), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n503), .A2(new_n598), .A3(new_n504), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n663), .A2(new_n664), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  OR2_X1    g486(.A1(new_n452), .A2(new_n453), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n377), .B(new_n673), .C1(new_n592), .C2(new_n593), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT101), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n375), .A2(new_n617), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NAND3_X1  g492(.A1(new_n375), .A2(new_n623), .A3(new_n675), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT102), .B(G116), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G18));
  NOR2_X1   g495(.A1(new_n669), .A2(new_n674), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n663), .A2(new_n632), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT103), .B(G119), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n363), .B2(new_n340), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n362), .A2(KEYINPUT28), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n338), .A2(new_n339), .ZN(new_n689));
  OAI211_X1 g503(.A(KEYINPUT104), .B(new_n688), .C1(new_n689), .C2(KEYINPUT28), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n690), .A3(new_n316), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n368), .B1(new_n691), .B2(new_n337), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n589), .A2(new_n590), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n607), .A3(new_n659), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n675), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(KEYINPUT105), .A3(new_n675), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  NAND4_X1  g515(.A1(new_n589), .A2(new_n636), .A3(new_n665), .A4(new_n693), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n605), .A2(new_n377), .A3(new_n458), .A4(new_n673), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT106), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n631), .B(new_n692), .C1(new_n588), .C2(G472), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n682), .A3(new_n706), .A4(new_n665), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n373), .B2(KEYINPUT32), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n348), .A2(KEYINPUT108), .A3(new_n351), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n374), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT107), .B1(new_n656), .B2(new_n468), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n503), .A2(new_n715), .A3(new_n603), .A4(new_n504), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n714), .A2(new_n594), .A3(new_n377), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n713), .A2(new_n718), .A3(new_n590), .A4(new_n665), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n375), .A2(new_n718), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n282), .ZN(G33));
  NAND3_X1  g538(.A1(new_n375), .A2(new_n643), .A3(new_n718), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  NOR2_X1   g540(.A1(new_n610), .A2(new_n614), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n631), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n587), .A2(new_n589), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(KEYINPUT44), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n714), .A2(new_n716), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n453), .B1(new_n462), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n736), .B2(new_n462), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n458), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n377), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n647), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n730), .A2(new_n731), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n735), .B(new_n747), .C1(KEYINPUT44), .C2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  NOR4_X1   g564(.A1(new_n663), .A2(new_n733), .A3(new_n590), .A4(new_n666), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n745), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  NAND2_X1  g571(.A1(new_n616), .A2(new_n622), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(new_n505), .A3(new_n606), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n587), .A3(new_n595), .A4(new_n589), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n585), .A2(new_n633), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n585), .A2(new_n633), .A3(new_n763), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n733), .A2(new_n574), .A3(new_n642), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n638), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n702), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT112), .B1(new_n768), .B2(new_n718), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n702), .A2(new_n717), .A3(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n725), .B(new_n767), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n723), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n676), .A2(new_n679), .A3(new_n683), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n699), .B2(new_n698), .ZN(new_n775));
  AND4_X1   g589(.A1(KEYINPUT53), .A2(new_n765), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n594), .A2(new_n377), .A3(new_n641), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n667), .A2(new_n621), .A3(new_n610), .A4(new_n668), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n655), .A2(new_n631), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n708), .A2(new_n645), .A3(new_n671), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n708), .A2(new_n645), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n671), .A2(new_n782), .A3(KEYINPUT52), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT113), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n704), .A2(new_n707), .B1(new_n638), .B2(new_n644), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n778), .B1(new_n638), .B2(new_n670), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n782), .A4(new_n789), .ZN(new_n790));
  AOI221_X4 g604(.A(new_n777), .B1(new_n778), .B2(new_n783), .C1(new_n786), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n783), .A2(new_n778), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT114), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n776), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n765), .A2(new_n773), .A3(new_n775), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n787), .A2(new_n782), .A3(new_n789), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n795), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n729), .A2(new_n578), .A3(new_n694), .ZN(new_n805));
  INV_X1    g619(.A(new_n658), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n603), .A3(new_n674), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n809));
  AND2_X1   g623(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n655), .A2(new_n250), .A3(new_n578), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n733), .A2(new_n674), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n549), .A3(new_n614), .A4(new_n813), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n729), .A2(new_n578), .A3(new_n674), .A4(new_n733), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n808), .A2(new_n809), .B1(new_n815), .B2(new_n705), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n805), .A2(new_n734), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n458), .A2(new_n673), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT110), .Z(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n377), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n754), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n804), .B1(new_n817), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n713), .A2(new_n590), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT48), .Z(new_n828));
  NAND2_X1  g642(.A1(new_n805), .A2(new_n682), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n812), .A2(new_n813), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n576), .B(new_n829), .C1(new_n830), .C2(new_n616), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n817), .A2(new_n824), .A3(new_n804), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n798), .A2(new_n801), .A3(new_n797), .ZN(new_n836));
  INV_X1    g650(.A(new_n798), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n791), .B2(new_n794), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n838), .B2(new_n797), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n803), .B(new_n835), .C1(new_n839), .C2(new_n796), .ZN(new_n840));
  INV_X1    g654(.A(G952), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n224), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n821), .B(KEYINPUT49), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n590), .A2(new_n727), .A3(new_n377), .A4(new_n603), .ZN(new_n845));
  OR4_X1    g659(.A1(new_n655), .A2(new_n844), .A3(new_n806), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(KEYINPUT117), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(G75));
  NAND2_X1  g665(.A1(new_n482), .A2(new_n484), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(new_n488), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n765), .A2(new_n773), .A3(new_n775), .A4(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n792), .A2(new_n793), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n777), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n792), .A2(KEYINPUT114), .A3(new_n793), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n802), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n360), .B(new_n502), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n861), .B2(new_n862), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n854), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n841), .A2(G953), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT119), .Z(new_n869));
  AOI211_X1 g683(.A(new_n235), .B(new_n501), .C1(new_n795), .C2(new_n802), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n863), .B1(new_n870), .B2(KEYINPUT56), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n853), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n867), .A2(new_n869), .A3(new_n873), .ZN(G51));
  INV_X1    g688(.A(new_n869), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n795), .A2(new_n802), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n803), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n876), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n739), .B(KEYINPUT120), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT57), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n591), .ZN(new_n884));
  INV_X1    g698(.A(new_n876), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n885), .A2(new_n235), .A3(new_n738), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n875), .B1(new_n884), .B2(new_n886), .ZN(G54));
  NAND4_X1  g701(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .A4(new_n360), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n888), .A2(KEYINPUT122), .A3(new_n540), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n869), .B1(new_n888), .B2(new_n540), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT122), .B1(new_n888), .B2(new_n540), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT59), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n612), .A2(new_n879), .A3(new_n880), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n803), .B1(new_n839), .B2(new_n796), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n612), .B1(new_n896), .B2(new_n894), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n875), .A3(new_n897), .ZN(G63));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT123), .Z(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT60), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n876), .A2(new_n629), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n875), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n233), .ZN(new_n909));
  INV_X1    g723(.A(new_n901), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n885), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n906), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n906), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(G66));
  INV_X1    g728(.A(G224), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n582), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n765), .A2(new_n775), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n852), .B1(G898), .B2(new_n224), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  INV_X1    g735(.A(new_n780), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n747), .A2(new_n826), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n749), .A2(new_n725), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n754), .A2(new_n755), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n723), .B1(new_n925), .B2(new_n752), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n787), .A2(new_n671), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(G953), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n333), .A2(new_n334), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n511), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n639), .B2(new_n224), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n648), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n375), .A2(new_n934), .A3(new_n734), .A4(new_n758), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n749), .A2(new_n756), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n661), .A2(new_n927), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n931), .B1(new_n940), .B2(new_n224), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n439), .B2(new_n639), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G72));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n928), .B2(new_n917), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n356), .A2(new_n317), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT126), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n875), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(new_n940), .B2(new_n917), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n356), .A2(new_n317), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n955));
  INV_X1    g769(.A(new_n946), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n357), .B2(new_n650), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n955), .B1(new_n839), .B2(new_n958), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n839), .A2(new_n955), .A3(new_n958), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(G57));
endmodule


