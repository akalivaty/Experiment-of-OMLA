//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT39), .ZN(new_n202));
  AND2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n207));
  OAI21_X1  g006(.A(G162gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n205), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT78), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n213), .A3(G141gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n210), .A2(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT77), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(new_n210), .B2(G141gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT76), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n204), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G155gat), .A3(G162gat), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G148gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n215), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  OR3_X1    g038(.A1(new_n239), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n233), .A4(new_n240), .ZN(new_n241));
  AND4_X1   g040(.A1(new_n220), .A2(new_n232), .A3(new_n236), .A4(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n220), .A2(new_n232), .B1(new_n241), .B2(new_n236), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT80), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n202), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n248), .A2(KEYINPUT88), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n232), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n240), .A2(new_n233), .A3(new_n238), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n254), .A2(new_n237), .B1(new_n255), .B2(new_n234), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n209), .A2(new_n219), .B1(new_n227), .B2(new_n231), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT4), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(new_n251), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n247), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n248), .A2(KEYINPUT88), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n264), .B2(new_n202), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT40), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n252), .B1(new_n250), .B2(new_n251), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n257), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n263), .A2(new_n247), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n246), .B1(new_n242), .B2(new_n243), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n259), .A2(KEYINPUT5), .A3(new_n247), .A4(new_n263), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n271), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n267), .A2(KEYINPUT40), .A3(new_n272), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n275), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(G211gat), .A2(G218gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G211gat), .A2(G218gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n296), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT27), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT28), .A4(new_n308), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT66), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n309), .A2(new_n322), .A3(new_n310), .ZN(new_n323));
  AND4_X1   g122(.A1(new_n303), .A2(new_n313), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n303), .ZN(new_n326));
  NAND3_X1  g125(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  INV_X1    g128(.A(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT25), .A4(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n315), .B2(KEYINPUT23), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n332), .A2(G169gat), .A3(G176gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT65), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n331), .A2(new_n333), .A3(new_n340), .A4(new_n334), .ZN(new_n341));
  NAND4_X1  g140(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n336), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n324), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n302), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n324), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n347), .ZN(new_n355));
  INV_X1    g154(.A(new_n336), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n313), .A2(new_n321), .A3(new_n303), .A4(new_n323), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT72), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n352), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n351), .B1(new_n360), .B2(new_n350), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n353), .B1(new_n324), .B2(new_n348), .ZN(new_n362));
  INV_X1    g161(.A(new_n350), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n325), .A2(new_n303), .B1(new_n327), .B2(new_n343), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n342), .A2(new_n364), .B1(new_n365), .B2(KEYINPUT65), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT25), .B1(new_n366), .B2(new_n341), .ZN(new_n367));
  OAI211_X1 g166(.A(KEYINPUT72), .B(new_n358), .C1(new_n367), .C2(new_n336), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n302), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n357), .A2(new_n358), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n352), .A3(new_n350), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n289), .B1(new_n361), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n371), .B2(new_n363), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n362), .B2(new_n368), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n363), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n288), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT30), .A4(new_n288), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT73), .B(new_n289), .C1(new_n361), .C2(new_n373), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n376), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT87), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n385), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n383), .A4(new_n376), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n285), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(KEYINPUT89), .B(KEYINPUT38), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n288), .B1(new_n379), .B2(new_n380), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT37), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n288), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n379), .B2(new_n380), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n281), .A2(new_n271), .A3(new_n282), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n283), .A2(new_n400), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n271), .B1(new_n281), .B2(new_n282), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n381), .B(new_n402), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n369), .A2(new_n302), .A3(new_n372), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n378), .A2(new_n363), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n370), .B1(new_n349), .B2(new_n350), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(KEYINPUT37), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(new_n392), .C1(new_n394), .C2(new_n396), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n399), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n302), .B1(new_n262), .B2(new_n352), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n297), .B2(new_n301), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n261), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n297), .C2(new_n301), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n250), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(KEYINPUT83), .B(new_n250), .C1(new_n418), .C2(new_n419), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n257), .B2(new_n261), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n370), .B1(new_n425), .B2(KEYINPUT85), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  AOI211_X1 g226(.A(new_n427), .B(KEYINPUT29), .C1(new_n257), .C2(new_n261), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n250), .B1(KEYINPUT3), .B2(new_n416), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n250), .B(KEYINPUT84), .C1(KEYINPUT3), .C2(new_n416), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n414), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(G22gat), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n437));
  INV_X1    g236(.A(new_n415), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n423), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n413), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n432), .A2(new_n414), .A3(new_n433), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n427), .B1(new_n443), .B2(KEYINPUT29), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n425), .A2(KEYINPUT85), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n370), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n436), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n439), .A2(new_n413), .B1(new_n442), .B2(new_n446), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n441), .ZN(new_n452));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G50gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n449), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n448), .A3(new_n450), .A4(new_n455), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n412), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n391), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT74), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n385), .A2(new_n384), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n394), .A2(KEYINPUT73), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n404), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n283), .A3(new_n400), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n467), .A2(new_n402), .B1(new_n381), .B2(new_n382), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n376), .A2(KEYINPUT74), .A3(new_n384), .A4(new_n385), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n457), .A2(new_n458), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT70), .ZN(new_n475));
  INV_X1    g274(.A(G15gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(G43gat), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n256), .B(new_n358), .C1(new_n367), .C2(new_n336), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT69), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n357), .A2(new_n481), .A3(new_n256), .A4(new_n358), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n251), .B1(new_n324), .B2(new_n348), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n478), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n256), .B1(new_n357), .B2(new_n358), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(KEYINPUT69), .B2(new_n479), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n485), .B2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n485), .A3(new_n482), .A4(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n480), .A2(new_n485), .A3(new_n482), .A4(new_n483), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT33), .B1(new_n484), .B2(new_n486), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n495), .B(new_n497), .C1(new_n502), .C2(new_n478), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n499), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n473), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n499), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n500), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT36), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n472), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR4_X1   g314(.A1(new_n471), .A2(new_n504), .A3(new_n515), .A4(new_n505), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n387), .A2(new_n390), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n504), .A2(new_n505), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n459), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT35), .B1(new_n520), .B2(new_n470), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n461), .A2(new_n512), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n523), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n524), .A3(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G8gat), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n539));
  AOI21_X1  g338(.A(G36gat), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n536), .A2(new_n541), .A3(G29gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n545));
  OAI221_X1 g344(.A(new_n535), .B1(new_n540), .B2(new_n542), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n540), .A2(new_n542), .B1(KEYINPUT15), .B2(new_n534), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n540), .B2(new_n542), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n543), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT17), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT17), .B1(new_n546), .B2(new_n549), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n531), .B(new_n533), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT93), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n531), .A2(new_n533), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n546), .A3(new_n549), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT94), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n552), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n556), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n549), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n531), .A3(new_n533), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n554), .B(KEYINPUT13), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n557), .A2(new_n569), .A3(new_n558), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n560), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n572));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G197gat), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT11), .B(G169gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT90), .B(KEYINPUT12), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n571), .A2(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n559), .A2(new_n578), .A3(new_n567), .A4(new_n561), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT95), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n580), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n522), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT107), .B(KEYINPUT10), .Z(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n588), .B1(new_n595), .B2(KEYINPUT105), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n594), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT105), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n588), .A3(new_n594), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n590), .A2(KEYINPUT104), .A3(new_n588), .A4(new_n594), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n596), .A2(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G64gat), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n605), .A2(G57gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT99), .B(G57gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(G64gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G71gat), .B(G78gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n610), .A2(new_n611), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n605), .A2(G57gat), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT96), .B1(new_n606), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G57gat), .B(G64gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n614), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT98), .B1(new_n623), .B2(new_n615), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(KEYINPUT98), .A3(new_n615), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n604), .B(new_n617), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n617), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n603), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n588), .B2(new_n595), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n625), .A2(new_n624), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n633), .A2(new_n604), .A3(KEYINPUT106), .A4(new_n617), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n587), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n627), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n586), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n586), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n632), .A2(new_n642), .A3(new_n634), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT108), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n632), .A2(KEYINPUT108), .A3(new_n642), .A4(new_n634), .ZN(new_n646));
  AND4_X1   g445(.A1(new_n638), .A2(new_n641), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n641), .B1(new_n638), .B2(new_n643), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT109), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n641), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n596), .A2(new_n599), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n628), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n631), .B1(new_n627), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n627), .A2(new_n629), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n634), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n587), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n637), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n642), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n643), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n651), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n638), .A2(new_n641), .A3(new_n645), .A4(new_n646), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT109), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n650), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT21), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n531), .B(new_n533), .C1(new_n627), .C2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT102), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n627), .A2(new_n667), .ZN(new_n670));
  XOR2_X1   g469(.A(G127gat), .B(G155gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n669), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G231gat), .A2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT101), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G183gat), .B(G211gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n673), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n629), .A2(new_n562), .ZN(new_n681));
  AND2_X1   g480(.A1(G232gat), .A2(G233gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(KEYINPUT41), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n629), .B1(new_n550), .B2(new_n551), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(G190gat), .B(G218gat), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n685), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n682), .A2(KEYINPUT41), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT103), .ZN(new_n690));
  XOR2_X1   g489(.A(G134gat), .B(G162gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n688), .B(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n666), .A2(new_n680), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n585), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n513), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n526), .ZN(G1324gat));
  INV_X1    g496(.A(new_n695), .ZN(new_n698));
  INV_X1    g497(.A(new_n517), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n532), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT16), .B(G8gat), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n695), .A2(new_n517), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT42), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(KEYINPUT42), .B2(new_n702), .ZN(G1325gat));
  AOI21_X1  g503(.A(G15gat), .B1(new_n698), .B2(new_n519), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n511), .A2(new_n476), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT110), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n698), .B2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n695), .A2(new_n459), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n472), .B(new_n511), .C1(new_n391), .C2(new_n460), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n513), .A2(new_n383), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n376), .A2(new_n384), .A3(new_n385), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n462), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n717), .A2(new_n459), .A3(new_n519), .A4(new_n469), .ZN(new_n718));
  AOI22_X1  g517(.A1(KEYINPUT35), .A2(new_n718), .B1(new_n516), .B2(new_n517), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n712), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n518), .A2(new_n521), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(KEYINPUT111), .A3(new_n713), .ZN(new_n722));
  INV_X1    g521(.A(new_n693), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(KEYINPUT44), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT44), .B1(new_n522), .B2(new_n723), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n665), .A2(new_n680), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n584), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT112), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  INV_X1    g530(.A(new_n729), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n731), .B(new_n732), .C1(new_n725), .C2(new_n726), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n513), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n537), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n522), .A2(new_n732), .A3(new_n723), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n537), .A3(new_n735), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT45), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT113), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n730), .A2(new_n733), .A3(new_n513), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n742), .B(new_n739), .C1(new_n743), .C2(new_n537), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(G1328gat));
  NAND3_X1  g544(.A1(new_n737), .A2(new_n541), .A3(new_n699), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n733), .A3(new_n517), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n541), .ZN(G1329gat));
  NAND2_X1  g548(.A1(new_n727), .A2(new_n729), .ZN(new_n750));
  OAI21_X1  g549(.A(G43gat), .B1(new_n750), .B2(new_n511), .ZN(new_n751));
  INV_X1    g550(.A(new_n519), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(G43gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n754), .ZN(new_n756));
  INV_X1    g555(.A(new_n511), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n734), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n758), .B2(G43gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g559(.A(G50gat), .B1(new_n750), .B2(new_n459), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n723), .A2(G50gat), .A3(new_n459), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n522), .A2(new_n584), .A3(new_n728), .A4(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n734), .A2(new_n471), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n767), .B2(G50gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g568(.A(new_n583), .B1(new_n579), .B2(new_n571), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n571), .A2(new_n572), .A3(new_n579), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n680), .A2(new_n772), .A3(new_n693), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n720), .A2(new_n666), .A3(new_n722), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n513), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(new_n607), .ZN(G1332gat));
  AOI211_X1 g575(.A(new_n517), .B(new_n774), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT114), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT115), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n777), .B(new_n780), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n774), .B2(new_n511), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n752), .A2(G71gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g584(.A1(new_n774), .A2(new_n459), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g586(.A1(new_n522), .A2(new_n723), .ZN(new_n788));
  INV_X1    g587(.A(new_n680), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n772), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n788), .A2(new_n790), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n795), .A2(new_n592), .A3(new_n735), .A4(new_n666), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n727), .A2(new_n666), .A3(new_n790), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n513), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n592), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT117), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n796), .B(new_n801), .C1(new_n592), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1336gat));
  INV_X1    g602(.A(new_n797), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n517), .A2(new_n593), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n804), .A2(new_n805), .B1(KEYINPUT118), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n808));
  INV_X1    g607(.A(new_n792), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n788), .A2(new_n790), .B1(KEYINPUT116), .B2(KEYINPUT51), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n699), .B(new_n666), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n593), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n807), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n808), .B1(new_n807), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n797), .B2(new_n511), .ZN(new_n816));
  INV_X1    g615(.A(G99gat), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n665), .A2(new_n752), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n795), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(G1338gat));
  NOR2_X1   g619(.A1(new_n459), .A2(G106gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n795), .A2(new_n666), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n797), .A2(new_n459), .ZN(new_n823));
  INV_X1    g622(.A(G106gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n658), .A2(new_n642), .A3(new_n659), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n638), .A3(KEYINPUT54), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n651), .B1(new_n638), .B2(KEYINPUT54), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n641), .B1(new_n660), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n829), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n772), .A2(new_n832), .A3(new_n663), .A4(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n552), .A2(new_n556), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n837), .A2(new_n554), .B1(new_n564), .B2(new_n566), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n576), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n582), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n650), .B2(new_n664), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT119), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n846), .A3(new_n723), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n693), .A3(new_n835), .A4(new_n663), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n840), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n789), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n773), .A2(new_n665), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n513), .ZN(new_n855));
  INV_X1    g654(.A(new_n520), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n517), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(new_n584), .ZN(new_n858));
  INV_X1    g657(.A(G113gat), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n836), .A2(new_n842), .A3(new_n845), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n845), .B1(new_n836), .B2(new_n842), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n860), .A2(new_n861), .A3(new_n693), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n680), .B1(new_n862), .B2(new_n849), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n852), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n517), .A2(new_n735), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n520), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n584), .A2(new_n859), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n858), .A2(new_n859), .B1(new_n868), .B2(new_n869), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n867), .B2(new_n665), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n665), .A2(G120gat), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT120), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n857), .B2(new_n873), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n867), .B2(new_n680), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n680), .A2(G127gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n857), .B2(new_n876), .ZN(G1342gat));
  NAND3_X1  g676(.A1(new_n864), .A2(new_n735), .A3(new_n856), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n699), .A2(new_n723), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(G134gat), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT121), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n855), .A2(new_n884), .A3(new_n856), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G134gat), .B1(new_n867), .B2(new_n723), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT56), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G1343gat));
  NOR2_X1   g690(.A1(new_n865), .A2(new_n757), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n584), .A2(new_n229), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n864), .B2(new_n471), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n459), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n835), .A2(new_n663), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n832), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n834), .A2(new_n829), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(KEYINPUT122), .A3(new_n827), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n899), .A2(new_n901), .A3(new_n903), .A4(new_n772), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n693), .B1(new_n904), .B2(new_n842), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n680), .B1(new_n905), .B2(new_n849), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n897), .B1(new_n906), .B2(new_n852), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n757), .A2(new_n459), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n864), .A2(new_n735), .A3(new_n517), .A4(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n229), .B1(new_n910), .B2(new_n584), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(KEYINPUT58), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1344gat));
  OAI21_X1  g715(.A(KEYINPUT59), .B1(new_n910), .B2(new_n665), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n211), .A3(new_n213), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n649), .B1(new_n647), .B2(new_n648), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT109), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n840), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT122), .B1(new_n902), .B2(new_n827), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n900), .B(KEYINPUT55), .C1(new_n834), .C2(new_n829), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n898), .A2(new_n584), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n848), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n841), .B1(new_n848), .B2(new_n927), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n926), .A2(new_n693), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n853), .B1(new_n930), .B2(new_n680), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n895), .B1(new_n931), .B2(new_n459), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n896), .B1(new_n851), .B2(new_n853), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n666), .A3(new_n892), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n892), .B1(new_n894), .B2(new_n907), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n665), .A2(KEYINPUT59), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n918), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(G1345gat));
  OAI22_X1  g738(.A1(new_n937), .A2(new_n680), .B1(new_n207), .B2(new_n206), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n680), .A2(new_n207), .A3(new_n206), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n910), .B2(new_n941), .ZN(G1346gat));
  OAI21_X1  g741(.A(G162gat), .B1(new_n937), .B2(new_n723), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n855), .A2(new_n222), .A3(new_n879), .A4(new_n909), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n517), .A2(new_n735), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n864), .A2(new_n856), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n584), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(new_n329), .ZN(G1348gat));
  INV_X1    g748(.A(new_n946), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n854), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n471), .B1(KEYINPUT124), .B2(new_n330), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n818), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n330), .A2(KEYINPUT124), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1349gat));
  OAI21_X1  g754(.A(new_n304), .B1(new_n947), .B2(new_n680), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n305), .A2(new_n307), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n951), .A2(new_n957), .A3(new_n856), .A4(new_n789), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1350gat));
  OAI22_X1  g761(.A1(new_n947), .A2(new_n723), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n963), .B(new_n964), .ZN(G1351gat));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n757), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n967), .A2(new_n584), .ZN(new_n968));
  XOR2_X1   g767(.A(KEYINPUT125), .B(G197gat), .Z(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n928), .A2(new_n929), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n680), .B1(new_n972), .B2(new_n905), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n852), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT57), .B1(new_n974), .B2(new_n471), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n897), .B1(new_n863), .B2(new_n852), .ZN(new_n976));
  OAI21_X1  g775(.A(KEYINPUT126), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n932), .A2(new_n933), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n971), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n854), .A2(new_n459), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n970), .B1(new_n981), .B2(new_n968), .ZN(new_n982));
  OAI21_X1  g781(.A(KEYINPUT127), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n971), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n932), .A2(new_n933), .A3(new_n978), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n978), .B1(new_n932), .B2(new_n933), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  INV_X1    g787(.A(new_n982), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n983), .A2(new_n990), .ZN(G1352gat));
  OAI211_X1 g790(.A(new_n666), .B(new_n966), .C1(new_n985), .C2(new_n986), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G204gat), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n665), .A2(G204gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n981), .A2(new_n966), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n996));
  OR2_X1    g795(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(G1353gat));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n966), .ZN(new_n999));
  OR3_X1    g798(.A1(new_n999), .A2(G211gat), .A3(new_n680), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n934), .A2(new_n789), .A3(new_n966), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(G211gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G1354gat));
  INV_X1    g803(.A(new_n999), .ZN(new_n1005));
  AOI21_X1  g804(.A(G218gat), .B1(new_n1005), .B2(new_n693), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n967), .B1(new_n977), .B2(new_n979), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n693), .A2(G218gat), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(G1355gat));
endmodule


