

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  NOR2_X1 U322 ( .A1(n469), .A2(n468), .ZN(n563) );
  INV_X1 U323 ( .A(n546), .ZN(n559) );
  XNOR2_X1 U324 ( .A(n307), .B(n306), .ZN(n527) );
  XNOR2_X1 U325 ( .A(n445), .B(KEYINPUT38), .ZN(n499) );
  XOR2_X1 U326 ( .A(n297), .B(n296), .Z(n290) );
  INV_X1 U327 ( .A(n416), .ZN(n417) );
  XNOR2_X1 U328 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U329 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U330 ( .A(n298), .B(n290), .ZN(n299) );
  NOR2_X1 U331 ( .A1(n516), .A2(n464), .ZN(n567) );
  XNOR2_X1 U332 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U333 ( .A(n300), .B(n299), .ZN(n305) );
  XNOR2_X1 U334 ( .A(n429), .B(n428), .ZN(n572) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n470) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n446) );
  XNOR2_X1 U337 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U338 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U339 ( .A(n473), .B(n472), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n449), .B(n448), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G176GAT), .B(KEYINPUT20), .Z(n292) );
  XNOR2_X1 U342 ( .A(KEYINPUT81), .B(G169GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n307) );
  XOR2_X1 U344 ( .A(KEYINPUT82), .B(G99GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(G43GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U347 ( .A(n295), .B(KEYINPUT80), .Z(n300) );
  XOR2_X1 U348 ( .A(KEYINPUT0), .B(G127GAT), .Z(n353) );
  XNOR2_X1 U349 ( .A(n353), .B(G120GAT), .ZN(n298) );
  XOR2_X1 U350 ( .A(G71GAT), .B(G15GAT), .Z(n297) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U352 ( .A(G134GAT), .B(G190GAT), .Z(n400) );
  XOR2_X1 U353 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U354 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(G183GAT), .B(n303), .Z(n328) );
  XNOR2_X1 U357 ( .A(n400), .B(n328), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U359 ( .A(KEYINPUT2), .B(G162GAT), .Z(n309) );
  XNOR2_X1 U360 ( .A(G155GAT), .B(G148GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(n310), .Z(n347) );
  XOR2_X1 U363 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(G106GAT), .B(G78GAT), .Z(n416) );
  XOR2_X1 U367 ( .A(n313), .B(n416), .Z(n315) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(G22GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U370 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n317) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U373 ( .A(n319), .B(n318), .Z(n325) );
  XNOR2_X1 U374 ( .A(G204GAT), .B(KEYINPUT85), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n320), .B(G197GAT), .ZN(n321) );
  XOR2_X1 U376 ( .A(n321), .B(KEYINPUT21), .Z(n323) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n327) );
  XNOR2_X1 U379 ( .A(G141GAT), .B(n327), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n347), .B(n326), .ZN(n361) );
  XNOR2_X1 U382 ( .A(KEYINPUT28), .B(n361), .ZN(n529) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n339) );
  XOR2_X1 U384 ( .A(G8GAT), .B(G169GAT), .Z(n435) );
  XOR2_X1 U385 ( .A(KEYINPUT92), .B(KEYINPUT77), .Z(n330) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U388 ( .A(n435), .B(n331), .Z(n333) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U391 ( .A(n334), .B(KEYINPUT90), .Z(n337) );
  XNOR2_X1 U392 ( .A(G92GAT), .B(G64GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n335), .B(G176GAT), .ZN(n414) );
  XNOR2_X1 U394 ( .A(n414), .B(KEYINPUT91), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n483) );
  XNOR2_X1 U397 ( .A(n483), .B(KEYINPUT93), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n340), .B(KEYINPUT27), .ZN(n363) );
  XOR2_X1 U399 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n342) );
  NAND2_X1 U400 ( .A1(G225GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n343), .B(KEYINPUT1), .Z(n349) );
  XOR2_X1 U403 ( .A(KEYINPUT6), .B(KEYINPUT88), .Z(n345) );
  XNOR2_X1 U404 ( .A(G134GAT), .B(G85GAT), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n352) );
  XOR2_X1 U408 ( .A(G1GAT), .B(G113GAT), .Z(n351) );
  XNOR2_X1 U409 ( .A(G29GAT), .B(G141GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n439) );
  XOR2_X1 U411 ( .A(n352), .B(n439), .Z(n355) );
  XOR2_X1 U412 ( .A(G120GAT), .B(G57GAT), .Z(n423) );
  XNOR2_X1 U413 ( .A(n353), .B(n423), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n366) );
  XNOR2_X1 U415 ( .A(KEYINPUT89), .B(n366), .ZN(n516) );
  NAND2_X1 U416 ( .A1(n363), .A2(n516), .ZN(n525) );
  NOR2_X1 U417 ( .A1(n529), .A2(n525), .ZN(n356) );
  XOR2_X1 U418 ( .A(KEYINPUT94), .B(n356), .Z(n357) );
  NOR2_X1 U419 ( .A1(n527), .A2(n357), .ZN(n370) );
  INV_X1 U420 ( .A(n527), .ZN(n469) );
  NOR2_X1 U421 ( .A1(n469), .A2(n483), .ZN(n358) );
  XOR2_X1 U422 ( .A(KEYINPUT95), .B(n358), .Z(n359) );
  NOR2_X1 U423 ( .A1(n361), .A2(n359), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n360), .B(KEYINPUT25), .ZN(n365) );
  INV_X1 U425 ( .A(n361), .ZN(n465) );
  NOR2_X1 U426 ( .A1(n527), .A2(n465), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n362), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U428 ( .A1(n363), .A2(n566), .ZN(n364) );
  NAND2_X1 U429 ( .A1(n365), .A2(n364), .ZN(n367) );
  NAND2_X1 U430 ( .A1(n367), .A2(n366), .ZN(n368) );
  XOR2_X1 U431 ( .A(KEYINPUT96), .B(n368), .Z(n369) );
  NOR2_X1 U432 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n371), .B(KEYINPUT97), .ZN(n477) );
  XOR2_X1 U434 ( .A(G183GAT), .B(G211GAT), .Z(n373) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G57GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U437 ( .A(n374), .B(G78GAT), .Z(n376) );
  XOR2_X1 U438 ( .A(G71GAT), .B(KEYINPUT13), .Z(n415) );
  XNOR2_X1 U439 ( .A(G155GAT), .B(n415), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n381) );
  XNOR2_X1 U441 ( .A(G22GAT), .B(G15GAT), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n377), .B(KEYINPUT69), .ZN(n434) );
  XOR2_X1 U443 ( .A(n434), .B(KEYINPUT12), .Z(n379) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U446 ( .A(n381), .B(n380), .Z(n389) );
  XOR2_X1 U447 ( .A(KEYINPUT77), .B(G8GAT), .Z(n383) );
  XNOR2_X1 U448 ( .A(G1GAT), .B(G64GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U450 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n385) );
  XNOR2_X1 U451 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n576) );
  NAND2_X1 U455 ( .A1(n477), .A2(n576), .ZN(n409) );
  XNOR2_X1 U456 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n390), .B(G36GAT), .ZN(n391) );
  XOR2_X1 U458 ( .A(n391), .B(KEYINPUT8), .Z(n393) );
  XNOR2_X1 U459 ( .A(G50GAT), .B(KEYINPUT68), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n433) );
  XOR2_X1 U461 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n395) );
  XNOR2_X1 U462 ( .A(G106GAT), .B(G92GAT), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n433), .B(n396), .ZN(n408) );
  XOR2_X1 U465 ( .A(KEYINPUT11), .B(G218GAT), .Z(n398) );
  XNOR2_X1 U466 ( .A(G162GAT), .B(G29GAT), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U468 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U469 ( .A1(G232GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U471 ( .A(n403), .B(KEYINPUT75), .Z(n406) );
  XNOR2_X1 U472 ( .A(G85GAT), .B(KEYINPUT72), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n404), .B(G99GAT), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n411), .B(KEYINPUT10), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n554) );
  XNOR2_X1 U477 ( .A(KEYINPUT36), .B(n554), .ZN(n580) );
  NOR2_X1 U478 ( .A1(n409), .A2(n580), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n410), .B(KEYINPUT37), .ZN(n514) );
  XNOR2_X1 U480 ( .A(n411), .B(KEYINPUT73), .ZN(n413) );
  AND2_X1 U481 ( .A1(G230GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U482 ( .A(n413), .B(n412), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n418) );
  INV_X1 U484 ( .A(G204GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n429) );
  XNOR2_X1 U486 ( .A(G148GAT), .B(n423), .ZN(n427) );
  XOR2_X1 U487 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n425) );
  XNOR2_X1 U488 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U490 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n431) );
  XNOR2_X1 U491 ( .A(G197GAT), .B(KEYINPUT30), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n443) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U497 ( .A(n438), .B(KEYINPUT65), .Z(n441) );
  XNOR2_X1 U498 ( .A(n439), .B(KEYINPUT67), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n501) );
  XNOR2_X1 U501 ( .A(n501), .B(KEYINPUT70), .ZN(n556) );
  NAND2_X1 U502 ( .A1(n572), .A2(n556), .ZN(n444) );
  XNOR2_X1 U503 ( .A(KEYINPUT74), .B(n444), .ZN(n480) );
  NOR2_X1 U504 ( .A1(n514), .A2(n480), .ZN(n445) );
  NAND2_X1 U505 ( .A1(n499), .A2(n527), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n447) );
  XOR2_X1 U507 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n467) );
  NAND2_X1 U508 ( .A1(n554), .A2(n576), .ZN(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n452) );
  INV_X1 U510 ( .A(KEYINPUT41), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n450), .B(n572), .ZN(n546) );
  NAND2_X1 U512 ( .A1(n501), .A2(n559), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U514 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n455), .B(KEYINPUT47), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n576), .A2(n580), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT45), .B(n456), .Z(n457) );
  NOR2_X1 U518 ( .A1(n556), .A2(n457), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n458), .A2(n572), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT64), .B(KEYINPUT48), .Z(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n524) );
  NOR2_X1 U523 ( .A1(n483), .A2(n524), .ZN(n463) );
  XOR2_X1 U524 ( .A(n463), .B(KEYINPUT54), .Z(n464) );
  NAND2_X1 U525 ( .A1(n567), .A2(n465), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n468) );
  INV_X1 U527 ( .A(n554), .ZN(n537) );
  NAND2_X1 U528 ( .A1(n563), .A2(n537), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n471) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT99), .B(n475), .Z(n482) );
  NOR2_X1 U533 ( .A1(n576), .A2(n537), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT16), .B(n476), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n479), .B(KEYINPUT98), .ZN(n503) );
  NOR2_X1 U537 ( .A1(n480), .A2(n503), .ZN(n490) );
  NAND2_X1 U538 ( .A1(n490), .A2(n516), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1324GAT) );
  XOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT101), .Z(n485) );
  INV_X1 U541 ( .A(n483), .ZN(n518) );
  NAND2_X1 U542 ( .A1(n490), .A2(n518), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n487) );
  NAND2_X1 U545 ( .A1(n490), .A2(n527), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n489) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT102), .Z(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n492) );
  NAND2_X1 U550 ( .A1(n490), .A2(n529), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT106), .Z(n495) );
  NAND2_X1 U554 ( .A1(n499), .A2(n516), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n497) );
  XOR2_X1 U556 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n518), .A2(n499), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n529), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT109), .Z(n505) );
  INV_X1 U563 ( .A(n501), .ZN(n568) );
  NAND2_X1 U564 ( .A1(n568), .A2(n559), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT110), .ZN(n515) );
  NOR2_X1 U566 ( .A1(n503), .A2(n515), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n511), .A2(n516), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT111), .Z(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n518), .A2(n511), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(KEYINPUT112), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n527), .A2(n511), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U577 ( .A1(n511), .A2(n529), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n521), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n527), .A2(n521), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n529), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT114), .ZN(n543) );
  NAND2_X1 U591 ( .A1(n527), .A2(n543), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n538), .A2(n556), .ZN(n531) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT115), .Z(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n533) );
  NAND2_X1 U597 ( .A1(n538), .A2(n559), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  INV_X1 U600 ( .A(n576), .ZN(n564) );
  NAND2_X1 U601 ( .A1(n564), .A2(n538), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT117), .Z(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n566), .A2(n543), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n568), .A2(n553), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n553), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(KEYINPUT52), .B(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n576), .A2(n553), .ZN(n552) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n563), .ZN(n557) );
  XOR2_X1 U624 ( .A(n557), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  NAND2_X1 U627 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n568), .A2(n579), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n579), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n577), .Z(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

