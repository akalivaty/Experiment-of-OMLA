//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT66), .Z(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT65), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n209), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n212), .B1(new_n215), .B2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G13), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n214), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G250), .B1(G257), .B2(G264), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n222), .B2(KEYINPUT0), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT67), .Z(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n215), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n223), .B(new_n231), .C1(KEYINPUT0), .C2(new_n222), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n208), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  INV_X1    g0054(.A(G58), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n209), .A2(G33), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n251), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n250), .B1(new_n213), .B2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(G50), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G274), .ZN(new_n274));
  INV_X1    g0074(.A(new_n273), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  OAI211_X1 g0076(.A(G1), .B(G13), .C1(new_n276), .C2(new_n271), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1698), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n284), .A2(G222), .B1(new_n287), .B2(G77), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n282), .B2(new_n283), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n288), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n280), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n269), .A2(new_n270), .B1(G190), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT10), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(new_n268), .B2(KEYINPUT9), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n300), .B1(new_n296), .B2(new_n301), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n257), .A2(new_n263), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n257), .B2(new_n266), .ZN(new_n306));
  INV_X1    g0106(.A(G68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n282), .A2(new_n209), .A3(new_n283), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n283), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n255), .A2(new_n307), .ZN(new_n313));
  OAI21_X1  g0113(.A(G20), .B1(new_n313), .B2(new_n202), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n260), .A2(G159), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT16), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n287), .B2(new_n209), .ZN(new_n318));
  INV_X1    g0118(.A(new_n311), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT16), .ZN(new_n321));
  INV_X1    g0121(.A(new_n316), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n306), .B1(new_n324), .B2(new_n250), .ZN(new_n325));
  OAI211_X1 g0125(.A(G223), .B(new_n290), .C1(new_n285), .C2(new_n286), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n282), .A2(new_n283), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n329), .A2(KEYINPUT78), .A3(G223), .A4(new_n290), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n291), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n277), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n274), .B1(new_n278), .B2(new_n236), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n297), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  INV_X1    g0136(.A(new_n334), .ZN(new_n337));
  OAI211_X1 g0137(.A(G226), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n338));
  INV_X1    g0138(.A(G87), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n276), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n328), .B2(new_n330), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n336), .B(new_n337), .C1(new_n341), .C2(new_n277), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n325), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n347));
  OAI211_X1 g0147(.A(G179), .B(new_n337), .C1(new_n341), .C2(new_n277), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT18), .B1(new_n349), .B2(new_n325), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n312), .A2(KEYINPUT16), .A3(new_n316), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n250), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n306), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT18), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(new_n348), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n325), .A2(new_n343), .A3(KEYINPUT17), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n346), .A2(new_n350), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n269), .B1(G169), .B2(new_n295), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G179), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n362), .A2(new_n363), .B1(new_n365), .B2(new_n295), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n284), .A2(G232), .B1(new_n287), .B2(G107), .ZN(new_n368));
  INV_X1    g0168(.A(G238), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n292), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n294), .ZN(new_n371));
  INV_X1    g0171(.A(G244), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n274), .C1(new_n372), .C2(new_n278), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n297), .B2(new_n373), .ZN(new_n375));
  INV_X1    g0175(.A(new_n260), .ZN(new_n376));
  INV_X1    g0176(.A(G77), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n252), .A2(new_n376), .B1(new_n209), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT70), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n378), .A2(new_n379), .B1(new_n258), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n250), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n266), .A2(new_n377), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n263), .B2(new_n377), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n373), .A2(G169), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n365), .B2(new_n373), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n387), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n304), .A2(new_n361), .A3(new_n367), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(KEYINPUT76), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n274), .B1(new_n278), .B2(new_n369), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n284), .A2(KEYINPUT73), .A3(G226), .ZN(new_n399));
  OAI211_X1 g0199(.A(G226), .B(new_n290), .C1(new_n285), .C2(new_n286), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT73), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G97), .ZN(new_n403));
  OAI211_X1 g0203(.A(G232), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n399), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n398), .B1(new_n405), .B2(new_n294), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n403), .B(new_n404), .C1(new_n400), .C2(new_n401), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT73), .B1(new_n284), .B2(G226), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n294), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n398), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT74), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n415), .A3(new_n407), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n408), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G169), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n397), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n411), .A2(new_n412), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n406), .B2(new_n407), .ZN(new_n422));
  AND4_X1   g0222(.A1(new_n415), .A2(new_n411), .A3(new_n407), .A4(new_n412), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(G169), .A3(new_n396), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(G179), .A3(new_n413), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n217), .A2(G1), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G20), .A3(new_n307), .ZN(new_n433));
  XOR2_X1   g0233(.A(new_n433), .B(KEYINPUT12), .Z(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(G68), .B2(new_n263), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n376), .A2(new_n264), .B1(new_n209), .B2(G68), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n258), .A2(new_n377), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n250), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n439));
  XNOR2_X1  g0239(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n431), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n408), .A2(new_n336), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n443), .B2(new_n413), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n297), .B2(new_n417), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n394), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n329), .A2(G250), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n290), .B1(new_n448), .B2(KEYINPUT4), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT4), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(G244), .C1(new_n286), .C2(new_n285), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n372), .B1(new_n282), .B2(new_n283), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(KEYINPUT4), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n294), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n272), .A2(G1), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  AND2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(G274), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n458), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n277), .ZN(new_n462));
  INV_X1    g0262(.A(G257), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(G190), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n260), .A2(G77), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n472), .A2(KEYINPUT6), .A3(G97), .ZN(new_n473));
  XNOR2_X1  g0273(.A(G97), .B(G107), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT6), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n471), .B1(new_n476), .B2(new_n209), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n472), .B1(new_n310), .B2(new_n311), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n250), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n480));
  OAI21_X1  g0280(.A(G107), .B1(new_n318), .B2(new_n319), .ZN(new_n481));
  AND2_X1   g0281(.A1(G97), .A2(G107), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G97), .A2(G107), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n475), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n472), .A2(KEYINPUT6), .A3(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n250), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n266), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n213), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n266), .A2(new_n493), .A3(new_n208), .A4(new_n249), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G97), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n480), .A2(new_n490), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n466), .A2(G200), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n470), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G250), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n282), .B2(new_n283), .ZN(new_n504));
  OAI21_X1  g0304(.A(G1698), .B1(new_n504), .B2(new_n450), .ZN(new_n505));
  OAI21_X1  g0305(.A(G244), .B1(new_n285), .B2(new_n286), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n450), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n505), .A2(new_n452), .A3(new_n507), .A4(new_n453), .ZN(new_n508));
  AOI211_X1 g0308(.A(KEYINPUT81), .B(new_n464), .C1(new_n508), .C2(new_n294), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n468), .B1(new_n456), .B2(new_n465), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n418), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n499), .A2(new_n492), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n489), .B1(new_n488), .B2(new_n250), .ZN(new_n513));
  AOI211_X1 g0313(.A(KEYINPUT79), .B(new_n251), .C1(new_n481), .C2(new_n487), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n456), .A2(new_n365), .A3(new_n465), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n502), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(G250), .B1(new_n272), .B2(G1), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n457), .A2(G274), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n294), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G238), .B(new_n290), .C1(new_n285), .C2(new_n286), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n506), .C2(new_n290), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n336), .B(new_n523), .C1(new_n526), .C2(new_n294), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n526), .B2(new_n294), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n527), .B1(G200), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT19), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n209), .B1(new_n403), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n339), .A2(new_n491), .A3(new_n472), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n209), .B(G68), .C1(new_n285), .C2(new_n286), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n531), .B1(new_n403), .B2(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n266), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n537), .A2(new_n250), .B1(new_n538), .B2(new_n380), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n496), .A2(G87), .A3(new_n497), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n380), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n496), .A2(new_n542), .A3(new_n497), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n539), .A2(new_n543), .B1(new_n528), .B2(new_n365), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n528), .A2(G169), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n530), .A2(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n502), .A2(new_n517), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(KEYINPUT82), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n276), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(new_n551), .B2(new_n453), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n209), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n250), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(KEYINPUT20), .B(new_n250), .C1(new_n552), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n494), .A2(G116), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G116), .B2(new_n538), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n418), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G270), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n460), .B1(new_n462), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G264), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n566));
  OAI211_X1 g0366(.A(G257), .B(new_n290), .C1(new_n285), .C2(new_n286), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(new_n294), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n569), .B2(new_n294), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n562), .A2(new_n573), .A3(KEYINPUT21), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT21), .B1(new_n562), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT84), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n559), .A2(new_n561), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G179), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n572), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n569), .A2(new_n570), .A3(new_n294), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n564), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT84), .A3(G179), .A4(new_n578), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n336), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n584), .B2(G200), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n579), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n576), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT87), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n496), .A2(G107), .A3(new_n497), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n432), .A2(G20), .A3(new_n472), .ZN(new_n593));
  XOR2_X1   g0393(.A(new_n593), .B(KEYINPUT25), .Z(new_n594));
  AND2_X1   g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n553), .B2(new_n258), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT23), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(new_n472), .A3(G20), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(KEYINPUT85), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(KEYINPUT85), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n209), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n603), .A2(KEYINPUT22), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(KEYINPUT22), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n602), .B(KEYINPUT24), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n250), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n603), .B(KEYINPUT22), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT24), .B1(new_n608), .B2(new_n602), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n595), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(G33), .A2(G294), .ZN(new_n611));
  OAI211_X1 g0411(.A(G257), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n612));
  OAI211_X1 g0412(.A(G250), .B(new_n290), .C1(new_n285), .C2(new_n286), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT86), .B1(new_n504), .B2(new_n290), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n294), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n462), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G264), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n460), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G169), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n620), .A2(new_n365), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n610), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n617), .A2(new_n619), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n336), .A3(new_n460), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n297), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n591), .B(new_n624), .C1(new_n628), .C2(new_n610), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n610), .B1(new_n627), .B2(new_n626), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(G179), .A3(new_n460), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT24), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n250), .A3(new_n606), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n631), .A2(new_n621), .B1(new_n635), .B2(new_n595), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT87), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n590), .B1(new_n629), .B2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n447), .A2(new_n520), .A3(new_n550), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n545), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT88), .B1(new_n528), .B2(G169), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n544), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n527), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n645), .B(new_n541), .C1(new_n297), .C2(new_n528), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n549), .A2(new_n630), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n576), .A2(new_n586), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n636), .A2(KEYINPUT89), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n624), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n644), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n516), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n480), .A2(new_n490), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n512), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n547), .A2(new_n657), .A3(new_n511), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n658), .A2(KEYINPUT90), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT90), .B1(new_n658), .B2(new_n659), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n657), .A2(new_n511), .A3(new_n646), .A4(new_n643), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n447), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n349), .A2(new_n325), .A3(KEYINPUT18), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT91), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n350), .A2(new_n670), .A3(new_n358), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n431), .A2(new_n441), .B1(new_n445), .B2(new_n392), .ZN(new_n673));
  INV_X1    g0473(.A(new_n359), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT17), .B1(new_n325), .B2(new_n343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n672), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n678), .A2(new_n304), .B1(new_n364), .B2(new_n366), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n666), .A2(new_n679), .ZN(G369));
  INV_X1    g0480(.A(new_n432), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .A3(G20), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT27), .B1(new_n681), .B2(G20), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n578), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n576), .B2(new_n586), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n576), .A2(new_n586), .A3(new_n589), .A4(new_n687), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g0492(.A(G330), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n629), .A2(new_n637), .B1(new_n610), .B2(new_n686), .ZN(new_n694));
  INV_X1    g0494(.A(new_n686), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n624), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n649), .A2(new_n686), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n652), .A2(new_n650), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n694), .A2(new_n700), .B1(new_n701), .B2(new_n695), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n220), .A2(G41), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n213), .ZN(new_n705));
  NOR4_X1   g0505(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(new_n207), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT26), .B1(new_n517), .B2(new_n647), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n547), .A2(new_n657), .A3(new_n659), .A4(new_n511), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(KEYINPUT95), .A3(new_n643), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n630), .A2(new_n647), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n576), .A2(new_n624), .A3(new_n586), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n518), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n644), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT95), .B1(new_n716), .B2(new_n710), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT29), .B(new_n695), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n686), .B1(new_n654), .B2(new_n664), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT29), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n638), .A2(new_n550), .A3(new_n520), .A4(new_n695), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n509), .A2(new_n510), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n625), .A2(new_n528), .ZN(new_n723));
  INV_X1    g0523(.A(new_n580), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT30), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n466), .A2(new_n620), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  NAND3_X1  g0530(.A1(new_n573), .A2(new_n365), .A3(new_n529), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n727), .B(new_n728), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n686), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n736));
  OAI211_X1 g0536(.A(new_n721), .B(new_n735), .C1(new_n733), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n720), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n708), .B1(new_n740), .B2(G1), .ZN(G364));
  INV_X1    g0541(.A(new_n693), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n217), .A2(G20), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G45), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n705), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n690), .A2(new_n692), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(G330), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n745), .B(KEYINPUT96), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(G1), .B(G13), .C1(new_n209), .C2(G169), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT99), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT99), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(G20), .A2(G190), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n365), .A3(new_n297), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n336), .A2(G20), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT32), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n329), .B1(new_n759), .B2(new_n264), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n365), .A2(new_n297), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n209), .B1(new_n762), .B2(G190), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n307), .B1(new_n771), .B2(new_n491), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT100), .ZN(new_n773));
  INV_X1    g0573(.A(new_n757), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G179), .A3(new_n297), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n760), .A2(new_n365), .A3(G200), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n776), .A2(G58), .B1(new_n777), .B2(G77), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n760), .A2(G179), .A3(new_n297), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n472), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n757), .A2(new_n297), .A3(G179), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G87), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n768), .A2(new_n773), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n759), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n777), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT33), .B(G317), .Z(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n788), .B1(new_n770), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n786), .B(new_n790), .C1(G322), .C2(new_n776), .ZN(new_n791));
  INV_X1    g0591(.A(new_n771), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G294), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n329), .B1(new_n779), .B2(G283), .ZN(new_n794));
  INV_X1    g0594(.A(new_n763), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G329), .B1(G303), .B2(new_n782), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n791), .A2(new_n793), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n756), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT97), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n209), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT98), .Z(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n756), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n220), .A2(new_n329), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n244), .A2(new_n272), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n207), .A2(G45), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n219), .A2(G355), .A3(new_n329), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n553), .B2(new_n220), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n804), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n751), .A2(new_n798), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n748), .B2(new_n803), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n749), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  AOI21_X1  g0615(.A(new_n695), .B1(new_n384), .B2(new_n386), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n391), .B1(new_n388), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n392), .A2(new_n695), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n719), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n719), .A2(new_n819), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n745), .B1(new_n825), .B2(new_n738), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(KEYINPUT103), .B1(new_n738), .B2(new_n825), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT103), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n745), .C1(new_n825), .C2(new_n738), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n777), .A2(G159), .B1(new_n758), .B2(G137), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n775), .C1(new_n833), .C2(new_n770), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n782), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n329), .B1(new_n838), .B2(new_n264), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n780), .A2(new_n307), .B1(new_n763), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G58), .C2(new_n792), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n836), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n287), .B1(new_n838), .B2(new_n472), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT101), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n795), .A2(G311), .B1(new_n779), .B2(G87), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n777), .A2(G116), .B1(new_n758), .B2(G303), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n770), .A2(new_n848), .B1(new_n775), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G97), .B2(new_n792), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n756), .B1(new_n843), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n755), .A2(new_n799), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n853), .B(new_n751), .C1(new_n377), .C2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n819), .B2(new_n800), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n830), .A2(new_n856), .ZN(G384));
  OAI211_X1 g0657(.A(G116), .B(new_n210), .C1(new_n486), .C2(KEYINPUT35), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(KEYINPUT35), .B2(new_n486), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n207), .B(G77), .C1(new_n255), .C2(new_n307), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n201), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n213), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n822), .A2(new_n818), .ZN(new_n865));
  INV_X1    g0665(.A(new_n441), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n695), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n442), .A2(KEYINPUT104), .A3(new_n445), .A4(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n419), .A2(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n869));
  OAI211_X1 g0669(.A(KEYINPUT104), .B(new_n445), .C1(new_n869), .C2(new_n866), .ZN(new_n870));
  INV_X1    g0670(.A(new_n867), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n355), .A2(new_n357), .ZN(new_n876));
  INV_X1    g0676(.A(new_n684), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n251), .B1(new_n317), .B2(new_n323), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n306), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n344), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n876), .A2(new_n344), .A3(new_n882), .A4(new_n879), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n879), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n360), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n875), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n886), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(KEYINPUT105), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n874), .A2(new_n896), .B1(new_n672), .B2(new_n877), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n892), .B2(new_n893), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n669), .A2(new_n676), .A3(new_n671), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(new_n885), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n884), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n901), .B2(new_n885), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n891), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT107), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT107), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(new_n891), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n893), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n900), .B1(new_n910), .B2(KEYINPUT39), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n442), .A2(new_n686), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n897), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n447), .B(new_n718), .C1(KEYINPUT29), .C2(new_n719), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n679), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n736), .B1(new_n732), .B2(new_n686), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n721), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n733), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n734), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n868), .A2(new_n872), .A3(new_n819), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n721), .A2(new_n917), .B1(new_n919), .B2(new_n734), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n868), .A2(new_n872), .A3(new_n819), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n895), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n910), .A2(new_n924), .B1(new_n927), .B2(new_n923), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n447), .A2(new_n925), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT108), .Z(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n916), .A2(new_n933), .B1(new_n213), .B2(new_n743), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n916), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n864), .B1(new_n934), .B2(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n694), .A2(new_n700), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n518), .B1(new_n500), .B2(new_n695), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n937), .A2(KEYINPUT42), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT42), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n517), .B1(new_n938), .B2(new_n624), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n695), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT43), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n695), .A2(new_n541), .ZN(new_n945));
  MUX2_X1   g0745(.A(new_n647), .B(new_n643), .S(new_n945), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n944), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n657), .A2(new_n511), .A3(new_n686), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n938), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n698), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n704), .B(new_n954), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n693), .A2(new_n697), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n957), .A2(new_n698), .B1(new_n649), .B2(new_n686), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n699), .A2(new_n700), .A3(new_n956), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n958), .A2(new_n959), .A3(new_n720), .A4(new_n738), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n701), .A2(new_n695), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n937), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n951), .ZN(new_n964));
  NOR2_X1   g0764(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n702), .B2(new_n951), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n702), .A2(new_n951), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(new_n974), .C1(KEYINPUT111), .C2(new_n699), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n699), .A2(KEYINPUT111), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n972), .B(KEYINPUT45), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n966), .A2(new_n968), .B1(KEYINPUT110), .B2(KEYINPUT44), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n961), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT112), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n961), .A2(new_n975), .A3(new_n982), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n955), .B1(new_n984), .B2(new_n740), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n744), .A2(G1), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n953), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n803), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n946), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n805), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n990), .A2(new_n240), .B1(new_n219), .B2(new_n380), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n750), .B1(new_n804), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n329), .B1(new_n838), .B2(new_n255), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n780), .A2(new_n377), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G137), .C2(new_n795), .ZN(new_n996));
  INV_X1    g0796(.A(new_n770), .ZN(new_n997));
  INV_X1    g0797(.A(new_n201), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n997), .A2(G159), .B1(new_n998), .B2(new_n777), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n776), .A2(G150), .B1(new_n758), .B2(G143), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n771), .A2(new_n307), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n782), .A2(G116), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT113), .Z(new_n1007));
  OAI22_X1  g0807(.A1(new_n780), .A2(new_n491), .B1(new_n787), .B2(new_n848), .ZN(new_n1008));
  INV_X1    g0808(.A(G303), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n287), .B1(new_n775), .B2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1004), .A2(new_n1005), .B1(new_n472), .B2(new_n771), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n997), .A2(G294), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n795), .A2(G317), .B1(new_n758), .B2(G311), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1007), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT47), .B1(new_n1003), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1003), .A2(KEYINPUT47), .A3(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n755), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n989), .B(new_n993), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n987), .A2(new_n1019), .ZN(G387));
  AOI22_X1  g0820(.A1(new_n792), .A2(G283), .B1(G294), .B2(new_n782), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n777), .A2(G303), .B1(new_n758), .B2(G322), .ZN(new_n1022));
  INV_X1    g0822(.A(G317), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1022), .B1(new_n788), .B2(new_n770), .C1(new_n1023), .C2(new_n775), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT115), .Z(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT49), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n287), .B1(new_n763), .B2(new_n785), .C1(new_n780), .C2(new_n553), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT116), .Z(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n838), .A2(new_n377), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G159), .B2(new_n758), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n287), .B1(new_n779), .B2(G97), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n795), .A2(G150), .B1(new_n777), .B2(G68), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n771), .A2(new_n380), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G50), .B2(new_n776), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT114), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n257), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1038), .B(new_n1041), .C1(new_n1042), .C2(new_n997), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n755), .B1(new_n1033), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n237), .A2(G45), .A3(new_n287), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n252), .A2(G50), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT50), .Z(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n1047), .C1(G68), .C2(G77), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n706), .B1(new_n1048), .B2(new_n329), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n219), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n804), .B1(G107), .B2(new_n220), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n751), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n697), .B2(new_n988), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n958), .A2(new_n959), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1055), .B1(new_n1057), .B2(new_n986), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n739), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(new_n704), .A3(new_n960), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT117), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1058), .A2(new_n1063), .A3(new_n1060), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(G393));
  AOI22_X1  g0865(.A1(new_n776), .A2(G159), .B1(new_n758), .B2(G150), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n838), .A2(new_n307), .B1(new_n763), .B2(new_n832), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n787), .A2(new_n252), .B1(new_n201), .B2(new_n770), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n771), .A2(new_n377), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n329), .C1(new_n339), .C2(new_n780), .ZN(new_n1072));
  OR4_X1    g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n329), .B(new_n781), .C1(G116), .C2(new_n792), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n759), .A2(new_n1023), .B1(new_n775), .B2(new_n788), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G303), .A2(new_n997), .B1(new_n795), .B2(G322), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n777), .A2(G294), .B1(new_n782), .B2(G283), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n756), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n990), .A2(new_n247), .B1(new_n491), .B2(new_n219), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n804), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n751), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n951), .B2(new_n803), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n971), .A2(new_n974), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(new_n698), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n986), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n704), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1086), .B2(new_n960), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n984), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(G390));
  INV_X1    g0892(.A(new_n854), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n750), .B1(new_n1042), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n782), .A2(G150), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT53), .Z(new_n1096));
  AOI22_X1  g0896(.A1(new_n997), .A2(G137), .B1(new_n998), .B2(new_n779), .ZN(new_n1097));
  INV_X1    g0897(.A(G125), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(new_n763), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n287), .B1(new_n776), .B2(G132), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT54), .B(G143), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n777), .B1(G128), .B2(new_n758), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1100), .B(new_n1103), .C1(new_n764), .C2(new_n771), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n287), .B1(new_n838), .B2(new_n339), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT119), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n795), .A2(G294), .B1(new_n776), .B2(G116), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n997), .A2(G107), .B1(new_n758), .B2(G283), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G68), .A2(new_n779), .B1(new_n777), .B2(G97), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1071), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1099), .A2(new_n1104), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1094), .B1(new_n1111), .B2(new_n755), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n911), .B2(new_n800), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n912), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n719), .A2(new_n817), .B1(new_n392), .B2(new_n695), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n873), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1117), .B(new_n900), .C1(new_n910), .C2(KEYINPUT39), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n737), .A2(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n926), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n695), .B(new_n817), .C1(new_n715), .C2(new_n717), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n818), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n912), .B1(new_n1122), .B2(new_n873), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT118), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n909), .A2(new_n893), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n901), .A2(new_n885), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT106), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n884), .A3(new_n903), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n908), .B1(new_n1128), .B2(new_n891), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1123), .B(new_n1124), .C1(new_n1125), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1124), .B1(new_n910), .B2(new_n1123), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1118), .B(new_n1120), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n899), .B1(new_n1134), .B2(new_n898), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1123), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT118), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1135), .A2(new_n1117), .B1(new_n1137), .B2(new_n1130), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n925), .A2(G330), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(new_n922), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1113), .B1(new_n1142), .B2(new_n1087), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n930), .A2(G330), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n679), .A3(new_n914), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n873), .B1(new_n1119), .B2(new_n819), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n865), .B1(new_n1146), .B2(new_n1140), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n925), .A2(G330), .A3(new_n819), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1116), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1120), .A2(new_n1149), .A3(new_n818), .A4(new_n1121), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1145), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1133), .B(new_n1151), .C1(new_n1138), .C2(new_n1141), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1089), .B1(new_n1142), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1143), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(G378));
  NOR2_X1   g0956(.A1(new_n672), .A2(new_n877), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n895), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1135), .B2(new_n1114), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n304), .A2(new_n367), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n269), .A3(new_n877), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n304), .B(new_n367), .C1(new_n268), .C2(new_n684), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n928), .B2(G330), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n924), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n927), .A2(new_n923), .ZN(new_n1169));
  AND4_X1   g0969(.A1(G330), .A2(new_n1168), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1160), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(G330), .A3(new_n1169), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1166), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n928), .A2(G330), .A3(new_n1166), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n913), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n801), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n746), .B1(new_n1093), .B2(new_n998), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n759), .A2(new_n1098), .B1(new_n770), .B2(new_n840), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n776), .A2(G128), .B1(new_n1102), .B2(new_n782), .ZN(new_n1181));
  INV_X1    g0981(.A(G137), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n787), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1180), .B(new_n1183), .C1(G150), .C2(new_n792), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n276), .B(new_n271), .C1(new_n780), .C2(new_n764), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G124), .B2(new_n795), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n775), .A2(new_n472), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n542), .A2(new_n777), .B1(G116), .B2(new_n758), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n848), .C2(new_n763), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n287), .A2(new_n271), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1034), .A2(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n780), .A2(new_n255), .B1(new_n491), .B2(new_n770), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1194), .A2(new_n1001), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT58), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(KEYINPUT58), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1195), .B(new_n264), .C1(G33), .C2(G41), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1190), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1179), .B1(new_n1202), .B2(new_n755), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1177), .A2(new_n986), .B1(new_n1178), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1145), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1152), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT121), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1206), .A2(new_n1208), .A3(KEYINPUT121), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1152), .A2(new_n1205), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n704), .B1(new_n1214), .B2(KEYINPUT57), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1204), .B1(new_n1213), .B2(new_n1215), .ZN(G375));
  INV_X1    g1016(.A(new_n955), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1147), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1153), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n986), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n759), .A2(new_n840), .B1(new_n775), .B2(new_n1182), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n329), .B1(new_n780), .B2(new_n255), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G50), .C2(new_n792), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n787), .A2(new_n833), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n838), .A2(new_n764), .B1(new_n770), .B2(new_n1101), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(G128), .C2(new_n795), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n787), .A2(new_n472), .B1(new_n759), .B2(new_n849), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n838), .A2(new_n491), .B1(new_n763), .B2(new_n1009), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n770), .A2(new_n553), .B1(new_n775), .B2(new_n848), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n995), .A2(new_n1231), .A3(new_n329), .A4(new_n1039), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1224), .A2(new_n1227), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n750), .B1(G68), .B2(new_n1093), .C1(new_n1233), .C2(new_n756), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1116), .B2(new_n799), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1219), .A2(new_n1221), .A3(new_n1236), .ZN(G381));
  INV_X1    g1037(.A(new_n1204), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1206), .A2(KEYINPUT121), .A3(new_n1208), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT121), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1206), .A2(new_n1177), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1089), .B1(new_n1242), .B2(new_n1207), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1238), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1155), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n856), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n827), .B2(new_n829), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1091), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1062), .A2(new_n814), .A3(new_n1064), .ZN(new_n1249));
  OR2_X1    g1049(.A1(G381), .A2(new_n1249), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G387), .A2(new_n1245), .A3(new_n1248), .A4(new_n1250), .ZN(G407));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND3_X1  g1052(.A1(new_n987), .A2(new_n1019), .A3(G390), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1058), .A2(new_n1063), .A3(new_n1060), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1063), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1257));
  OAI21_X1  g1057(.A(G396), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1258), .A2(new_n1249), .A3(KEYINPUT124), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT124), .B1(new_n1258), .B2(new_n1249), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1253), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n987), .B2(new_n1019), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1255), .B(new_n1261), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1253), .C1(new_n1254), .C2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT122), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1089), .B(new_n1151), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1221), .A2(new_n1236), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1247), .B(new_n1270), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1151), .A2(new_n1089), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT122), .B1(new_n1278), .B2(G384), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(G384), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G2897), .ZN(new_n1282));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1282), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1275), .A2(new_n1279), .A3(new_n1280), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1204), .B1(new_n1242), .B2(new_n955), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1155), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1244), .B2(G378), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1293), .B2(new_n1284), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G378), .B(new_n1204), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1291), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1281), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1285), .A4(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1294), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1284), .B(new_n1281), .C1(new_n1295), .C2(new_n1291), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1302), .A2(new_n1297), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1269), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1268), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1296), .A2(new_n1285), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n1289), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT123), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1302), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  OAI211_X1 g1111(.A(KEYINPUT123), .B(new_n1311), .C1(new_n1307), .C2(new_n1281), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1308), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1304), .A2(new_n1313), .ZN(G405));
  NAND2_X1  g1114(.A1(G375), .A2(G378), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1269), .A2(new_n1245), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1245), .A2(new_n1315), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1268), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1316), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


