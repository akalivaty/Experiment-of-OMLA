//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G250), .B1(G257), .B2(G264), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT66), .B(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n215), .A2(KEYINPUT0), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT67), .B(G238), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n222), .A2(G68), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G87), .A2(G250), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n221), .B1(KEYINPUT0), .B2(new_n215), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G107), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n245), .B(new_n250), .Z(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n217), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n254), .B2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G20), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n204), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT8), .B(G58), .Z(new_n265));
  NAND2_X1  g0065(.A1(new_n216), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n253), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n256), .B1(G50), .B2(new_n259), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(KEYINPUT70), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n205), .ZN(new_n285));
  MUX2_X1   g0085(.A(G222), .B(G223), .S(G1698), .Z(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n274), .B1(new_n287), .B2(KEYINPUT71), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(KEYINPUT71), .B2(new_n287), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n274), .A2(G274), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n274), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G226), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT69), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n289), .A2(G190), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n289), .A2(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n271), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n271), .A2(new_n304), .A3(new_n299), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n270), .B1(new_n300), .B2(G179), .ZN(new_n307));
  AOI21_X1  g0107(.A(G169), .B1(new_n289), .B2(new_n298), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n293), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n295), .B2(KEYINPUT74), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n314));
  OR3_X1    g0114(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n292), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G226), .A2(G1698), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n235), .B2(G1698), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n278), .A2(new_n318), .A3(new_n283), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n314), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT13), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n316), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(G190), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT11), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n263), .A2(new_n247), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n266), .A2(new_n205), .B1(new_n260), .B2(G68), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT76), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI221_X1 g0135(.A(KEYINPUT76), .B1(new_n260), .B2(G68), .C1(new_n266), .C2(new_n205), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n331), .B1(new_n337), .B2(new_n269), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT12), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n259), .B2(G68), .ZN(new_n340));
  INV_X1    g0140(.A(new_n259), .ZN(new_n341));
  INV_X1    g0141(.A(G68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(KEYINPUT12), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n255), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n340), .B(new_n343), .C1(new_n344), .C2(new_n342), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n269), .B1(new_n335), .B2(new_n336), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(KEYINPUT11), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n330), .A2(new_n338), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n329), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n328), .B1(new_n316), .B2(new_n325), .ZN(new_n350));
  OAI21_X1  g0150(.A(G200), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n327), .A2(new_n329), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT75), .A3(G200), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n348), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n338), .A2(new_n347), .ZN(new_n357));
  OAI21_X1  g0157(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n327), .A2(G179), .A3(new_n329), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT14), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n361), .A3(G169), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n356), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n284), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n222), .A2(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n365), .B(new_n366), .C1(new_n235), .C2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n314), .C1(G107), .C2(new_n365), .ZN(new_n368));
  INV_X1    g0168(.A(new_n295), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n311), .B1(G244), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G190), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n265), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n376), .B1(new_n205), .B2(new_n216), .C1(new_n263), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT72), .B1(new_n267), .B2(new_n375), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n253), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n259), .A2(G77), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n255), .B2(G77), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n371), .A2(G200), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n373), .A2(new_n380), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n382), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n386), .B(new_n387), .C1(G179), .C2(new_n371), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n306), .A2(new_n310), .A3(new_n364), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT78), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n260), .B1(new_n203), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n262), .A2(G159), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n392), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n202), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT78), .A3(new_n394), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT66), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G20), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n281), .A2(new_n403), .A3(new_n405), .A4(new_n282), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n276), .A2(new_n277), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(G20), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n402), .B1(new_n412), .B2(G68), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n406), .A2(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n414), .A2(KEYINPUT77), .A3(new_n342), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n401), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT7), .A2(G20), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n278), .B2(new_n283), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n407), .B1(new_n409), .B2(new_n216), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n420), .A2(new_n421), .A3(new_n342), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n393), .A2(new_n395), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n416), .A2(new_n425), .A3(new_n253), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n377), .A2(new_n341), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n344), .B2(new_n377), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n296), .A2(G1698), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n430), .B1(G223), .B2(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n274), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n293), .B1(new_n295), .B2(new_n235), .ZN(new_n434));
  OAI21_X1  g0234(.A(G200), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n434), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n432), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n314), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n426), .A2(new_n429), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT77), .B1(new_n414), .B2(new_n342), .ZN(new_n446));
  INV_X1    g0246(.A(new_n411), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT7), .B1(new_n409), .B2(new_n216), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n402), .B(G68), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n269), .B1(new_n450), .B2(new_n401), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n428), .B1(new_n451), .B2(new_n425), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n442), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n426), .A2(new_n429), .ZN(new_n458));
  INV_X1    g0258(.A(G179), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n433), .A2(new_n434), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(G169), .B2(new_n439), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n457), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(KEYINPUT18), .B(new_n461), .C1(new_n426), .C2(new_n429), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT79), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n426), .B2(new_n429), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n457), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT18), .B1(new_n452), .B2(new_n461), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n456), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n390), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(G244), .B(new_n474), .C1(new_n276), .C2(new_n277), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n476));
  AOI22_X1  g0276(.A1(new_n475), .A2(new_n476), .B1(G33), .B2(G283), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(KEYINPUT4), .A3(G244), .ZN(new_n478));
  INV_X1    g0278(.A(G250), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n474), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n278), .A3(new_n283), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n274), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n291), .A2(G1), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n485), .C1(KEYINPUT5), .C2(new_n290), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n254), .A2(G45), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT84), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G257), .A3(new_n274), .ZN(new_n492));
  INV_X1    g0292(.A(G274), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n272), .B2(new_n273), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n486), .A2(new_n489), .A3(new_n494), .A4(new_n490), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n483), .A2(new_n459), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n492), .ZN(new_n497));
  INV_X1    g0297(.A(new_n495), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n497), .A2(new_n482), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(G169), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n341), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n254), .A2(G33), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n269), .A2(new_n259), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(new_n501), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n284), .A2(new_n418), .B1(KEYINPUT7), .B2(new_n406), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G107), .B1(G77), .B2(new_n262), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n509), .A2(new_n208), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n209), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g0315(.A(new_n216), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n510), .A2(new_n512), .A3(new_n517), .A4(new_n513), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n505), .B1(new_n520), .B2(new_n253), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n500), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  INV_X1    g0323(.A(G200), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n499), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n483), .A2(new_n492), .A3(new_n495), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(KEYINPUT85), .A3(G200), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n499), .A2(G190), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n521), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n281), .A2(new_n282), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n312), .A2(new_n474), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(G244), .C2(new_n474), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n314), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n274), .A2(G274), .A3(new_n484), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT86), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT86), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n494), .A2(new_n538), .A3(new_n484), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n488), .A2(G250), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n314), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT87), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT87), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n545), .B(new_n542), .C1(new_n537), .C2(new_n539), .ZN(new_n546));
  OAI211_X1 g0346(.A(G179), .B(new_n535), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n494), .A2(new_n538), .A3(new_n484), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n538), .B1(new_n494), .B2(new_n484), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n543), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n545), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n540), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n551), .A2(new_n552), .B1(new_n314), .B2(new_n534), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n547), .B1(new_n553), .B2(new_n385), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n504), .A2(new_n374), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n555), .B(KEYINPUT88), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n266), .A2(new_n501), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n530), .A2(new_n216), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n557), .A2(KEYINPUT19), .B1(new_n342), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n321), .A2(KEYINPUT19), .A3(new_n322), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(new_n216), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n253), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n341), .A2(new_n374), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n554), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n535), .B1(new_n544), .B2(new_n546), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  INV_X1    g0368(.A(new_n504), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G87), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n563), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G190), .B(new_n535), .C1(new_n544), .C2(new_n546), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n522), .A2(new_n529), .A3(new_n566), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n259), .A2(G116), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n504), .B2(new_n244), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n280), .A2(G97), .ZN(new_n578));
  INV_X1    g0378(.A(G283), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n216), .B(new_n578), .C1(new_n280), .C2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n252), .A2(new_n217), .B1(G20), .B2(new_n244), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT20), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(KEYINPUT20), .A3(new_n581), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g0386(.A1(G257), .A2(G1698), .ZN(new_n587));
  OAI221_X1 g0387(.A(new_n587), .B1(G264), .B2(new_n474), .C1(new_n276), .C2(new_n277), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G303), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n278), .B2(new_n283), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n314), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n491), .A2(G270), .A3(new_n274), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n495), .A3(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n586), .A2(new_n594), .A3(new_n459), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n575), .B1(new_n569), .B2(G116), .ZN(new_n596));
  INV_X1    g0396(.A(new_n585), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT20), .B1(new_n580), .B2(new_n581), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n594), .A3(G169), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT21), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n599), .A2(new_n594), .A3(new_n602), .A4(G169), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n595), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT22), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n216), .A2(G87), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n284), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n533), .A2(G20), .ZN(new_n609));
  INV_X1    g0409(.A(G107), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(KEYINPUT23), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(KEYINPUT23), .A2(G107), .ZN(new_n613));
  NAND2_X1  g0413(.A1(KEYINPUT22), .A2(G87), .ZN(new_n614));
  OAI221_X1 g0414(.A(new_n612), .B1(new_n216), .B2(new_n613), .C1(new_n558), .C2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT24), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n216), .B2(new_n613), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n558), .A2(new_n614), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT24), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n607), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n253), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n491), .A2(G264), .A3(new_n274), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n479), .A2(new_n474), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(G257), .B2(new_n474), .ZN(new_n626));
  INV_X1    g0426(.A(G294), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n626), .A2(new_n409), .B1(new_n280), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n314), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(G190), .A3(new_n495), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n258), .A2(G20), .A3(new_n610), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT25), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT25), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n633), .B(new_n634), .C1(new_n610), .C2(new_n504), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n624), .A2(new_n495), .A3(new_n629), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G200), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n623), .A2(new_n631), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n599), .B1(new_n594), .B2(G200), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n440), .B2(new_n594), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(G169), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n459), .B2(new_n637), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n269), .B1(new_n616), .B2(new_n621), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n635), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n604), .A2(new_n639), .A3(new_n641), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n574), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n473), .A2(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n467), .A2(new_n468), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n362), .A2(new_n360), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n361), .B1(new_n354), .B2(G169), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n357), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n356), .B2(new_n388), .ZN(new_n653));
  INV_X1    g0453(.A(new_n456), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT90), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n655), .A2(KEYINPUT90), .B1(new_n303), .B2(new_n305), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n309), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n604), .A2(new_n645), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n639), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n574), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n500), .A2(new_n521), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n566), .A2(new_n662), .A3(new_n573), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n566), .A2(new_n662), .A3(new_n573), .A4(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n566), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n661), .B1(new_n668), .B2(KEYINPUT89), .ZN(new_n669));
  INV_X1    g0469(.A(new_n566), .ZN(new_n670));
  AOI211_X1 g0470(.A(KEYINPUT89), .B(new_n670), .C1(new_n665), .C2(new_n666), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n473), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n658), .A2(new_n674), .ZN(G369));
  INV_X1    g0475(.A(new_n604), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n216), .A2(new_n258), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n586), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n604), .A2(new_n641), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT91), .Z(new_n687));
  OR2_X1    g0487(.A1(new_n645), .A2(new_n681), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT93), .ZN(new_n689));
  INV_X1    g0489(.A(new_n681), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n644), .B2(new_n635), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n639), .A2(new_n645), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n604), .A2(new_n690), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n645), .A2(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  NOR2_X1   g0504(.A1(new_n213), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G1), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n560), .A2(new_n244), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n219), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n592), .A2(new_n495), .A3(new_n593), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n499), .A2(new_n713), .A3(new_n630), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n714), .B2(new_n547), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT95), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n594), .A2(new_n459), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n553), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n567), .A2(KEYINPUT95), .A3(new_n459), .A4(new_n594), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(new_n526), .A4(new_n637), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n712), .B(new_n722), .C1(new_n714), .C2(new_n547), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n716), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n690), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n647), .A2(new_n681), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n711), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n690), .B1(new_n669), .B2(new_n672), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n670), .B1(new_n665), .B2(new_n666), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n522), .A2(new_n529), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n566), .A2(new_n573), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n639), .A4(new_n659), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n690), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n729), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n710), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n516), .A2(new_n257), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n707), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n217), .B1(G20), .B2(new_n385), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n216), .A2(new_n459), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n440), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n216), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(G322), .B1(G329), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n524), .A2(G179), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n516), .A2(new_n440), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n579), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n747), .A2(new_n440), .A3(new_n524), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT96), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n755), .B1(new_n762), .B2(G311), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n440), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n216), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n627), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n753), .A2(G20), .A3(G190), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n284), .B1(new_n590), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n747), .A2(new_n440), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n766), .B(new_n768), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n763), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n765), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G97), .ZN(new_n777));
  INV_X1    g0577(.A(G87), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n365), .C1(new_n778), .C2(new_n767), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n247), .A2(new_n774), .B1(new_n769), .B2(new_n342), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n749), .A2(new_n249), .B1(new_n754), .B2(new_n610), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n751), .A2(G159), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT32), .Z(new_n784));
  OAI211_X1 g0584(.A(new_n782), .B(new_n784), .C1(new_n205), .C2(new_n761), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n746), .B1(new_n775), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n745), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n284), .A2(new_n213), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G355), .B1(new_n244), .B2(new_n213), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n250), .A2(G45), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n213), .A2(new_n530), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G45), .B2(new_n219), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n792), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n744), .B(new_n786), .C1(new_n790), .C2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT97), .Z(new_n798));
  INV_X1    g0598(.A(new_n789), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n685), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT98), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n687), .B(new_n744), .C1(G330), .C2(new_n685), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n387), .A2(new_n690), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n384), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n388), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n388), .A2(new_n690), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n730), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT89), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n735), .B1(new_n732), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n681), .B(new_n810), .C1(new_n813), .C2(new_n671), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n729), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n743), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n811), .A2(new_n729), .A3(new_n814), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n745), .A2(new_n787), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT99), .ZN(new_n821));
  INV_X1    g0621(.A(new_n754), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G87), .ZN(new_n823));
  INV_X1    g0623(.A(new_n751), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n627), .B2(new_n749), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n284), .B1(new_n610), .B2(new_n767), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G97), .B2(new_n776), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n579), .B2(new_n769), .C1(new_n590), .C2(new_n774), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n829), .C1(G116), .C2(new_n762), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n770), .A2(G150), .B1(new_n750), .B2(G143), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G159), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n774), .C1(new_n761), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT34), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n754), .A2(new_n342), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n530), .B1(new_n247), .B2(new_n767), .C1(new_n765), .C2(new_n249), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G132), .C2(new_n751), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n830), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n743), .B1(G77), .B2(new_n821), .C1(new_n839), .C2(new_n746), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n787), .B2(new_n809), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  NOR2_X1   g0642(.A1(new_n819), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G384));
  INV_X1    g0644(.A(KEYINPUT106), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n458), .A2(new_n462), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n406), .A2(KEYINPUT7), .ZN(new_n847));
  OAI211_X1 g0647(.A(G68), .B(new_n847), .C1(new_n365), .C2(new_n419), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n848), .B2(new_n423), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n400), .B1(new_n446), .B2(new_n449), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n849), .A2(new_n850), .A3(new_n269), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n680), .B1(new_n851), .B2(new_n428), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n846), .A2(new_n852), .A3(new_n443), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n428), .B(new_n441), .C1(new_n451), .C2(new_n425), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n466), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n852), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n852), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n445), .A2(new_n467), .A3(new_n455), .A4(new_n468), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n859), .A2(KEYINPUT104), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n854), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n450), .A2(new_n396), .A3(new_n399), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n417), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n428), .B1(new_n867), .B2(new_n451), .ZN(new_n868));
  INV_X1    g0668(.A(new_n680), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n443), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n461), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n858), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n868), .A2(new_n869), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT38), .B(new_n873), .C1(new_n471), .C2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n845), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n857), .B1(new_n856), .B2(new_n852), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n857), .A2(new_n846), .A3(new_n852), .A4(new_n443), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT104), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n861), .A2(new_n860), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n864), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT106), .A3(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n725), .A2(new_n726), .ZN(new_n887));
  AND4_X1   g0687(.A1(new_n604), .A2(new_n641), .A3(new_n639), .A4(new_n645), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n888), .A2(new_n733), .A3(new_n734), .A4(new_n681), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n728), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n357), .B(new_n690), .C1(new_n356), .C2(new_n363), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n338), .A2(new_n347), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT75), .B1(new_n354), .B2(G200), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n352), .B(new_n524), .C1(new_n327), .C2(new_n329), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n892), .B(new_n330), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n357), .A2(new_n690), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n652), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  AND4_X1   g0698(.A1(KEYINPUT40), .A2(new_n890), .A3(new_n810), .A4(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n873), .B1(new_n471), .B2(new_n874), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n883), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT103), .A3(new_n875), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT103), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n903), .A3(new_n883), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n890), .A2(new_n810), .A3(new_n898), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n886), .A2(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n473), .A2(new_n890), .ZN(new_n910));
  OAI21_X1  g0710(.A(G330), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n814), .A2(new_n808), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n913), .A2(new_n904), .A3(new_n902), .A4(new_n898), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n649), .A2(new_n869), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n363), .A2(new_n357), .A3(new_n681), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n918));
  XNOR2_X1  g0718(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n884), .A2(new_n875), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n473), .B(new_n737), .C1(new_n730), .C2(KEYINPUT29), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n658), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n912), .A2(new_n925), .B1(new_n254), .B2(new_n740), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n912), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n515), .A2(new_n518), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(G116), .B(new_n218), .C1(new_n929), .C2(KEYINPUT35), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT101), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(KEYINPUT101), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT36), .Z(new_n936));
  NOR3_X1   g0736(.A1(new_n219), .A2(new_n205), .A3(new_n397), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(KEYINPUT102), .ZN(new_n938));
  INV_X1    g0738(.A(new_n201), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(G68), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(KEYINPUT102), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n254), .B(G13), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n927), .A2(new_n936), .A3(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n733), .B1(new_n521), .B2(new_n681), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(new_n645), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n690), .B1(new_n945), .B2(new_n522), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n662), .A2(new_n690), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n695), .A2(new_n699), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n946), .B1(new_n949), .B2(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT42), .B2(new_n949), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n571), .A2(new_n681), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n734), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n566), .B2(new_n952), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n697), .A2(new_n948), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n962));
  XOR2_X1   g0762(.A(new_n705), .B(new_n962), .Z(new_n963));
  NAND3_X1  g0763(.A1(new_n700), .A2(new_n701), .A3(new_n948), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT45), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT44), .B1(new_n703), .B2(new_n948), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  INV_X1    g0768(.A(new_n948), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n702), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n698), .A3(new_n967), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n700), .A2(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n700), .A2(KEYINPUT109), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  INV_X1    g0775(.A(new_n699), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(new_n696), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n695), .A2(KEYINPUT108), .A3(new_n699), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n687), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n974), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n974), .B2(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n967), .A2(new_n970), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n697), .B1(new_n984), .B2(new_n965), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n971), .A2(new_n983), .A3(new_n738), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n963), .B1(new_n986), .B2(new_n738), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n742), .A2(new_n254), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n960), .B(new_n961), .C1(new_n987), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n239), .A2(new_n794), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n745), .B(new_n789), .C1(new_n213), .C2(new_n375), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n744), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n767), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(G116), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n409), .C1(new_n610), .C2(new_n765), .ZN(new_n997));
  INV_X1    g0797(.A(new_n774), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(G311), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n822), .A2(G97), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n590), .B2(new_n749), .C1(new_n824), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n762), .B2(G283), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n999), .B(new_n1003), .C1(new_n627), .C2(new_n769), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n998), .A2(G143), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n770), .A2(G159), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n776), .A2(G68), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n284), .B1(G58), .B2(new_n994), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n822), .A2(G77), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n750), .A2(G150), .B1(G137), .B2(new_n751), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n761), .C2(new_n939), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1004), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n993), .B1(new_n799), .B2(new_n954), .C1(new_n1014), .C2(new_n746), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n983), .A2(new_n738), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n738), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n982), .A3(new_n981), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n705), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n409), .B1(new_n824), .B2(new_n773), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n998), .A2(G322), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n770), .A2(G311), .B1(new_n750), .B2(G317), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n761), .C2(new_n590), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n776), .A2(G283), .B1(G294), .B2(new_n994), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT49), .Z(new_n1030));
  AOI211_X1 g0830(.A(new_n1021), .B(new_n1030), .C1(G116), .C2(new_n822), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n761), .A2(new_n342), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n776), .A2(new_n375), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n409), .B1(new_n994), .B2(G77), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1000), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n824), .A2(new_n261), .B1(new_n247), .B2(new_n749), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n833), .A2(new_n774), .B1(new_n769), .B2(new_n377), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n745), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n794), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n236), .B2(G45), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n708), .B2(new_n791), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n265), .A2(new_n247), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n291), .B1(new_n342), .B2(new_n205), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1044), .A2(new_n708), .A3(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1042), .A2(new_n1046), .B1(G107), .B2(new_n212), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n744), .B1(new_n1047), .B2(new_n790), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1039), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n696), .B2(new_n789), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n983), .B2(new_n989), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1020), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT110), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1020), .A2(KEYINPUT110), .A3(new_n1051), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(G393));
  AND2_X1   g0856(.A1(new_n986), .A2(new_n705), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n971), .A2(new_n985), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n1017), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n971), .A2(new_n989), .A3(new_n985), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n245), .A2(new_n1040), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n790), .B1(new_n501), .B2(new_n212), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n769), .A2(new_n590), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n822), .A2(G107), .B1(G322), .B2(new_n751), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n365), .B1(G283), .B2(new_n994), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n244), .C2(new_n765), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1064), .B(new_n1067), .C1(G294), .C2(new_n762), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n774), .A2(new_n1001), .B1(new_n749), .B2(new_n825), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n769), .A2(new_n939), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n751), .A2(G143), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n776), .A2(G77), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n409), .B1(new_n994), .B2(G68), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n823), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1071), .B(new_n1075), .C1(new_n762), .C2(new_n265), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n774), .A2(new_n261), .B1(new_n749), .B2(new_n833), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1068), .A2(new_n1070), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n743), .B1(new_n1062), .B2(new_n1063), .C1(new_n1079), .C2(new_n746), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT111), .Z(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n799), .B2(new_n948), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1061), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1060), .B1(new_n1085), .B2(new_n1086), .ZN(G390));
  INV_X1    g0887(.A(new_n917), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n681), .B(new_n806), .C1(new_n668), .C2(new_n661), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n808), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n891), .A2(new_n897), .A3(KEYINPUT113), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT113), .B1(new_n891), .B2(new_n897), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1088), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n884), .A2(KEYINPUT106), .A3(new_n875), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT106), .B1(new_n884), .B2(new_n875), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n918), .A2(new_n920), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1088), .B1(new_n913), .B2(new_n898), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n890), .A2(G330), .A3(new_n810), .A4(new_n898), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n989), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n743), .B1(new_n821), .B2(new_n265), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT117), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  INV_X1    g0908(.A(G132), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n824), .A2(new_n1108), .B1(new_n1109), .B2(new_n749), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1111), .A2(new_n774), .B1(new_n769), .B2(new_n832), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n767), .A2(KEYINPUT53), .A3(new_n261), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT53), .B1(new_n767), .B2(new_n261), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n833), .B2(new_n765), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n365), .B1(new_n754), .B2(new_n939), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT118), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1116), .B(new_n1118), .C1(new_n761), .C2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G107), .A2(new_n770), .B1(new_n998), .B2(G283), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n761), .B2(new_n501), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT119), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n836), .B1(G294), .B2(new_n751), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n750), .A2(G116), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n365), .B1(G87), .B2(new_n994), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n1073), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1107), .B1(new_n1128), .B2(new_n745), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1098), .B2(new_n788), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1105), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT120), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n473), .A2(new_n729), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n923), .A2(new_n658), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1093), .B1(new_n729), .B2(new_n810), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n807), .B1(new_n736), .B2(new_n806), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1101), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT114), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n890), .A2(G330), .A3(new_n810), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT114), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n1101), .A4(new_n1137), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n898), .B1(new_n729), .B2(new_n810), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n913), .B1(new_n1145), .B2(new_n1102), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1135), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1103), .A2(new_n1104), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n705), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT115), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1147), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT116), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(KEYINPUT115), .A3(new_n705), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1151), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1133), .A2(new_n1159), .ZN(G378));
  INV_X1    g0960(.A(new_n1135), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1148), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n908), .B(G330), .C1(new_n921), .C2(new_n916), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n906), .A2(new_n907), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n899), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(G330), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n921), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n902), .A2(new_n904), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n898), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n814), .B2(new_n808), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1168), .A2(new_n1170), .B1(new_n649), .B2(new_n869), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1166), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n306), .A2(new_n310), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1173), .B(new_n1174), .Z(new_n1175));
  AND2_X1   g0975(.A1(new_n270), .A2(new_n680), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1163), .A2(new_n1172), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1163), .B2(new_n1172), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1162), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n706), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1162), .B(KEYINPUT57), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT123), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1163), .A2(new_n1172), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1179), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1163), .A2(new_n1172), .A3(new_n1179), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT123), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(KEYINPUT57), .A4(new_n1162), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1184), .A2(new_n1186), .A3(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1177), .A2(new_n788), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n743), .B1(new_n821), .B2(new_n201), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n750), .A2(G107), .B1(G283), .B2(new_n751), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n822), .A2(G58), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G41), .B(new_n530), .C1(new_n994), .C2(G77), .ZN(new_n1199));
  AND4_X1   g0999(.A1(new_n1007), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G97), .A2(new_n770), .B1(new_n998), .B2(G116), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n374), .C2(new_n761), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT58), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n247), .B1(new_n276), .B2(G41), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n765), .A2(new_n261), .B1(new_n767), .B2(new_n1119), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n749), .A2(new_n1111), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G132), .C2(new_n770), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n1108), .B2(new_n774), .C1(new_n832), .C2(new_n761), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n280), .B(new_n290), .C1(new_n754), .C2(new_n833), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G124), .B2(new_n751), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1203), .B(new_n1204), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT121), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n746), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1196), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1191), .A2(new_n989), .B1(new_n1195), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1194), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n989), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n365), .B1(G97), .B2(new_n994), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n1033), .C1(new_n627), .C2(new_n774), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G116), .B2(new_n770), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1010), .B1(new_n824), .B2(new_n590), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G283), .B2(new_n750), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(new_n610), .C2(new_n761), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n409), .B1(new_n994), .B2(G159), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1198), .B(new_n1229), .C1(new_n247), .C2(new_n765), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n824), .A2(new_n1111), .B1(new_n832), .B2(new_n749), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1109), .A2(new_n774), .B1(new_n769), .B2(new_n1119), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n261), .B2(new_n761), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n746), .B1(new_n1235), .B2(KEYINPUT125), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(KEYINPUT125), .B2(new_n1235), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n821), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n744), .B1(new_n1238), .B2(new_n342), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(new_n1093), .C2(new_n788), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1222), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n963), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1153), .A2(new_n1243), .A3(new_n1156), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1144), .A2(new_n1135), .A3(new_n1146), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT124), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT124), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1242), .B1(new_n1244), .B2(new_n1248), .ZN(G381));
  INV_X1    g1049(.A(new_n1086), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1250), .A2(new_n1084), .B1(new_n1059), .B2(new_n1057), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n843), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1054), .A2(new_n801), .A3(new_n802), .A4(new_n1055), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1252), .A2(G387), .A3(G381), .A4(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1133), .A2(new_n1159), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1219), .A4(new_n1194), .ZN(G407));
  INV_X1    g1056(.A(G213), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(G343), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G407), .B(G213), .C1(G375), .C2(new_n1259), .ZN(G409));
  NAND3_X1  g1060(.A1(new_n1194), .A2(G378), .A3(new_n1219), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1219), .B1(new_n963), .B2(new_n1182), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1255), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT126), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1258), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1245), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n706), .B1(new_n1267), .B2(KEYINPUT60), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1152), .A2(KEYINPUT60), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1248), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1242), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n843), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(G384), .A3(new_n1242), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1261), .A2(new_n1263), .A3(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1265), .A2(new_n1266), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1265), .A2(new_n1266), .A3(new_n1277), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1258), .A2(G2897), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1274), .A2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1274), .A2(new_n1282), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1251), .A2(G387), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1253), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G390), .A2(new_n990), .A3(new_n1015), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1288), .A2(new_n1290), .B1(new_n1291), .B2(new_n1287), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  AND4_X1   g1093(.A1(new_n1293), .A2(new_n1290), .A3(new_n1287), .A4(new_n1291), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(KEYINPUT61), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1258), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1275), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1280), .A2(new_n1286), .A3(new_n1296), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1301), .B2(new_n1297), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1278), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1297), .A2(KEYINPUT62), .A3(new_n1275), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1295), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1299), .B1(new_n1306), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1255), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1261), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1275), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1295), .ZN(G402));
endmodule


