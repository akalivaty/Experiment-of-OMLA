//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n188), .B2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n194), .B2(new_n190), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT72), .B(G110), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT16), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G125), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(G146), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n196), .A2(G110), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n191), .A2(new_n192), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(G125), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n203), .B1(new_n213), .B2(new_n201), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(new_n205), .ZN(new_n215));
  AOI21_X1  g029(.A(G146), .B1(new_n200), .B2(new_n203), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n208), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(G137), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n207), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n207), .B2(new_n217), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT74), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(KEYINPUT74), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n225), .A2(new_n226), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n207), .A2(new_n217), .ZN(new_n232));
  INV_X1    g046(.A(new_n222), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n207), .A2(new_n217), .A3(new_n222), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n226), .A3(new_n230), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(G217), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(G234), .B2(new_n226), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n231), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n225), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g057(.A(new_n243), .B(KEYINPUT75), .Z(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  INV_X1    g060(.A(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G134), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n247), .A2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n250), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n246), .B(new_n254), .C1(new_n257), .C2(new_n253), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n205), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n205), .A2(G143), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n187), .B1(KEYINPUT1), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G143), .B(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n251), .A2(G134), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n246), .B1(new_n252), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI211_X1 g087(.A(KEYINPUT66), .B(new_n246), .C1(new_n252), .C2(new_n270), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n258), .B(new_n268), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n265), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT0), .B(G128), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n262), .A2(new_n280), .A3(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n249), .A2(G134), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n285));
  OAI21_X1  g099(.A(G137), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n255), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n253), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n254), .ZN(new_n289));
  OAI21_X1  g103(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n283), .B1(new_n290), .B2(new_n258), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n245), .B1(new_n276), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n258), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT65), .B(G134), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n287), .B1(new_n294), .B2(new_n251), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT11), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n246), .B1(new_n296), .B2(new_n254), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n282), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n265), .B2(G128), .ZN(new_n301));
  AND4_X1   g115(.A1(new_n266), .A2(new_n259), .A3(new_n261), .A4(G128), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n269), .B1(new_n294), .B2(new_n251), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT66), .B1(new_n306), .B2(new_n246), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n271), .A2(new_n272), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n309), .A3(new_n258), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n298), .A2(KEYINPUT30), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT2), .A2(G113), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT67), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT2), .A3(G113), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n317));
  INV_X1    g131(.A(G113), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G116), .B(G119), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n313), .A2(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n321), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT68), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT68), .B1(new_n323), .B2(new_n325), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n292), .A2(new_n311), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n325), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n326), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n298), .A2(new_n334), .A3(new_n310), .ZN(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G210), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n330), .A2(new_n335), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n335), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n298), .A2(new_n334), .A3(new_n310), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n334), .B1(new_n298), .B2(new_n275), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n335), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n341), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(KEYINPUT32), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n345), .A2(new_n346), .B1(new_n341), .B2(new_n354), .ZN(new_n360));
  INV_X1    g174(.A(new_n357), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n348), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n329), .B1(new_n276), .B2(new_n291), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(new_n335), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n335), .A2(new_n352), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n342), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n330), .A2(new_n335), .A3(new_n341), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n334), .B1(new_n298), .B2(new_n310), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT28), .B1(new_n349), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n341), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n353), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n226), .ZN(new_n376));
  OAI21_X1  g190(.A(G472), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT71), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT71), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G472), .C1(new_n370), .C2(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n244), .B1(new_n363), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n387), .A2(new_n390), .A3(new_n394), .A4(new_n391), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(G101), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n387), .A2(new_n390), .A3(new_n338), .A4(new_n391), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n393), .A2(KEYINPUT4), .A3(G101), .A4(new_n395), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n385), .B1(new_n401), .B2(new_n334), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n386), .A2(G107), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n389), .A2(G104), .ZN(new_n404));
  OAI21_X1  g218(.A(G101), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n407));
  INV_X1    g221(.A(G116), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n408), .A2(KEYINPUT5), .A3(G119), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(G113), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n325), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n399), .A2(new_n400), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n329), .A2(KEYINPUT81), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G122), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT82), .Z(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n402), .A2(new_n413), .A3(new_n418), .A4(new_n411), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n421), .A3(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n268), .A2(new_n211), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n282), .A2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n218), .A2(G224), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n425), .B(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n420), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n416), .B(KEYINPUT8), .Z(new_n434));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n406), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n410), .A2(new_n325), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n425), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT86), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n425), .A2(new_n442), .A3(new_n432), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n419), .A2(new_n433), .A3(new_n439), .A4(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n445), .A2(new_n226), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n430), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n430), .A2(new_n448), .A3(new_n446), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n384), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n412), .A2(new_n282), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT78), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n301), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n300), .B(KEYINPUT78), .C1(new_n265), .C2(G128), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n267), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n406), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT10), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n290), .A2(new_n258), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n406), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n453), .A2(new_n460), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G140), .ZN(new_n465));
  INV_X1    g279(.A(G227), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(G953), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n465), .B(new_n467), .Z(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT80), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n453), .A2(new_n460), .A3(new_n463), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(KEYINPUT80), .A3(new_n468), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT79), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n268), .A2(new_n406), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n406), .B2(new_n457), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n478), .B(new_n479), .C1(new_n481), .C2(new_n462), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n458), .B1(new_n268), .B2(new_n406), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(new_n476), .A3(new_n477), .A4(new_n461), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n484), .A3(new_n464), .ZN(new_n485));
  INV_X1    g299(.A(new_n468), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(G469), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  AND4_X1   g303(.A1(new_n464), .A2(new_n482), .A3(new_n484), .A4(new_n468), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n468), .B1(new_n473), .B2(new_n464), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n489), .B(new_n226), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n489), .A2(new_n226), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT9), .B(G234), .Z(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G221), .B1(new_n497), .B2(G902), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT76), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n497), .A2(new_n238), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n408), .A2(KEYINPUT89), .A3(G122), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT89), .B1(new_n408), .B2(G122), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n408), .A2(G122), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(G116), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n408), .A2(KEYINPUT89), .A3(G122), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT92), .B1(new_n519), .B2(new_n511), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n514), .A3(new_n518), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n522), .A2(new_n523), .A3(G107), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n522), .B2(G107), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n518), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n389), .A3(new_n512), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT90), .B1(new_n187), .B2(G143), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n260), .A3(G128), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n260), .A2(G128), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n532), .A2(new_n294), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n256), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n527), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n524), .A2(new_n525), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n527), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n389), .B1(new_n526), .B2(new_n512), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT91), .B(new_n535), .C1(new_n532), .C2(KEYINPUT13), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(KEYINPUT13), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT13), .B1(new_n528), .B2(new_n530), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n533), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n534), .B(new_n541), .C1(new_n547), .C2(G134), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n506), .B1(new_n538), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n541), .B1(new_n547), .B2(G134), .ZN(new_n550));
  INV_X1    g364(.A(new_n534), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n522), .A2(G107), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n522), .A2(new_n523), .A3(G107), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n552), .B(new_n505), .C1(new_n556), .C2(new_n537), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n504), .B1(new_n558), .B2(new_n226), .ZN(new_n559));
  AOI211_X1 g373(.A(G902), .B(new_n503), .C1(new_n549), .C2(new_n557), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G952), .ZN(new_n563));
  AOI211_X1 g377(.A(G953), .B(new_n563), .C1(G234), .C2(G237), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT21), .B(G898), .Z(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n226), .B(new_n218), .C1(G234), .C2(G237), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT18), .A2(G131), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n572));
  AOI21_X1  g386(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n569), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n213), .A2(G146), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n206), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n572), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n577), .B2(KEYINPUT87), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(KEYINPUT87), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n574), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G131), .B1(new_n572), .B2(new_n573), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n582));
  INV_X1    g396(.A(G237), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(new_n218), .A3(G214), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n260), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n246), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n581), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n214), .A2(new_n205), .ZN(new_n589));
  OAI211_X1 g403(.A(KEYINPUT17), .B(G131), .C1(new_n572), .C2(new_n573), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n204), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G113), .B(G122), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT88), .B(G104), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n580), .A2(new_n597), .A3(new_n591), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n226), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G475), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n581), .A2(new_n587), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n213), .A2(KEYINPUT19), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n213), .A2(KEYINPUT19), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n603), .B(new_n204), .C1(new_n606), .C2(G146), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n580), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n595), .ZN(new_n609));
  AOI21_X1  g423(.A(G475), .B1(new_n609), .B2(new_n598), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n602), .B1(new_n610), .B2(new_n226), .ZN(new_n611));
  INV_X1    g425(.A(G475), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n580), .A2(new_n597), .A3(new_n591), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n597), .B1(new_n580), .B2(new_n607), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n612), .B(new_n226), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(KEYINPUT20), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n601), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n562), .A2(new_n568), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n382), .A2(new_n452), .A3(new_n501), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  INV_X1    g434(.A(new_n568), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n430), .A2(new_n448), .A3(new_n446), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n448), .B1(new_n430), .B2(new_n446), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n383), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n549), .A2(KEYINPUT33), .A3(new_n557), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT33), .B1(new_n549), .B2(new_n557), .ZN(new_n626));
  OAI21_X1  g440(.A(G478), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n558), .A2(new_n502), .A3(new_n226), .ZN(new_n628));
  NAND2_X1  g442(.A1(G478), .A2(G902), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n627), .A2(new_n617), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT94), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n630), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n452), .A2(new_n632), .A3(new_n633), .A4(new_n621), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n361), .B1(new_n347), .B2(new_n355), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n360), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n244), .A2(new_n639), .A3(new_n500), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  OAI21_X1  g457(.A(KEYINPUT95), .B1(new_n611), .B2(new_n616), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n610), .A2(new_n602), .A3(new_n226), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n615), .A2(KEYINPUT20), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n644), .A2(new_n648), .B1(G475), .B2(new_n600), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n562), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n640), .A2(new_n452), .A3(new_n621), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n232), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n241), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n240), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n240), .A2(KEYINPUT96), .A3(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n383), .B(new_n661), .C1(new_n622), .C2(new_n623), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n639), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n501), .A3(new_n618), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G12));
  AOI21_X1  g482(.A(new_n341), .B1(new_n351), .B2(new_n353), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n330), .A2(new_n335), .A3(new_n341), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n373), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n375), .A2(new_n226), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n379), .B1(new_n673), .B2(G472), .ZN(new_n674));
  INV_X1    g488(.A(new_n380), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n362), .B(new_n358), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n564), .B1(new_n567), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n562), .A2(new_n649), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n676), .A2(new_n663), .A3(new_n501), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XOR2_X1   g496(.A(KEYINPUT99), .B(KEYINPUT39), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n678), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n501), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT100), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n450), .A2(new_n451), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT38), .Z(new_n689));
  INV_X1    g503(.A(new_n371), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n335), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(KEYINPUT98), .A3(new_n341), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n343), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT98), .B1(new_n691), .B2(new_n341), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n226), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G472), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n358), .A2(new_n362), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n689), .A2(new_n657), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n617), .A2(new_n383), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n561), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n687), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NOR2_X1   g517(.A1(new_n630), .A2(new_n678), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n676), .A2(new_n663), .A3(new_n501), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(new_n244), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n490), .A2(new_n491), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n226), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n498), .A3(new_n492), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n676), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n713), .A2(new_n635), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n714), .B1(new_n713), .B2(new_n635), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT41), .B(G113), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  OAI21_X1  g533(.A(new_n383), .B1(new_n622), .B2(new_n623), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n711), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n382), .A2(new_n621), .A3(new_n650), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n676), .A3(new_n618), .A4(new_n661), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  OAI21_X1  g539(.A(new_n701), .B1(new_n622), .B2(new_n623), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT102), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT102), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n701), .B(new_n728), .C1(new_n622), .C2(new_n623), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n367), .B1(new_n691), .B2(KEYINPUT28), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n347), .B1(new_n342), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n357), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n243), .A3(new_n638), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n621), .A3(new_n712), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AND3_X1   g550(.A1(new_n733), .A2(new_n638), .A3(new_n657), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n721), .A2(new_n704), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n495), .A2(new_n498), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n688), .A2(new_n384), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n704), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT104), .B1(new_n636), .B2(KEYINPUT32), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n360), .A2(new_n744), .A3(new_n359), .A4(new_n361), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n362), .A2(KEYINPUT105), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n636), .A2(KEYINPUT105), .A3(KEYINPUT32), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n381), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT106), .B1(new_n749), .B2(new_n243), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n381), .B1(new_n743), .B2(new_n745), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n747), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT106), .B(new_n243), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT42), .B(new_n742), .C1(new_n750), .C2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n741), .A2(new_n676), .A3(new_n707), .A4(new_n704), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT103), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT103), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND3_X1  g578(.A1(new_n382), .A2(new_n680), .A3(new_n741), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  AND2_X1   g580(.A1(new_n627), .A2(new_n629), .ZN(new_n767));
  INV_X1    g581(.A(new_n617), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n628), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT43), .ZN(new_n770));
  INV_X1    g584(.A(new_n657), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n770), .A2(new_n664), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT108), .Z(new_n775));
  NOR2_X1   g589(.A1(new_n688), .A2(new_n384), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n778));
  INV_X1    g592(.A(new_n487), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n475), .A2(KEYINPUT45), .A3(new_n487), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n494), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n492), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT46), .B1(new_n784), .B2(new_n494), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n498), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n684), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n773), .B2(new_n772), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(new_n776), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NAND2_X1  g607(.A1(new_n789), .A2(KEYINPUT47), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n676), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n244), .A3(new_n704), .A4(new_n776), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NAND2_X1  g613(.A1(new_n776), .A2(new_n712), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n776), .A2(new_n712), .A3(KEYINPUT115), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n244), .A2(new_n697), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n564), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n617), .B1(new_n767), .B2(new_n628), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT117), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n802), .A2(new_n564), .A3(new_n803), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n770), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n737), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n710), .A2(new_n492), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n794), .B(new_n796), .C1(new_n499), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n734), .A2(new_n564), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n770), .A2(new_n822), .A3(new_n384), .A4(new_n688), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n689), .A2(new_n384), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n770), .A2(new_n711), .A3(new_n822), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT50), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT114), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT114), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n821), .A2(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n563), .B(G953), .C1(new_n809), .C2(new_n632), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT51), .B1(new_n827), .B2(new_n828), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n821), .B2(new_n823), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n819), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n813), .B1(new_n750), .B2(new_n754), .ZN(new_n840));
  NAND2_X1  g654(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n834), .A2(new_n839), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n826), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n720), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT119), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n681), .A2(new_n738), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  INV_X1    g665(.A(new_n740), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n697), .A2(new_n771), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n730), .A2(new_n853), .A3(new_n679), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n850), .A2(new_n851), .A3(new_n705), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n681), .A2(new_n705), .A3(new_n738), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n730), .A2(new_n853), .A3(new_n679), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT52), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n855), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n649), .A2(new_n863), .A3(new_n561), .A4(new_n679), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(new_n661), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n649), .A2(new_n561), .A3(new_n679), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n676), .A2(new_n865), .A3(new_n501), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n737), .A2(new_n704), .A3(new_n852), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n776), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n765), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n735), .A2(new_n722), .A3(new_n724), .ZN(new_n874));
  INV_X1    g688(.A(new_n716), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n713), .A2(new_n635), .A3(new_n714), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT110), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n624), .B2(new_n630), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n452), .A2(new_n632), .A3(KEYINPUT110), .A4(new_n621), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n561), .A2(new_n617), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n624), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n640), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n619), .A3(new_n665), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n763), .A2(new_n873), .A3(new_n877), .A4(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n849), .B1(new_n862), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n717), .A2(new_n886), .A3(new_n874), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n872), .B1(new_n755), .B2(new_n762), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n855), .A2(new_n858), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n892), .A3(new_n894), .A4(KEYINPUT53), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n849), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT112), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n763), .A2(new_n873), .A3(new_n877), .A4(new_n887), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(KEYINPUT113), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT112), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n905), .A3(new_n849), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n896), .B1(new_n907), .B2(KEYINPUT54), .ZN(new_n908));
  INV_X1    g722(.A(new_n838), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n835), .B(new_n844), .C1(new_n909), .C2(new_n818), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT51), .B1(new_n819), .B2(new_n831), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n913));
  INV_X1    g727(.A(new_n847), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(new_n842), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n848), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n563), .A2(new_n218), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT109), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n243), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n769), .B(new_n921), .C1(KEYINPUT49), .C2(new_n820), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n499), .A2(new_n383), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n698), .A3(new_n689), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n918), .A2(new_n924), .ZN(G75));
  AOI21_X1  g739(.A(new_n226), .B1(new_n889), .B2(new_n895), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G210), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT55), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n420), .A2(new_n422), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n429), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n218), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(G51));
  NAND3_X1  g754(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n889), .A2(new_n895), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n889), .A2(KEYINPUT121), .A3(new_n890), .A4(new_n895), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n494), .A2(KEYINPUT57), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n494), .A2(KEYINPUT57), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n708), .ZN(new_n951));
  INV_X1    g765(.A(new_n784), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n926), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n938), .B1(new_n951), .B2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(KEYINPUT122), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n926), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT122), .B1(KEYINPUT58), .B2(G475), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n609), .A2(new_n598), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n938), .ZN(G60));
  OR2_X1    g775(.A1(new_n625), .A2(new_n626), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n629), .B(KEYINPUT59), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n947), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n962), .B1(new_n908), .B2(new_n963), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n947), .A2(KEYINPUT123), .A3(new_n964), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n967), .A2(new_n939), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(new_n963), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n897), .A2(new_n905), .A3(new_n849), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n905), .B1(new_n897), .B2(new_n849), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n890), .B1(new_n975), .B2(new_n904), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n972), .B1(new_n976), .B2(new_n896), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n938), .B1(new_n977), .B2(new_n962), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n978), .A2(new_n979), .A3(new_n967), .A4(new_n969), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n971), .A2(new_n980), .ZN(G63));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT60), .Z(new_n983));
  AND2_X1   g797(.A1(new_n944), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n938), .B1(new_n984), .B2(new_n655), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n225), .B2(new_n984), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT61), .Z(G66));
  INV_X1    g801(.A(new_n891), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n218), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n218), .B1(new_n565), .B2(G224), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n933), .B1(G898), .B2(new_n218), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n992), .B(new_n993), .Z(G69));
  INV_X1    g808(.A(new_n856), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n702), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT62), .Z(new_n997));
  NAND2_X1  g811(.A1(new_n883), .A2(new_n630), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n686), .A2(new_n382), .A3(new_n776), .A4(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n997), .A2(new_n792), .A3(new_n798), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n292), .A2(new_n311), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT126), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(new_n606), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1000), .A2(new_n218), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n218), .A2(G900), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n730), .B1(new_n750), .B2(new_n754), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n763), .B(new_n765), .C1(new_n790), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n792), .A2(new_n798), .A3(new_n995), .A4(new_n1008), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n1005), .B(new_n1003), .C1(new_n1009), .C2(new_n218), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(G953), .B1(new_n466), .B2(new_n677), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n1000), .B2(new_n988), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n341), .B1(new_n330), .B2(new_n335), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1019), .B(new_n1015), .C1(new_n1000), .C2(new_n988), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1009), .B2(new_n988), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n938), .B1(new_n1022), .B2(new_n670), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n907), .A2(new_n369), .A3(new_n1015), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n1024), .A2(new_n1018), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .ZN(G57));
endmodule


