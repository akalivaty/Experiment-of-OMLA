//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n209), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n212), .A2(new_n213), .B1(new_n202), .B2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n216), .A2(new_n217), .B1(new_n205), .B2(new_n218), .ZN(new_n219));
  NOR3_X1   g0019(.A1(new_n211), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT67), .B(G238), .Z(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(new_n201), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n220), .A2(new_n222), .B1(G1), .B2(G20), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n212), .A2(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  OAI22_X1  g0035(.A1(new_n223), .A2(new_n224), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(G1), .ZN(new_n237));
  NOR3_X1   g0037(.A1(new_n237), .A2(new_n225), .A3(G13), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n238), .B(G250), .C1(G257), .C2(G264), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(KEYINPUT64), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT0), .ZN(new_n241));
  AOI211_X1 g0041(.A(new_n236), .B(new_n241), .C1(new_n224), .C2(new_n223), .ZN(G361));
  XOR2_X1   g0042(.A(G238), .B(G244), .Z(new_n243));
  XNOR2_X1  g0043(.A(G226), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G250), .B(G257), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G264), .B(G270), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G358));
  NAND2_X1  g0052(.A1(G68), .A2(G77), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n203), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n254), .B(KEYINPUT70), .Z(new_n255));
  XNOR2_X1  g0055(.A(G50), .B(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(G87), .B(G97), .Z(new_n258));
  XNOR2_X1  g0058(.A(G107), .B(G116), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n257), .B(new_n260), .Z(G351));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n266), .A2(G223), .B1(G77), .B2(new_n264), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n231), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n237), .B1(G41), .B2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n237), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n231), .B2(new_n271), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n272), .A2(new_n275), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n274), .B(new_n286), .C1(new_n217), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G179), .B2(new_n288), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n237), .A2(G13), .A3(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n230), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n237), .B2(G20), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(new_n296), .B2(G50), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G50), .A2(G58), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n225), .B1(new_n299), .B2(new_n201), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n302), .A2(new_n212), .A3(KEYINPUT8), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT65), .B(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(G150), .ZN(new_n308));
  INV_X1    g0108(.A(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n225), .A2(new_n309), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n305), .A2(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI221_X1 g0113(.A(KEYINPUT74), .B1(new_n308), .B2(new_n310), .C1(new_n305), .C2(new_n307), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n298), .B1(new_n315), .B2(new_n295), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n291), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n288), .A2(G200), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n288), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n311), .A2(new_n312), .ZN(new_n322));
  INV_X1    g0122(.A(new_n300), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n322), .A2(new_n314), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n294), .A2(new_n230), .ZN(new_n325));
  OAI211_X1 g0125(.A(KEYINPUT9), .B(new_n297), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT80), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT80), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n316), .A2(new_n328), .A3(KEYINPUT9), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n321), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT10), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n297), .B1(new_n324), .B2(new_n325), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(KEYINPUT79), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT79), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n316), .B2(KEYINPUT9), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n330), .A2(new_n331), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n331), .B1(new_n330), .B2(new_n337), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n318), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G20), .A2(G33), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n307), .B2(new_n202), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n344), .A2(new_n295), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(KEYINPUT11), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(KEYINPUT11), .ZN(new_n347));
  OR3_X1    g0147(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT12), .B1(new_n292), .B2(G68), .ZN(new_n349));
  AOI22_X1  g0149(.A1(G68), .A2(new_n296), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n272), .A2(G238), .A3(new_n275), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n286), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n268), .A2(G226), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n266), .A2(G232), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT81), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT81), .A4(new_n359), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n273), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n356), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n356), .B2(new_n364), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n353), .B(G169), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n356), .A2(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(G179), .A3(new_n366), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n366), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n353), .B1(new_n374), .B2(G169), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n352), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(G200), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(G190), .A3(new_n366), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n351), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT82), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n286), .B1(new_n214), .B2(new_n287), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n268), .A2(G232), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT3), .B(G33), .ZN(new_n386));
  INV_X1    g0186(.A(new_n266), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n385), .B1(new_n206), .B2(new_n386), .C1(new_n221), .C2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n383), .A2(new_n384), .B1(new_n273), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n286), .B(KEYINPUT75), .C1(new_n214), .C2(new_n287), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n289), .ZN(new_n392));
  INV_X1    g0192(.A(G179), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT15), .B(G87), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT77), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n399), .A2(new_n307), .B1(new_n202), .B2(new_n306), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n301), .B(KEYINPUT76), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n342), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n325), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n296), .A2(G77), .ZN(new_n404));
  XOR2_X1   g0204(.A(new_n404), .B(KEYINPUT78), .Z(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G77), .B2(new_n292), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n392), .B(new_n394), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n389), .B2(new_n390), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n403), .A2(new_n406), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n389), .A2(G190), .A3(new_n390), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n262), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT83), .B(G33), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n306), .C1(new_n417), .C2(KEYINPUT3), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n386), .B2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n201), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT84), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n225), .B1(new_n234), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G159), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n310), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n422), .ZN(new_n427));
  NOR2_X1   g0227(.A1(G58), .A2(G68), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n342), .A2(G159), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT84), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n414), .B1(new_n420), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT85), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n432), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT83), .A2(G33), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT83), .A2(G33), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT3), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n263), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT7), .B1(new_n441), .B2(G20), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n306), .A2(new_n415), .ZN(new_n444));
  OAI21_X1  g0244(.A(G68), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n436), .B(KEYINPUT16), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(KEYINPUT85), .B(new_n414), .C1(new_n420), .C2(new_n432), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n435), .A2(new_n295), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n305), .A2(new_n292), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n305), .B2(new_n296), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n263), .B1(new_n417), .B2(KEYINPUT3), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n217), .A2(G1698), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(G223), .B2(G1698), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G87), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n309), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n273), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT86), .B1(new_n287), .B2(new_n213), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT86), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n272), .A2(new_n460), .A3(G232), .A4(new_n275), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n286), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G169), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n393), .B2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n451), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT18), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT18), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n451), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(new_n408), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n286), .A2(new_n458), .A3(new_n320), .A4(new_n462), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n448), .A3(new_n450), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT17), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n472), .A2(new_n448), .A3(KEYINPUT17), .A4(new_n450), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n467), .A2(new_n469), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n413), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n376), .A2(KEYINPUT82), .A3(new_n379), .ZN(new_n479));
  AND4_X1   g0279(.A1(new_n341), .A2(new_n382), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G303), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n386), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n218), .B1(new_n439), .B2(new_n440), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n265), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT90), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G264), .A2(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n441), .B2(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(KEYINPUT90), .B(new_n487), .C1(new_n439), .C2(new_n440), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n485), .B(KEYINPUT91), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT90), .B1(new_n452), .B2(new_n487), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n441), .A2(new_n486), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT91), .B1(new_n495), .B2(new_n485), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n273), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT92), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT91), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n489), .A2(new_n490), .ZN(new_n500));
  INV_X1    g0300(.A(new_n483), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n441), .A2(G257), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G1698), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n491), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT92), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n273), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(new_n272), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G270), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n281), .B(new_n510), .C1(new_n512), .C2(new_n511), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n508), .A2(G190), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n205), .B2(G33), .ZN(new_n521));
  OAI221_X1 g0321(.A(new_n295), .B1(new_n225), .B2(G116), .C1(new_n229), .C2(new_n521), .ZN(new_n522));
  XOR2_X1   g0322(.A(new_n522), .B(KEYINPUT20), .Z(new_n523));
  NOR2_X1   g0323(.A1(new_n292), .A2(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n325), .B(new_n292), .C1(G1), .C2(new_n309), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n526), .B2(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n517), .B1(new_n498), .B2(new_n507), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n519), .B(new_n529), .C1(new_n408), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(G169), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n506), .B1(new_n505), .B2(new_n273), .ZN(new_n535));
  AOI211_X1 g0335(.A(KEYINPUT92), .B(new_n272), .C1(new_n504), .C2(new_n491), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n518), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n533), .A2(new_n532), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n517), .A2(new_n393), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(new_n538), .B1(new_n508), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n531), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n292), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT25), .B1(new_n543), .B2(new_n206), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n545), .A2(new_n546), .B1(new_n525), .B2(new_n206), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n229), .A2(new_n548), .A3(new_n206), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n417), .A2(new_n225), .A3(G116), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT23), .B1(new_n225), .B2(G107), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n441), .A2(KEYINPUT22), .A3(G87), .A4(new_n306), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n386), .A2(new_n306), .A3(G87), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT24), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n547), .B1(new_n558), .B2(new_n295), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n441), .A2(G250), .A3(new_n265), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n417), .A2(G294), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n502), .C2(new_n265), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n273), .B1(G264), .B2(new_n514), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n516), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(G190), .A3(new_n516), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT93), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n564), .B2(new_n393), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n289), .B1(new_n563), .B2(new_n516), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n563), .A2(KEYINPUT93), .A3(G179), .A4(new_n516), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n325), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n575), .B2(new_n547), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n567), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g0377(.A(KEYINPUT87), .B(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n207), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n205), .A2(G107), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n582), .A2(new_n306), .B1(new_n202), .B2(new_n310), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n206), .B1(new_n418), .B2(new_n419), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n295), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n292), .A2(G97), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n526), .B2(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n214), .B1(new_n439), .B2(new_n440), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT4), .B1(new_n589), .B2(new_n265), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n386), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n386), .A2(G250), .A3(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n520), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n273), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n513), .A2(new_n272), .A3(G257), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n516), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT88), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT88), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n516), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n588), .B1(new_n600), .B2(G200), .ZN(new_n601));
  INV_X1    g0401(.A(new_n600), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G190), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(G1698), .B1(new_n439), .B2(new_n440), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(G238), .B1(G116), .B2(new_n417), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n441), .A2(G244), .A3(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n272), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n272), .B(G250), .C1(G1), .C2(new_n509), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n281), .A2(new_n510), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n289), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n441), .A2(G238), .A3(new_n265), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n417), .A2(G116), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n607), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n273), .ZN(new_n616));
  INV_X1    g0416(.A(new_n611), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n393), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n441), .A2(G68), .A3(new_n306), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n306), .B1(new_n620), .B2(new_n359), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n456), .A2(new_n205), .A3(new_n206), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n306), .A2(G33), .A3(G97), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n620), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n295), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n292), .B1(new_n397), .B2(new_n398), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n399), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n526), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n612), .A2(new_n618), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n608), .B2(new_n611), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n616), .A2(G190), .A3(new_n617), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n525), .A2(new_n456), .ZN(new_n636));
  AOI211_X1 g0436(.A(new_n636), .B(new_n628), .C1(new_n626), .C2(new_n295), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n600), .A2(new_n289), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n594), .A2(new_n393), .A3(new_n597), .A4(new_n599), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n588), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n604), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n481), .A2(new_n542), .A3(new_n577), .A4(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n467), .A2(new_n469), .ZN(new_n645));
  INV_X1    g0445(.A(new_n379), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n376), .B1(new_n646), .B2(new_n407), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n475), .A2(new_n476), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n338), .A2(new_n339), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n317), .ZN(new_n653));
  INV_X1    g0453(.A(new_n642), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT26), .B1(new_n639), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n633), .A2(new_n638), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n642), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n633), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n576), .ZN(new_n660));
  INV_X1    g0460(.A(new_n570), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n661), .B(new_n568), .C1(new_n393), .C2(new_n564), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n541), .A2(new_n534), .A3(new_n663), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n567), .A2(new_n642), .A3(new_n604), .A4(new_n639), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n653), .B1(new_n481), .B2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n306), .A2(new_n237), .A3(G13), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT94), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n672));
  INV_X1    g0472(.A(G213), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n529), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n542), .B2(KEYINPUT95), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n540), .B1(new_n535), .B2(new_n536), .ZN(new_n680));
  INV_X1    g0480(.A(new_n538), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n530), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n533), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT21), .B1(new_n537), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT95), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n531), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n678), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n559), .A2(new_n677), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n577), .A2(new_n690), .B1(new_n663), .B2(new_n677), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n688), .A2(G330), .A3(new_n689), .A4(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n577), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n693), .B(new_n677), .C1(new_n684), .C2(new_n682), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n660), .A2(new_n662), .A3(new_n677), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT96), .Z(G399));
  INV_X1    g0499(.A(new_n238), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n622), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n704), .A2(KEYINPUT97), .B1(new_n235), .B2(new_n702), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(KEYINPUT97), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  NOR2_X1   g0507(.A1(new_n577), .A2(new_n643), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n685), .A2(new_n708), .A3(new_n531), .A4(new_n677), .ZN(new_n709));
  INV_X1    g0509(.A(new_n677), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n600), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n608), .A2(new_n611), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n539), .A3(new_n563), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n712), .B(new_n715), .C1(new_n535), .C2(new_n536), .ZN(new_n716));
  INV_X1    g0516(.A(new_n713), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n564), .A3(new_n393), .A4(new_n600), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n530), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n498), .B2(new_n507), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT30), .B1(new_n720), .B2(new_n602), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n710), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT31), .B(new_n710), .C1(new_n719), .C2(new_n721), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n709), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  OR3_X1    g0527(.A1(new_n666), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT29), .B1(new_n666), .B2(new_n710), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n707), .B1(new_n731), .B2(G1), .ZN(G364));
  NAND3_X1  g0532(.A1(new_n688), .A2(G330), .A3(new_n689), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n306), .A2(G13), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G1), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n701), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n689), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n679), .B2(new_n687), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n386), .A2(new_n238), .ZN(new_n749));
  INV_X1    g0549(.A(G355), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n749), .A2(new_n750), .B1(G116), .B2(new_n238), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n257), .A2(G45), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n441), .A2(new_n700), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n235), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(new_n509), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n751), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n230), .B1(G20), .B2(new_n289), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n737), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n408), .A2(G179), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G20), .A3(G190), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n264), .B1(new_n763), .B2(new_n482), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n306), .A2(G190), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G179), .A3(G200), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n306), .B1(G190), .B2(new_n769), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n306), .A2(new_n393), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n764), .B(new_n771), .C1(G311), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n408), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G322), .A2(new_n778), .B1(new_n779), .B2(G326), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n765), .A2(new_n769), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G329), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n765), .A2(new_n762), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT99), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G283), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n776), .A2(new_n780), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(G159), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(G107), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n386), .B1(new_n763), .B2(new_n456), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n775), .B2(G77), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G50), .A2(new_n779), .B1(new_n778), .B2(G58), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n770), .A2(new_n205), .ZN(new_n797));
  INV_X1    g0597(.A(new_n766), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(G68), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n793), .A2(new_n795), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n790), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n761), .B1(new_n801), .B2(new_n758), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n744), .B1(new_n748), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  NOR2_X1   g0604(.A1(new_n666), .A2(new_n710), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n407), .A2(new_n710), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n412), .A2(new_n409), .B1(new_n410), .B2(new_n677), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n407), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n805), .B(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n737), .B1(new_n809), .B2(new_n727), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n727), .B2(new_n809), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n758), .A2(new_n745), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n738), .B1(new_n202), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n758), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n441), .B1(new_n784), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT103), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n788), .A2(G68), .ZN(new_n818));
  INV_X1    g0618(.A(new_n770), .ZN(new_n819));
  INV_X1    g0619(.A(new_n763), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n819), .A2(G58), .B1(new_n820), .B2(G50), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n816), .A2(KEYINPUT103), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n798), .A2(G150), .B1(new_n775), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(new_n778), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  INV_X1    g0628(.A(new_n779), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n825), .B1(new_n826), .B2(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n779), .A2(G303), .B1(new_n775), .B2(G116), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n766), .A2(KEYINPUT100), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n766), .A2(KEYINPUT100), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT101), .B(G283), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT102), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n788), .A2(G87), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n785), .A2(G311), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n386), .B(new_n797), .C1(G107), .C2(new_n820), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n778), .A2(G294), .ZN(new_n842));
  AND4_X1   g0642(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n824), .A2(new_n831), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n813), .B1(new_n814), .B2(new_n844), .C1(new_n808), .C2(new_n746), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n811), .A2(new_n845), .ZN(G384));
  XOR2_X1   g0646(.A(new_n582), .B(KEYINPUT35), .Z(new_n847));
  INV_X1    g0647(.A(G116), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n847), .A2(new_n848), .A3(new_n233), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n755), .A2(G77), .A3(new_n422), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n216), .A2(G68), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n237), .B(G13), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n373), .A2(new_n375), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n352), .B(new_n710), .C1(new_n856), .C2(new_n646), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n376), .B(new_n379), .C1(new_n351), .C2(new_n677), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n806), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n654), .B1(new_n603), .B2(new_n601), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n567), .A3(new_n639), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n685), .B2(new_n663), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n677), .B(new_n808), .C1(new_n863), .C2(new_n659), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n859), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n446), .A2(new_n295), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n442), .B(G68), .C1(new_n441), .C2(new_n444), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n867), .B2(new_n436), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n450), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n465), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n676), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n473), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n451), .A2(new_n676), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n466), .A2(new_n874), .A3(new_n875), .A4(new_n473), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n477), .A2(new_n676), .A3(new_n869), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n873), .A2(new_n876), .A3(KEYINPUT105), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT38), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n865), .A2(new_n886), .B1(new_n645), .B2(new_n675), .ZN(new_n887));
  INV_X1    g0687(.A(new_n874), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n477), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n466), .A2(new_n874), .A3(new_n473), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n876), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT106), .B1(new_n477), .B2(new_n888), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n883), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n885), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n856), .A2(new_n352), .A3(new_n677), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n887), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n728), .A2(new_n729), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n480), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n653), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n903), .B(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n895), .A2(new_n885), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n857), .A2(new_n858), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n726), .A2(new_n909), .A3(new_n808), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT40), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n726), .A2(new_n909), .A3(new_n808), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT40), .B1(new_n884), .B2(new_n885), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n480), .A2(new_n726), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n740), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n907), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n237), .B2(new_n734), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n907), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n855), .B1(new_n920), .B2(new_n921), .ZN(G367));
  OAI22_X1  g0722(.A1(new_n835), .A2(new_n424), .B1(new_n784), .B2(new_n828), .ZN(new_n923));
  INV_X1    g0723(.A(new_n787), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(G77), .B1(new_n819), .B2(G68), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n264), .B1(new_n820), .B2(G58), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n926), .C1(new_n216), .C2(new_n774), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n827), .A2(new_n829), .B1(new_n826), .B2(new_n308), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT114), .Z(new_n930));
  XOR2_X1   g0730(.A(KEYINPUT112), .B(G317), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n785), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n452), .C1(new_n205), .C2(new_n787), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(KEYINPUT113), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT111), .B(G311), .Z(new_n935));
  OAI22_X1  g0735(.A1(new_n482), .A2(new_n826), .B1(new_n829), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n820), .A2(G116), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT46), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n206), .B2(new_n770), .C1(new_n774), .C2(new_n836), .ZN(new_n939));
  INV_X1    g0739(.A(new_n835), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n936), .B(new_n939), .C1(G294), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n933), .A2(KEYINPUT113), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n930), .B1(new_n934), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n758), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n639), .B1(new_n637), .B2(new_n677), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n633), .A2(new_n677), .A3(new_n637), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n747), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n251), .A2(new_n753), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n760), .B1(new_n630), .B2(new_n700), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n738), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n946), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT110), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n685), .A2(new_n710), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n694), .B1(new_n957), .B2(new_n691), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n742), .A2(G330), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n742), .B2(G330), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n956), .B1(new_n961), .B2(new_n730), .ZN(new_n962));
  INV_X1    g0762(.A(new_n958), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n733), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n742), .A2(G330), .A3(new_n958), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(KEYINPUT110), .A3(new_n731), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n710), .A2(new_n588), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n861), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n654), .A2(new_n710), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n694), .A2(new_n695), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  INV_X1    g0775(.A(new_n971), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT44), .B1(new_n696), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n978), .B(new_n971), .C1(new_n694), .C2(new_n695), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n974), .A2(new_n975), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n692), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n962), .A2(new_n967), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n731), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n701), .B(new_n984), .Z(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n736), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n957), .A2(new_n693), .A3(new_n971), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n642), .B1(new_n969), .B2(new_n663), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n989), .A2(KEYINPUT42), .B1(new_n677), .B2(new_n990), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n976), .A2(new_n694), .A3(KEYINPUT42), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n950), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n991), .A2(new_n994), .A3(new_n950), .A4(new_n992), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n692), .A2(new_n976), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n988), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n1000), .A3(KEYINPUT108), .A4(new_n998), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT107), .B1(new_n999), .B2(new_n1001), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1005), .A3(new_n1003), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n955), .B1(new_n987), .B2(new_n1009), .ZN(G387));
  OR3_X1    g0810(.A1(new_n691), .A2(G20), .A3(new_n746), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n749), .A2(new_n703), .B1(G107), .B2(new_n238), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n401), .A2(new_n216), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT50), .Z(new_n1014));
  NAND4_X1  g0814(.A1(new_n1014), .A2(new_n509), .A3(new_n253), .A4(new_n703), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n754), .B1(new_n247), .B2(G45), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n737), .B1(new_n1017), .B2(new_n760), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n788), .A2(G97), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n452), .B1(G77), .B2(new_n820), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n308), .C2(new_n784), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT115), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n305), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n798), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n399), .A2(new_n770), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G68), .B2(new_n775), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G50), .A2(new_n778), .B1(new_n779), .B2(G159), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n778), .A2(new_n931), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n482), .B2(new_n774), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G322), .B2(new_n779), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n835), .B2(new_n935), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n770), .A2(new_n836), .B1(new_n768), .B2(new_n763), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT116), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n785), .A2(G326), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n441), .B1(new_n924), .B2(G116), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT49), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1028), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1018), .B1(new_n1043), .B2(new_n758), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n966), .A2(new_n736), .B1(new_n1011), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n966), .A2(new_n731), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n701), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n966), .A2(new_n731), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(G393));
  INV_X1    g0849(.A(new_n692), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n980), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n972), .B(new_n973), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n692), .C1(new_n977), .C2(new_n979), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1053), .A3(new_n736), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n976), .A2(new_n747), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n940), .A2(G50), .B1(new_n785), .B2(G143), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n441), .B1(new_n201), .B2(new_n763), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n770), .A2(new_n202), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n401), .C2(new_n775), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n839), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G150), .A2(new_n779), .B1(new_n778), .B2(G159), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT51), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n940), .A2(G303), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n785), .A2(G322), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n264), .B1(new_n763), .B2(new_n836), .C1(new_n774), .C2(new_n768), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G116), .B2(new_n819), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n793), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G311), .A2(new_n778), .B1(new_n779), .B2(G317), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT52), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1060), .A2(new_n1062), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n758), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n759), .B1(new_n205), .B2(new_n238), .C1(new_n754), .C2(new_n260), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1055), .A2(new_n737), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1054), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n702), .B1(new_n1075), .B2(new_n1046), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(new_n982), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT117), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(G390));
  NAND2_X1  g0879(.A1(new_n807), .A2(new_n407), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n407), .B2(new_n710), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n666), .A2(new_n710), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n806), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n726), .A2(G330), .A3(new_n808), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n859), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n726), .A2(new_n909), .A3(G330), .A4(new_n808), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT119), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT118), .B1(new_n1082), .B2(new_n806), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT118), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n864), .A2(new_n1090), .A3(new_n860), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1085), .A2(new_n1089), .A3(new_n1091), .A4(new_n1086), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1083), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(KEYINPUT119), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1088), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1086), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n896), .A2(new_n899), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n909), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n909), .B1(new_n1082), .B2(new_n806), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n898), .A2(new_n901), .B1(new_n1101), .B2(new_n899), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1097), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n898), .A2(new_n901), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n899), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n859), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1086), .C1(new_n1107), .C2(new_n1098), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n480), .A2(G330), .A3(new_n726), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n905), .A2(new_n653), .A3(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1096), .A2(new_n1103), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1095), .A2(new_n1092), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1087), .A2(KEYINPUT119), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1111), .A2(new_n1116), .A3(new_n701), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1103), .A2(new_n1108), .A3(new_n736), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT120), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1103), .A2(new_n1108), .A3(new_n1120), .A4(new_n736), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1104), .A2(new_n745), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n812), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n737), .B1(new_n1023), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n820), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n787), .A2(new_n216), .B1(new_n770), .B2(new_n424), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n785), .C2(G125), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n828), .B2(new_n835), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n264), .B1(new_n775), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(new_n826), .B2(new_n815), .C1(new_n1134), .C2(new_n829), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n818), .B1(new_n784), .B2(new_n768), .C1(new_n206), .C2(new_n835), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G116), .A2(new_n778), .B1(new_n779), .B2(G283), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1058), .B1(G97), .B2(new_n775), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n264), .B1(new_n763), .B2(new_n456), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT121), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1130), .A2(new_n1135), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n1142), .B2(new_n758), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1123), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1117), .A2(new_n1122), .A3(new_n1144), .ZN(G378));
  NAND2_X1  g0945(.A1(new_n887), .A2(new_n902), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n316), .A2(new_n675), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT55), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n340), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n1150));
  INV_X1    g0950(.A(new_n1148), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n318), .B(new_n1151), .C1(new_n338), .C2(new_n339), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n915), .B2(G330), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n740), .B(new_n1155), .C1(new_n911), .C2(new_n914), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1146), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n896), .A2(new_n726), .A3(new_n808), .A4(new_n909), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1160), .A2(KEYINPUT40), .B1(new_n912), .B2(new_n913), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1155), .B1(new_n1161), .B2(new_n740), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n915), .A2(G330), .A3(new_n1156), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n903), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n736), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n738), .B1(new_n216), .B2(new_n812), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n441), .A2(G41), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(G33), .A2(G41), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT122), .Z(new_n1169));
  AND3_X1   g0969(.A1(new_n1167), .A2(new_n216), .A3(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G125), .A2(new_n779), .B1(new_n778), .B2(G128), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n819), .A2(G150), .B1(new_n820), .B2(new_n1132), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n798), .A2(G132), .B1(new_n775), .B2(G137), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n785), .A2(G124), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1169), .B1(new_n924), .B2(G159), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1178), .C1(new_n1174), .C2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n399), .A2(new_n774), .B1(new_n766), .B2(new_n205), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT123), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n785), .A2(G283), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n787), .A2(new_n212), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n770), .A2(new_n201), .B1(new_n202), .B2(new_n763), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n1167), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G107), .A2(new_n778), .B1(new_n779), .B2(G116), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1182), .A2(new_n1183), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1176), .A2(new_n1180), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1170), .B(new_n1190), .C1(new_n1189), .C2(new_n1188), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1166), .B1(new_n814), .B2(new_n1191), .C1(new_n1155), .C2(new_n746), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1165), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT125), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1110), .B(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1115), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n906), .A2(new_n1109), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1099), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1198), .A2(new_n1199), .B1(new_n1087), .B2(KEYINPUT119), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1197), .B1(new_n1200), .B2(new_n1088), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1195), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1159), .A2(KEYINPUT57), .A3(new_n1164), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n701), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1162), .A2(new_n903), .A3(new_n1163), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n903), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1110), .A2(new_n1194), .ZN(new_n1208));
  AND4_X1   g1008(.A1(new_n1194), .A2(new_n905), .A3(new_n653), .A4(new_n1109), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1193), .B1(new_n1204), .B2(new_n1212), .ZN(G375));
  NAND3_X1  g1013(.A1(new_n1200), .A2(new_n1197), .A3(new_n1088), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1114), .A3(new_n986), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n859), .A2(new_n745), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n737), .B1(G68), .B2(new_n1124), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n940), .A2(G116), .B1(G77), .B2(new_n788), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n482), .B2(new_n784), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n386), .B(new_n1025), .C1(G97), .C2(new_n820), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G283), .A2(new_n778), .B1(new_n779), .B2(G294), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n206), .C2(new_n774), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n452), .B(new_n1184), .C1(G159), .C2(new_n820), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n775), .A2(G150), .B1(new_n819), .B2(G50), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G132), .A2(new_n779), .B1(new_n778), .B2(G137), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n835), .A2(new_n1131), .B1(new_n784), .B2(new_n1134), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1219), .A2(new_n1222), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1217), .B1(new_n1228), .B2(new_n758), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1096), .A2(new_n736), .B1(new_n1216), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1215), .A2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT126), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(G381));
  XNOR2_X1  g1033(.A(G375), .B(KEYINPUT127), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n955), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n736), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1075), .B1(new_n956), .B2(new_n1046), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n730), .B1(new_n1238), .B2(new_n967), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1239), .B2(new_n985), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1002), .A2(new_n1005), .A3(new_n1003), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1005), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1236), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1117), .A2(new_n1122), .A3(new_n1144), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1235), .A2(new_n1244), .A3(new_n1245), .A4(new_n1232), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1234), .A2(new_n1246), .ZN(G407));
  NOR2_X1   g1047(.A1(new_n673), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(new_n1234), .C2(new_n1249), .ZN(G409));
  XNOR2_X1  g1050(.A(G393), .B(new_n803), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1244), .A2(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n982), .A2(new_n1076), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1074), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1078), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(KEYINPUT117), .B(new_n1074), .C1(new_n982), .C2(new_n1076), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G387), .A2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1252), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1244), .A2(G390), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(new_n1258), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1251), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G378), .B(new_n1193), .C1(new_n1204), .C2(new_n1212), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1207), .A2(new_n1211), .A3(new_n986), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1193), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1245), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1248), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1200), .A2(new_n1197), .A3(new_n1088), .A4(KEYINPUT60), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(new_n701), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1214), .B1(new_n1201), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1274), .A2(G384), .A3(new_n1230), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G384), .B1(new_n1274), .B2(new_n1230), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1269), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1264), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1274), .A2(new_n1230), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1274), .A2(G384), .A3(new_n1230), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1248), .A2(G2897), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1269), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1277), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1280), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G2897), .B(new_n1248), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1296), .B2(new_n1269), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1248), .ZN(new_n1300));
  AND4_X1   g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .A4(new_n1277), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1269), .B2(new_n1277), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1297), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1264), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1292), .B1(new_n1303), .B2(new_n1304), .ZN(G405));
  XNOR2_X1  g1105(.A(G375), .B(G378), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1277), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1264), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1310), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1304), .A3(new_n1308), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(G402));
endmodule


