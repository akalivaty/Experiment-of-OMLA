//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT67), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n207), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n215), .B(new_n218), .C1(new_n221), .C2(new_n225), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT69), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n219), .ZN(new_n246));
  NAND3_X1  g0046(.A1(KEYINPUT69), .A2(G33), .A3(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n248), .A2(new_n252), .A3(G226), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n248), .A2(G274), .A3(new_n251), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n246), .A2(new_n243), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n255), .B1(new_n260), .B2(new_n202), .ZN(new_n261));
  MUX2_X1   g0061(.A(G222), .B(G223), .S(G1698), .Z(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n253), .A2(new_n254), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(G179), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT70), .B1(new_n266), .B2(new_n219), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G50), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n220), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n220), .B1(new_n201), .B2(new_n203), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n269), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n275), .B(new_n282), .C1(G50), .C2(new_n271), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n264), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n265), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT9), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n264), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n283), .A2(new_n287), .B1(G200), .B2(new_n264), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(new_n295), .A3(new_n292), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n286), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n255), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT75), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n258), .B2(G33), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n256), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n302));
  AND2_X1   g0102(.A1(G226), .A2(G1698), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n259), .A4(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT77), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G87), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n259), .A3(new_n302), .ZN(new_n308));
  INV_X1    g0108(.A(G1698), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n303), .A2(KEYINPUT77), .B1(G223), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n299), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n248), .A2(new_n252), .A3(G232), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n254), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n289), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n304), .A2(new_n305), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n307), .C1(new_n308), .C2(new_n310), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n314), .B1(new_n318), .B2(new_n299), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(G200), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n278), .B1(new_n270), .B2(G20), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n273), .A2(new_n321), .B1(new_n272), .B2(new_n278), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  AND2_X1   g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n203), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n276), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n308), .A2(new_n220), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(KEYINPUT7), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n301), .A2(new_n302), .A3(new_n333), .A4(new_n259), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n332), .A3(new_n220), .A4(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n323), .B(new_n327), .C1(new_n330), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT3), .B(G33), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n332), .B1(new_n337), .B2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n327), .B1(new_n340), .B2(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n269), .B1(new_n341), .B2(KEYINPUT16), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n320), .B(new_n322), .C1(new_n336), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n346));
  INV_X1    g0146(.A(new_n322), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n266), .A2(new_n219), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n340), .A2(G68), .ZN(new_n353));
  INV_X1    g0153(.A(new_n327), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n355), .B2(new_n323), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n330), .A2(new_n335), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT16), .A3(new_n354), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n347), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n312), .A2(G179), .A3(new_n315), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n284), .B1(new_n312), .B2(new_n315), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n346), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n359), .A2(KEYINPUT17), .A3(new_n320), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n322), .B1(new_n336), .B2(new_n342), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n319), .A2(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n312), .A2(new_n315), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n346), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n345), .A2(new_n363), .A3(new_n364), .A4(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n248), .A2(new_n252), .A3(G238), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G226), .A2(G1698), .ZN(new_n377));
  INV_X1    g0177(.A(G232), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(G1698), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n379), .B2(new_n337), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n254), .B(new_n374), .C1(new_n380), .C2(new_n255), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G226), .B2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n375), .B1(new_n384), .B2(new_n260), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n299), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT13), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n254), .A4(new_n374), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(G190), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n220), .A2(G33), .A3(G77), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n328), .A2(G20), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n276), .A2(G50), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n269), .B(KEYINPUT11), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n271), .A2(G68), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT12), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n396), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(new_n394), .A3(new_n393), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT11), .B1(new_n403), .B2(new_n269), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT71), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n269), .B2(new_n272), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n352), .A2(KEYINPUT71), .A3(new_n271), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G68), .A4(new_n274), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n389), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G200), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n382), .B2(new_n388), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT74), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n403), .A2(new_n269), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT11), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND4_X1   g0216(.A1(new_n409), .A2(new_n416), .A3(new_n400), .A4(new_n397), .ZN(new_n417));
  INV_X1    g0217(.A(new_n412), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n389), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n417), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n382), .A2(new_n388), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(G169), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n382), .A2(G179), .A3(new_n388), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n423), .B2(G169), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n337), .A2(G238), .A3(G1698), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n337), .A2(G232), .A3(new_n309), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n432), .C1(new_n433), .C2(new_n337), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n299), .ZN(new_n435));
  INV_X1    g0235(.A(G179), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n248), .A2(new_n252), .A3(G244), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(new_n254), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT72), .Z(new_n440));
  INV_X1    g0240(.A(new_n278), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n279), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(new_n269), .B1(new_n202), .B2(new_n272), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n407), .A2(new_n408), .A3(G77), .A4(new_n274), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n435), .A2(new_n438), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n445), .A2(new_n446), .B1(new_n447), .B2(new_n284), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(G200), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n435), .A2(G190), .A3(new_n438), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n446), .A3(new_n445), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n298), .A2(new_n373), .A3(new_n430), .A4(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(G250), .A2(G1698), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(G257), .B2(new_n309), .ZN(new_n456));
  INV_X1    g0256(.A(G294), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n308), .A2(new_n456), .B1(new_n256), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n299), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n270), .A2(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT79), .A2(G41), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(KEYINPUT5), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(KEYINPUT79), .B2(G41), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n462), .A2(new_n248), .A3(G274), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n250), .A2(G1), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n248), .A3(G264), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n411), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT88), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n474), .A3(new_n411), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n459), .A2(new_n465), .A3(new_n470), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n289), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n272), .A2(new_n433), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT25), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n270), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n352), .A2(new_n271), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n433), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n301), .A2(new_n302), .A3(new_n220), .A4(new_n259), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT22), .A2(G87), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n220), .A2(G87), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n260), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G20), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n220), .B2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n433), .A2(KEYINPUT23), .A3(G20), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n487), .A2(new_n488), .A3(new_n491), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n491), .A2(new_n497), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n485), .A2(new_n486), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT24), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n484), .B1(new_n502), .B2(new_n269), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n478), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n471), .A2(new_n284), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n469), .A2(new_n248), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n299), .A2(new_n458), .B1(new_n507), .B2(G264), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n436), .A3(new_n465), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n505), .B1(new_n510), .B2(new_n503), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n506), .A2(new_n509), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n491), .A2(new_n497), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n488), .B1(new_n513), .B2(new_n487), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT24), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n269), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n484), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n512), .A2(new_n518), .A3(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n504), .A2(new_n511), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n270), .B2(G33), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n407), .A2(new_n408), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n272), .A2(new_n521), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  AOI221_X4 g0325(.A(new_n525), .B1(new_n521), .B2(G20), .C1(new_n266), .C2(new_n219), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(G20), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT84), .B1(new_n348), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n256), .A2(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n220), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT85), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT85), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n530), .A2(new_n534), .A3(new_n220), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT20), .B1(new_n529), .B2(new_n536), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n523), .B(new_n524), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G257), .A2(G1698), .ZN(new_n541));
  INV_X1    g0341(.A(G264), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(new_n301), .A3(new_n259), .A4(new_n302), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n260), .A2(G303), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n255), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n469), .A2(new_n248), .A3(G270), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n465), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(G200), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n546), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n540), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n284), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(KEYINPUT21), .B(G169), .C1(new_n546), .C2(new_n548), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n542), .A2(G1698), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G257), .B2(G1698), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n545), .B1(new_n308), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n299), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(G179), .A3(new_n465), .A4(new_n547), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT86), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(new_n539), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n563), .B2(new_n539), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n552), .B(new_n556), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n520), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n469), .A2(new_n248), .A3(G257), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n465), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT80), .ZN(new_n571));
  INV_X1    g0371(.A(G244), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n301), .A2(new_n302), .A3(new_n573), .A4(new_n259), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT4), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n257), .A2(new_n259), .A3(G250), .A4(G1698), .ZN(new_n577));
  AND2_X1   g0377(.A1(KEYINPUT4), .A2(G244), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n257), .A2(new_n259), .A3(new_n578), .A4(new_n309), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n579), .A3(new_n531), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n299), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT80), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n465), .A2(new_n582), .A3(new_n569), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n571), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT7), .B1(new_n260), .B2(new_n220), .ZN(new_n586));
  AOI211_X1 g0386(.A(new_n332), .B(G20), .C1(new_n257), .C2(new_n259), .ZN(new_n587));
  OAI21_X1  g0387(.A(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT6), .ZN(new_n589));
  AND2_X1   g0389(.A1(G97), .A2(G107), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n433), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n352), .B1(new_n588), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G97), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n483), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n271), .A2(G97), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n465), .A2(new_n569), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n581), .A2(new_n601), .A3(G190), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT81), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT81), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n581), .A2(new_n601), .A3(new_n604), .A4(G190), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n585), .A2(new_n600), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n598), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n594), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n276), .A2(G77), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n433), .B1(new_n338), .B2(new_n339), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n269), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n599), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n581), .A2(new_n601), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n284), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n571), .A2(new_n581), .A3(new_n583), .A4(new_n436), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(G250), .B1(new_n270), .B2(G45), .ZN(new_n620));
  INV_X1    g0420(.A(G274), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n468), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n572), .A2(G1698), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(G238), .B2(G1698), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n492), .B1(new_n308), .B2(new_n624), .ZN(new_n625));
  AOI221_X4 g0425(.A(G179), .B1(new_n622), .B2(new_n248), .C1(new_n625), .C2(new_n299), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n299), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(new_n248), .ZN(new_n628));
  AOI21_X1  g0428(.A(G169), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n485), .A2(new_n328), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT19), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n632), .A2(new_n220), .A3(G33), .A4(G97), .ZN(new_n633));
  INV_X1    g0433(.A(G87), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n597), .A3(new_n433), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n375), .A2(new_n220), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n637), .B2(KEYINPUT19), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n269), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n443), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n271), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n352), .A2(new_n271), .A3(new_n640), .A4(new_n482), .ZN(new_n643));
  AND4_X1   g0443(.A1(KEYINPUT82), .A2(new_n639), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n645), .A2(new_n633), .B1(new_n485), .B2(new_n328), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n641), .B1(new_n646), .B2(new_n269), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT82), .B1(new_n647), .B2(new_n643), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n630), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n627), .A2(G190), .A3(new_n628), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n411), .B1(new_n627), .B2(new_n628), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n273), .A2(G87), .A3(new_n482), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT83), .B1(new_n619), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n606), .A2(new_n618), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT83), .ZN(new_n660));
  INV_X1    g0460(.A(new_n657), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n454), .A2(new_n568), .A3(new_n658), .A4(new_n662), .ZN(G372));
  AND2_X1   g0463(.A1(new_n345), .A2(new_n364), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n449), .B1(new_n420), .B2(new_n413), .ZN(new_n665));
  INV_X1    g0465(.A(new_n429), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT91), .B1(new_n359), .B2(new_n362), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT91), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n365), .A2(new_n369), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(KEYINPUT18), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n294), .A2(new_n296), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n286), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n454), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n627), .A2(new_n436), .A3(new_n628), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n625), .A2(new_n299), .B1(new_n248), .B2(new_n622), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(G169), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT82), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n647), .A2(KEYINPUT82), .A3(new_n643), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n654), .A2(new_n650), .A3(new_n651), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT89), .B1(new_n649), .B2(new_n656), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n472), .A2(KEYINPUT88), .B1(new_n476), .B2(new_n289), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n518), .B1(new_n475), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n619), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n649), .A2(KEYINPUT89), .A3(new_n656), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n471), .A2(new_n474), .A3(new_n411), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n474), .B1(new_n471), .B2(new_n411), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n471), .A2(G190), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n618), .B(new_n606), .C1(new_n704), .C2(new_n518), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT90), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n563), .A2(new_n539), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n556), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n510), .A2(new_n503), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n697), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n649), .A3(new_n656), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n687), .B1(new_n714), .B2(KEYINPUT26), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT26), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n698), .A2(new_n699), .A3(new_n716), .A4(new_n713), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n678), .B1(new_n679), .B2(new_n720), .ZN(G369));
  NAND3_X1  g0521(.A1(new_n270), .A2(new_n220), .A3(G13), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G213), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT92), .B(G343), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n709), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT93), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n503), .A2(new_n728), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n520), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n520), .B2(new_n731), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(new_n709), .B2(new_n727), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n707), .A2(KEYINPUT86), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n563), .A2(new_n539), .A3(new_n564), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n556), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n728), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n729), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n540), .A2(new_n728), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n708), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n567), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n734), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n741), .A2(new_n747), .ZN(G399));
  NAND3_X1  g0548(.A1(new_n216), .A2(KEYINPUT95), .A3(new_n249), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT95), .B1(new_n216), .B2(new_n249), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n591), .A2(new_n634), .A3(new_n521), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n752), .A2(new_n270), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n225), .B2(new_n752), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  AOI211_X1 g0556(.A(KEYINPUT29), .B(new_n727), .C1(new_n712), .C2(new_n719), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT29), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n737), .A2(new_n511), .A3(new_n519), .A4(new_n556), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n692), .A3(new_n695), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n692), .A2(KEYINPUT97), .A3(KEYINPUT26), .A4(new_n713), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT97), .B1(new_n714), .B2(new_n716), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT26), .A4(new_n713), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n760), .A2(new_n761), .A3(new_n764), .A4(new_n649), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n758), .B1(new_n765), .B2(new_n728), .ZN(new_n766));
  INV_X1    g0566(.A(G330), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n550), .A2(G179), .A3(new_n508), .A4(new_n681), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT96), .B1(new_n768), .B2(new_n615), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT30), .ZN(new_n771));
  OAI211_X1 g0571(.A(KEYINPUT96), .B(new_n771), .C1(new_n768), .C2(new_n615), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n550), .A2(G179), .A3(new_n681), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n471), .A3(new_n584), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  AND3_X1   g0575(.A1(new_n775), .A2(KEYINPUT31), .A3(new_n727), .ZN(new_n776));
  AOI21_X1  g0576(.A(KEYINPUT31), .B1(new_n775), .B2(new_n727), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n568), .A2(new_n658), .A3(new_n662), .A4(new_n728), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n767), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n757), .A2(new_n766), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n756), .B1(new_n781), .B2(G1), .ZN(G364));
  AND2_X1   g0582(.A1(new_n220), .A2(G13), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n270), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n752), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n744), .B2(G330), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G330), .B2(new_n744), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n219), .B1(G20), .B2(new_n284), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n220), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT99), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n793), .A2(G179), .A3(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT32), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n220), .A2(new_n289), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n436), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n791), .A2(new_n798), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G58), .A2(new_n800), .B1(new_n802), .B2(G77), .ZN(new_n803));
  INV_X1    g0603(.A(G50), .ZN(new_n804));
  NAND3_X1  g0604(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n289), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n803), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT98), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G179), .A2(G200), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n220), .B1(new_n810), .B2(G190), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n597), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n797), .A2(new_n436), .A3(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n805), .A2(G190), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n337), .B1(new_n813), .B2(new_n634), .C1(new_n328), .C2(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n793), .A2(G179), .A3(new_n411), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n812), .B(new_n816), .C1(G107), .C2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n796), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n794), .A2(G329), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(G283), .ZN(new_n821));
  INV_X1    g0621(.A(new_n813), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n337), .B1(new_n822), .B2(G303), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G322), .A2(new_n800), .B1(new_n802), .B2(G311), .ZN(new_n824));
  AND4_X1   g0624(.A1(new_n820), .A2(new_n821), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n811), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(G294), .B1(G326), .B2(new_n806), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT33), .B(G317), .Z(new_n828));
  OAI211_X1 g0628(.A(new_n825), .B(new_n827), .C1(new_n815), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n790), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n216), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n260), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G355), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(G116), .B2(new_n216), .ZN(new_n834));
  MUX2_X1   g0634(.A(new_n224), .B(new_n241), .S(G45), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n331), .A2(new_n334), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(G13), .A2(G33), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G20), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n789), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n786), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n830), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n841), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n744), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n788), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  INV_X1    g0649(.A(new_n786), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n789), .A2(new_n839), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n202), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n812), .B1(new_n806), .B2(G303), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n815), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n813), .A2(new_n433), .B1(new_n799), .B2(new_n457), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n337), .B(new_n856), .C1(G116), .C2(new_n802), .ZN(new_n857));
  INV_X1    g0657(.A(new_n817), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n634), .B2(new_n858), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n855), .B(new_n859), .C1(G311), .C2(new_n794), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n817), .A2(G68), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n794), .A2(G132), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n822), .A2(G50), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n826), .A2(G58), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n836), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT100), .ZN(new_n868));
  AOI22_X1  g0668(.A1(G143), .A2(new_n800), .B1(new_n802), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(new_n815), .B2(new_n870), .C1(new_n871), .C2(new_n807), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT34), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n860), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n440), .A2(new_n448), .A3(new_n728), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n445), .A2(new_n446), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n727), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n440), .A2(new_n448), .B1(new_n452), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n852), .B1(new_n874), .B2(new_n790), .C1(new_n880), .C2(new_n840), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n452), .A2(new_n878), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n449), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n875), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n720), .B2(new_n727), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n712), .A2(new_n719), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n728), .A3(new_n880), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(KEYINPUT101), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT101), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n885), .C1(new_n720), .C2(new_n727), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n780), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(KEYINPUT102), .A3(new_n780), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n780), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n889), .A2(new_n898), .A3(new_n891), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n850), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n882), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(G384));
  OR2_X1    g0703(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(G116), .A3(new_n221), .A4(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT36), .Z(new_n907));
  OR3_X1    g0707(.A1(new_n224), .A2(new_n202), .A3(new_n324), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n201), .A2(G68), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n270), .B(G13), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n422), .A2(new_n727), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n421), .A2(new_n429), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n421), .B2(new_n429), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n888), .B2(new_n875), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n327), .B1(new_n330), .B2(new_n335), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n269), .B1(new_n918), .B2(KEYINPUT16), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n336), .B1(new_n919), .B2(KEYINPUT103), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n269), .C1(new_n918), .C2(KEYINPUT16), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n347), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n725), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n369), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n343), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n359), .B2(new_n725), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n365), .A2(KEYINPUT104), .A3(new_n924), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n365), .A2(new_n369), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT37), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n343), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n926), .A2(KEYINPUT37), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n923), .A2(new_n725), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n373), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n917), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n373), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n358), .A3(new_n922), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n322), .ZN(new_n941));
  INV_X1    g0741(.A(new_n925), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n932), .B1(new_n943), .B2(new_n343), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n343), .A2(new_n931), .A3(new_n932), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n928), .B2(new_n929), .ZN(new_n946));
  OAI211_X1 g0746(.A(KEYINPUT38), .B(new_n938), .C1(new_n944), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n916), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n343), .A2(KEYINPUT105), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT105), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n359), .A2(new_n952), .A3(new_n320), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n359), .A2(new_n362), .A3(KEYINPUT91), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n669), .B1(new_n365), .B2(new_n369), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n951), .B(new_n953), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n928), .A2(new_n929), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT37), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n946), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n668), .A2(KEYINPUT18), .A3(new_n670), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT18), .B1(new_n668), .B2(new_n670), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n664), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n957), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT38), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n947), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n950), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n666), .A2(new_n728), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n937), .A2(new_n947), .A3(KEYINPUT39), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n673), .A2(new_n674), .A3(new_n725), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n949), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n454), .B1(new_n757), .B2(new_n766), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n678), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n914), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n421), .A2(new_n429), .A3(new_n912), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n885), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT106), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT40), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND4_X1   g0782(.A1(new_n568), .A2(new_n658), .A3(new_n662), .A4(new_n728), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n775), .A2(new_n727), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT31), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n775), .A2(KEYINPUT31), .A3(new_n727), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n979), .B(new_n982), .C1(new_n983), .C2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n880), .B1(new_n913), .B2(new_n914), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n779), .B2(new_n778), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n948), .C1(KEYINPUT106), .C2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n979), .B1(new_n983), .B2(new_n988), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n930), .B1(new_n675), .B2(new_n664), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n671), .A2(new_n930), .A3(new_n953), .A4(new_n951), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n946), .B1(new_n995), .B2(KEYINPUT37), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n917), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n993), .B1(new_n947), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n992), .B1(new_n998), .B2(new_n981), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n679), .B1(new_n779), .B2(new_n778), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n767), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n999), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n976), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n270), .B2(new_n783), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n976), .A2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n911), .B1(new_n1004), .B2(new_n1005), .ZN(G367));
  NOR2_X1   g0806(.A1(new_n618), .A2(new_n728), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT107), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n659), .B1(new_n600), .B2(new_n728), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n734), .A2(new_n740), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n519), .A2(new_n511), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n618), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1013), .A2(KEYINPUT42), .B1(new_n728), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n655), .A2(new_n728), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n700), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n687), .A2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(KEYINPUT43), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1019), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1016), .A2(new_n1025), .A3(new_n1024), .A4(new_n1018), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n746), .A2(new_n1011), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1030), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n752), .B(KEYINPUT41), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n734), .A2(new_n745), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n746), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n740), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n740), .B1(new_n746), .B2(new_n1035), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n781), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n741), .A2(KEYINPUT44), .A3(new_n1011), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT44), .B1(new_n741), .B2(new_n1011), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n729), .B(new_n1010), .C1(new_n734), .C2(new_n740), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n747), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1047), .B(KEYINPUT45), .Z(new_n1050));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n1043), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1052), .A3(new_n746), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1042), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1034), .B1(new_n1054), .B2(new_n781), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1033), .B1(new_n1055), .B2(new_n785), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n837), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n842), .B1(new_n216), .B2(new_n443), .C1(new_n1057), .C2(new_n234), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n786), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n799), .A2(new_n870), .B1(new_n801), .B2(new_n201), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n260), .B(new_n1060), .C1(G58), .C2(new_n822), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n817), .A2(G77), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n794), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT108), .B(G137), .Z(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n826), .A2(G68), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n806), .A2(G143), .ZN(new_n1067));
  INV_X1    g0867(.A(G159), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1067), .C1(new_n1068), .C2(new_n815), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n794), .A2(G317), .ZN(new_n1070));
  INV_X1    g0870(.A(G303), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n799), .A2(new_n1071), .B1(new_n801), .B2(new_n854), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G107), .B2(new_n826), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n858), .C2(new_n597), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n813), .A2(new_n521), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT46), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G294), .B2(new_n814), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1075), .A2(KEYINPUT46), .B1(new_n806), .B2(G311), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n866), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1065), .A2(new_n1069), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT47), .Z(new_n1081));
  OAI221_X1 g0881(.A(new_n1059), .B1(new_n790), .B2(new_n1081), .C1(new_n1023), .C2(new_n846), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1056), .A2(new_n1082), .ZN(G387));
  INV_X1    g0883(.A(KEYINPUT112), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n781), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n781), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1040), .A2(KEYINPUT112), .A3(new_n1041), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n752), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n811), .A2(new_n443), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n822), .A2(G77), .B1(new_n800), .B2(G50), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n328), .B2(new_n801), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(new_n441), .C2(new_n814), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT109), .B(G150), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n817), .A2(G97), .B1(new_n794), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n806), .A2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT110), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n836), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n814), .A2(G311), .B1(new_n806), .B2(G322), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT111), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT111), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G317), .A2(new_n800), .B1(new_n802), .B2(G303), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT48), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n813), .A2(new_n457), .B1(new_n811), .B2(new_n854), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G116), .A2(new_n817), .B1(new_n794), .B2(G326), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n866), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT49), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1098), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n789), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n231), .A2(new_n250), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1114), .A2(new_n837), .B1(new_n753), .B2(new_n832), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT50), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n441), .B2(new_n804), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n278), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n250), .B1(new_n328), .B2(new_n202), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n753), .A4(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1115), .A2(new_n1120), .B1(G107), .B2(new_n216), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n842), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1113), .A2(new_n1122), .A3(new_n786), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n734), .B2(new_n841), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1085), .B2(new_n785), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1089), .A2(new_n1125), .ZN(G393));
  NAND2_X1  g0926(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1087), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(new_n752), .A3(new_n1054), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1049), .A2(new_n1053), .A3(new_n785), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n842), .B1(new_n597), .B2(new_n216), .C1(new_n1057), .C2(new_n238), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n786), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n800), .A2(G311), .B1(G317), .B2(new_n806), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G107), .A2(new_n817), .B1(new_n794), .B2(G322), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n260), .B1(new_n801), .B2(new_n457), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G283), .B2(new_n822), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n826), .A2(G116), .B1(G303), .B2(new_n814), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G87), .A2(new_n817), .B1(new_n794), .B2(G143), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n811), .A2(new_n202), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n813), .A2(new_n328), .B1(new_n801), .B2(new_n278), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n201), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1142), .C1(new_n1143), .C2(new_n814), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n836), .A3(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n800), .A2(G159), .B1(G150), .B2(new_n806), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT51), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1134), .A2(new_n1139), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1132), .B1(new_n1148), .B2(new_n789), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1010), .B2(new_n846), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1130), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1129), .A2(new_n1151), .ZN(G390));
  INV_X1    g0952(.A(new_n915), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n780), .A2(new_n880), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n727), .B(new_n885), .C1(new_n712), .C2(new_n719), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1153), .B1(new_n1156), .B2(new_n876), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1157), .A2(new_n968), .B1(new_n967), .B2(new_n970), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n997), .A2(new_n947), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n968), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n765), .A2(new_n728), .A3(new_n884), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n915), .B1(new_n1161), .B2(new_n875), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1155), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n969), .B1(new_n997), .B2(new_n947), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1161), .A2(new_n875), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n915), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n916), .A2(new_n969), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n970), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1159), .B2(new_n950), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1154), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1164), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1170), .A2(new_n840), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n851), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n786), .B1(new_n441), .B2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n260), .B1(new_n799), .B2(new_n521), .C1(new_n634), .C2(new_n813), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1141), .B(new_n1177), .C1(G283), .C2(new_n806), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n794), .A2(G294), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n802), .A2(G97), .B1(G107), .B2(new_n814), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT118), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n861), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT54), .B(G143), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n801), .A2(new_n1183), .B1(new_n811), .B2(new_n1068), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1064), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n814), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT116), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G125), .A2(new_n794), .B1(new_n817), .B2(new_n1143), .ZN(new_n1188));
  INV_X1    g0988(.A(G132), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n337), .B1(new_n799), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G128), .B2(new_n806), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n822), .A2(new_n1094), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1188), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1182), .B1(new_n1187), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1176), .B1(new_n1196), .B2(new_n789), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1173), .A2(new_n785), .B1(new_n1174), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n752), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n888), .A2(new_n875), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1153), .B1(new_n780), .B2(new_n880), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n1155), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n780), .A2(new_n880), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n915), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1166), .A2(new_n1204), .A3(new_n1154), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT114), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n454), .A2(new_n780), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n974), .A2(new_n678), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT113), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT113), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n974), .A2(new_n1211), .A3(new_n678), .A4(new_n1208), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1155), .A2(new_n1201), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(KEYINPUT114), .A3(new_n1166), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1207), .A2(new_n1210), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1199), .B1(new_n1172), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AND4_X1   g1018(.A1(KEYINPUT114), .A2(new_n1166), .A3(new_n1204), .A4(new_n1154), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT114), .B1(new_n1213), .B2(new_n1166), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n1202), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1221), .A3(new_n1164), .A4(new_n1171), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1216), .A2(new_n1222), .A3(KEYINPUT115), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT115), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1198), .B1(new_n1223), .B2(new_n1224), .ZN(G378));
  NAND2_X1  g1025(.A1(new_n1207), .A2(new_n1214), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1218), .B1(new_n1172), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n283), .A2(new_n924), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n297), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n297), .A2(new_n1228), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n991), .B1(new_n965), .B2(new_n966), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT40), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n767), .B(new_n1234), .C1(new_n1236), .C2(new_n992), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1234), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n999), .B2(G330), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n973), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n993), .A2(new_n980), .B1(new_n947), .B2(new_n937), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n989), .A2(new_n1241), .B1(new_n1235), .B2(KEYINPUT40), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1234), .B1(new_n1242), .B2(new_n767), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n949), .A2(new_n971), .A3(new_n972), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n999), .A2(G330), .A3(new_n1238), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1227), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT119), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1240), .A2(new_n1246), .A3(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT119), .A4(new_n1245), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1227), .A3(KEYINPUT57), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n752), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1234), .A2(new_n839), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n786), .B1(new_n1143), .B2(new_n1175), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n815), .A2(new_n1189), .B1(new_n811), .B2(new_n870), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n800), .A2(G128), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n871), .B2(new_n801), .C1(new_n813), .C2(new_n1183), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G125), .C2(new_n806), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n256), .B(new_n249), .C1(new_n858), .C2(new_n1068), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G124), .B2(new_n794), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n817), .A2(G58), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n799), .A2(new_n433), .B1(new_n801), .B2(new_n443), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n249), .B1(new_n813), .B2(new_n202), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1268), .B(new_n1271), .C1(new_n1063), .C2(new_n854), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1066), .B1(new_n815), .B2(new_n597), .C1(new_n521), .C2(new_n807), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1272), .A2(new_n836), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT58), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(KEYINPUT58), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n249), .B1(new_n866), .B2(new_n256), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n804), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1267), .A2(new_n1275), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1257), .B1(new_n1279), .B2(new_n789), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1247), .A2(new_n785), .B1(new_n1256), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1255), .A2(new_n1281), .ZN(G375));
  AOI21_X1  g1082(.A(new_n1034), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1226), .A2(new_n1217), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n786), .B1(G68), .B2(new_n1175), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1090), .B1(new_n806), .B2(G294), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n521), .B2(new_n815), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n794), .A2(G303), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n337), .B1(new_n822), .B2(G97), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(G283), .A2(new_n800), .B1(new_n802), .B2(G107), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1062), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n794), .A2(G128), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1185), .A2(new_n800), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n822), .A2(G159), .B1(new_n802), .B2(G150), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1268), .A2(new_n1293), .A3(new_n1294), .A4(new_n1295), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n826), .A2(G50), .B1(G132), .B2(new_n806), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n836), .B(new_n1297), .C1(new_n815), .C2(new_n1183), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n1288), .A2(new_n1292), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1286), .B1(new_n789), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1153), .B2(new_n840), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1226), .B2(new_n784), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1285), .A2(new_n1302), .ZN(G381));
  NAND3_X1  g1103(.A1(new_n1089), .A2(new_n848), .A3(new_n1125), .ZN(new_n1304));
  OR3_X1    g1104(.A1(G390), .A2(G384), .A3(new_n1304), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1305), .A2(G387), .A3(G381), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(new_n1198), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1306), .A2(new_n1255), .A3(new_n1281), .A4(new_n1308), .ZN(G407));
  NAND2_X1  g1109(.A1(new_n726), .A2(G213), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G407), .B(G213), .C1(G375), .C2(new_n1312), .ZN(G409));
  XOR2_X1   g1113(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1314));
  NAND3_X1  g1114(.A1(G378), .A2(new_n1255), .A3(new_n1281), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1252), .A2(new_n785), .A3(new_n1253), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1256), .A2(new_n1280), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1316), .B(new_n1317), .C1(new_n1034), .C2(new_n1248), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1308), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1315), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1310), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(G2897), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT122), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1322), .A2(KEYINPUT122), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT120), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1302), .B1(new_n902), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1215), .A2(KEYINPUT60), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1284), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1226), .A2(new_n1217), .A3(KEYINPUT60), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n752), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n1331));
  OAI21_X1  g1131(.A(KEYINPUT120), .B1(new_n1331), .B2(new_n882), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1326), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1326), .B2(new_n1330), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1323), .B(new_n1324), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1326), .A2(new_n1330), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1332), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1326), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1338), .A2(KEYINPUT122), .A3(new_n1322), .A4(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1314), .B1(new_n1321), .B2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1311), .B1(new_n1315), .B2(new_n1319), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1343), .A2(KEYINPUT62), .A3(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT62), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1342), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT126), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(G393), .A2(G396), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1304), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(KEYINPUT123), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1056), .A2(new_n1082), .A3(G390), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT124), .ZN(new_n1354));
  AOI21_X1  g1154(.A(G390), .B1(new_n1056), .B2(new_n1082), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1353), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1355), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(KEYINPUT124), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1352), .B1(new_n1356), .B2(new_n1358), .ZN(new_n1359));
  AOI211_X1 g1159(.A(new_n1355), .B(new_n1353), .C1(new_n1304), .C2(new_n1350), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1342), .B(KEYINPUT126), .C1(new_n1345), .C2(new_n1346), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1349), .A2(new_n1361), .A3(new_n1362), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1361), .A2(KEYINPUT61), .ZN(new_n1364));
  AOI22_X1  g1164(.A1(new_n1343), .A2(KEYINPUT121), .B1(new_n1340), .B2(new_n1335), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1365), .B1(KEYINPUT121), .B2(new_n1343), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(KEYINPUT63), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1367), .A2(KEYINPUT63), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1364), .A2(new_n1366), .A3(new_n1368), .A4(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1363), .A2(new_n1370), .ZN(G405));
  NOR2_X1   g1171(.A1(new_n1344), .A2(KEYINPUT127), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1361), .A2(new_n1373), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1372), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1344), .A2(KEYINPUT127), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(G375), .A2(new_n1308), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1377), .A2(new_n1315), .A3(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1376), .A2(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(new_n1379), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1374), .A2(new_n1381), .A3(new_n1375), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1380), .A2(new_n1382), .ZN(G402));
endmodule


