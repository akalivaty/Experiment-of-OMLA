//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1323, new_n1324, new_n1325, new_n1326, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n209), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT0), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n211), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n218), .A2(KEYINPUT0), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n219), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n206), .C2(new_n217), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n213), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n228), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n211), .A2(new_n255), .A3(KEYINPUT69), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G20), .B2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n259), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT8), .A2(G58), .ZN(new_n261));
  INV_X1    g0061(.A(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n261), .B1(new_n266), .B2(KEYINPUT8), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n211), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n260), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n223), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G20), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n272), .B1(new_n210), .B2(G20), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(G50), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(KEYINPUT9), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(KEYINPUT9), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n255), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G222), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(new_n230), .B2(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(G1698), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT67), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n292), .B1(new_n294), .B2(G223), .ZN(new_n295));
  AND2_X1   g0095(.A1(G1), .A2(G13), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G226), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n296), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT66), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n210), .C1(G41), .C2(G45), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT10), .B1(new_n310), .B2(G190), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT70), .B(G200), .Z(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n299), .B2(new_n309), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n281), .A2(new_n315), .A3(new_n282), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n284), .A2(new_n311), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OR3_X1    g0118(.A1(new_n299), .A2(new_n318), .A3(new_n309), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n283), .A3(new_n314), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n259), .A2(G50), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n259), .A2(KEYINPUT73), .A3(G50), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n269), .A2(new_n230), .B1(new_n211), .B2(G68), .ZN(new_n328));
  OAI211_X1 g0128(.A(KEYINPUT11), .B(new_n272), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n325), .B2(new_n326), .ZN(new_n331));
  INV_X1    g0131(.A(new_n272), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OR3_X1    g0133(.A1(new_n276), .A2(KEYINPUT12), .A3(G68), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT12), .B1(new_n276), .B2(G68), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(G68), .B2(new_n278), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n329), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n240), .A2(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(G226), .B2(G1698), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n338), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n298), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n301), .A2(G238), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n308), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n344), .A2(new_n345), .B1(new_n301), .B2(G238), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n308), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n352), .A3(G190), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n352), .A3(KEYINPUT72), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT72), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n350), .A2(new_n356), .A3(new_n351), .A4(new_n308), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n355), .A2(G200), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(G169), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT14), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n355), .A2(new_n362), .A3(G169), .A4(new_n357), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n349), .A2(new_n352), .A3(G179), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n337), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n299), .A2(G179), .A3(new_n309), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n280), .C1(G169), .C2(new_n310), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n278), .A2(G77), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G77), .B2(new_n276), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G20), .A2(G77), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT8), .B(G58), .Z(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n259), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n373), .B1(new_n269), .B2(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n372), .B1(new_n272), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n301), .A2(G244), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n380), .A2(new_n308), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n290), .A2(new_n240), .B1(new_n206), .B2(new_n288), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n294), .B2(G238), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n383), .B2(new_n298), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n379), .B1(new_n384), .B2(new_n318), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT67), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n293), .B(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G238), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n345), .B1(new_n389), .B2(new_n382), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n312), .B1(new_n390), .B2(new_n381), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n379), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G179), .B2(new_n384), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n322), .A2(new_n367), .A3(new_n370), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n298), .A2(G232), .A3(new_n300), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n308), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(G223), .A2(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G226), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(G1698), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n288), .B1(G33), .B2(G87), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n345), .B1(new_n405), .B2(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n407), .B1(new_n410), .B2(new_n343), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n318), .B(new_n401), .C1(new_n406), .C2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n298), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n405), .A2(KEYINPUT76), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n400), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(G200), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n268), .A2(new_n278), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n268), .A2(new_n276), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n286), .A2(new_n211), .A3(new_n287), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n287), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT75), .B1(new_n426), .B2(G68), .ZN(new_n427));
  INV_X1    g0227(.A(G68), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n263), .B2(new_n265), .ZN(new_n429));
  OAI21_X1  g0229(.A(G20), .B1(new_n429), .B2(new_n201), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT74), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n259), .B2(G159), .ZN(new_n432));
  INV_X1    g0232(.A(G159), .ZN(new_n433));
  AOI211_X1 g0233(.A(KEYINPUT74), .B(new_n433), .C1(new_n256), .C2(new_n258), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n428), .B1(new_n424), .B2(new_n425), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT75), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT16), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n259), .A2(G159), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT74), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n259), .A2(new_n431), .A3(G159), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT7), .B1(new_n343), .B2(new_n211), .ZN(new_n444));
  INV_X1    g0244(.A(new_n425), .ZN(new_n445));
  OAI21_X1  g0245(.A(G68), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(KEYINPUT16), .A3(new_n446), .A4(new_n430), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n272), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n418), .B(new_n421), .C1(new_n439), .C2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n398), .B1(new_n449), .B2(KEYINPUT77), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT68), .B(G58), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n220), .B1(new_n453), .B2(new_n428), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n441), .A2(new_n442), .B1(G20), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n455), .A3(new_n438), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT16), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n435), .A2(new_n437), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n332), .B1(new_n459), .B2(KEYINPUT16), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n458), .A2(new_n460), .B1(new_n420), .B2(new_n419), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n415), .A2(new_n416), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n393), .B1(new_n462), .B2(new_n401), .ZN(new_n463));
  INV_X1    g0263(.A(G179), .ZN(new_n464));
  AOI211_X1 g0264(.A(new_n464), .B(new_n400), .C1(new_n415), .C2(new_n416), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT18), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT77), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n461), .A2(new_n468), .A3(KEYINPUT17), .A4(new_n418), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n421), .B1(new_n439), .B2(new_n448), .ZN(new_n470));
  INV_X1    g0270(.A(new_n466), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT18), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n450), .A2(new_n467), .A3(new_n469), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n397), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n476));
  XNOR2_X1  g0276(.A(G97), .B(G107), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n479), .A2(new_n211), .B1(new_n377), .B2(new_n230), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n206), .B1(new_n424), .B2(new_n425), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n272), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n276), .A2(G97), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n210), .A2(KEYINPUT78), .A3(G33), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n255), .B2(G1), .ZN(new_n486));
  AND4_X1   g0286(.A1(new_n332), .A2(new_n276), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n487), .B2(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G257), .A3(new_n298), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT80), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n495), .A2(new_n498), .A3(G257), .A4(new_n298), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G244), .B(new_n289), .C1(new_n341), .C2(new_n342), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G250), .A2(G1698), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT4), .A2(G244), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G1698), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n288), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n345), .ZN(new_n511));
  AND2_X1   g0311(.A1(G33), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(G274), .B1(new_n512), .B2(new_n223), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT79), .B1(new_n495), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n210), .A2(G45), .ZN(new_n515));
  OR2_X1    g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n492), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n304), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n500), .A2(new_n511), .A3(new_n464), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n489), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n510), .A2(new_n345), .B1(new_n519), .B2(new_n514), .ZN(new_n523));
  AOI21_X1  g0323(.A(G169), .B1(new_n523), .B2(new_n500), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT81), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n500), .A2(new_n511), .A3(new_n520), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n393), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n489), .A4(new_n521), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n482), .A2(new_n488), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(G200), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n318), .C2(new_n526), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n525), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G200), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n495), .A2(new_n513), .A3(KEYINPUT79), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n518), .B1(new_n517), .B2(new_n304), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n495), .A2(G264), .A3(new_n298), .ZN(new_n538));
  INV_X1    g0338(.A(G294), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n255), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G250), .A2(G1698), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n216), .B2(G1698), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(new_n288), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n538), .B1(new_n543), .B2(new_n298), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n534), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n216), .A2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G250), .B2(G1698), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n343), .B1(new_n255), .B2(new_n539), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n516), .A2(new_n492), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(new_n491), .B1(new_n296), .B2(new_n297), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n548), .A2(new_n345), .B1(new_n550), .B2(G264), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n520), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n545), .B1(new_n552), .B2(G190), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n487), .A2(G107), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n211), .A2(G107), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n275), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(KEYINPUT87), .A3(KEYINPUT25), .ZN(new_n557));
  OR2_X1    g0357(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g0358(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n275), .A2(new_n555), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n288), .A2(new_n563), .A3(new_n211), .A4(G87), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n211), .B(G87), .C1(new_n341), .C2(new_n342), .ZN(new_n565));
  XOR2_X1   g0365(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT85), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(G20), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n211), .A2(KEYINPUT85), .A3(G33), .A4(G116), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n211), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n571), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(KEYINPUT86), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT86), .B1(new_n568), .B2(new_n576), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n568), .A2(new_n576), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n272), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n553), .B(new_n562), .C1(new_n581), .C2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n374), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n276), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n288), .A2(new_n211), .A3(G68), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n211), .B1(new_n338), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(G87), .B2(new_n207), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n269), .B2(new_n205), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n588), .B1(new_n594), .B2(new_n272), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n487), .A2(new_n587), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n231), .A2(G1698), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G238), .B2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n570), .B1(new_n599), .B2(new_n343), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n345), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n210), .A2(new_n303), .A3(G45), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n209), .B1(new_n490), .B2(G1), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n298), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n393), .ZN(new_n606));
  INV_X1    g0406(.A(new_n604), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n600), .B2(new_n345), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n464), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n597), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n313), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(G190), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n487), .A2(G87), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n595), .A4(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n586), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n533), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NOR2_X1   g0418(.A1(G257), .A2(G1698), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n217), .B2(G1698), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n286), .B2(new_n287), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n345), .B1(new_n288), .B2(G303), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n495), .A2(G270), .A3(new_n298), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n535), .B2(new_n536), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT82), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n520), .A2(KEYINPUT82), .A3(new_n624), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G116), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n276), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n487), .B2(new_n630), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n504), .B(new_n211), .C1(G33), .C2(new_n205), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT20), .ZN(new_n634));
  AOI22_X1  g0434(.A1(KEYINPUT83), .A2(new_n634), .B1(new_n630), .B2(G20), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n635), .A3(new_n272), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n634), .A2(KEYINPUT83), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G169), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n618), .B1(new_n629), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n629), .A2(G179), .A3(new_n639), .ZN(new_n642));
  INV_X1    g0442(.A(new_n623), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n520), .A2(KEYINPUT82), .A3(new_n624), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT82), .B1(new_n520), .B2(new_n624), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n393), .B1(new_n632), .B2(new_n638), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(KEYINPUT21), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT88), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n650), .B(G169), .C1(new_n537), .C2(new_n544), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n551), .A2(G179), .A3(new_n520), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n650), .B1(new_n552), .B2(G169), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n582), .A2(new_n583), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n577), .A3(KEYINPUT24), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n332), .B1(new_n579), .B2(new_n580), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n561), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n629), .A2(G190), .ZN(new_n662));
  INV_X1    g0462(.A(new_n639), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n662), .B(new_n663), .C1(new_n534), .C2(new_n629), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n475), .A2(new_n617), .A3(new_n661), .A4(new_n664), .ZN(G372));
  NAND2_X1  g0465(.A1(new_n467), .A2(new_n473), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n365), .A2(new_n366), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n359), .B2(new_n395), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n450), .A2(new_n469), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n322), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n370), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n475), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT89), .B1(new_n649), .B2(new_n660), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n617), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n661), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT90), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n525), .A2(new_n529), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n615), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n522), .A2(new_n524), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n615), .A2(new_n684), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n610), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n680), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n610), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n610), .A2(new_n614), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n527), .A2(new_n489), .A3(new_n521), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n688), .B1(new_n691), .B2(new_n681), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n525), .B2(new_n529), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n692), .B(KEYINPUT90), .C1(new_n681), .C2(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n677), .A2(new_n679), .B1(new_n687), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n674), .B1(new_n675), .B2(new_n695), .ZN(G369));
  OAI21_X1  g0496(.A(new_n562), .B1(new_n581), .B2(new_n585), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n654), .B2(new_n653), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n275), .A2(new_n211), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  OAI21_X1  g0500(.A(G213), .B1(new_n699), .B2(KEYINPUT27), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n703), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G343), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n649), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n586), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n659), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n698), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n706), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n664), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n705), .A2(new_n639), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n649), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n641), .A2(new_n715), .A3(new_n642), .A4(new_n648), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(KEYINPUT92), .A3(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n660), .A2(new_n708), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n712), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT93), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT93), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n729), .B(new_n726), .C1(new_n722), .C2(new_n723), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n713), .B1(new_n728), .B2(new_n730), .ZN(G399));
  INV_X1    g0531(.A(G41), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n214), .A2(KEYINPUT94), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT94), .B1(new_n214), .B2(new_n732), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n222), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n737), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  INV_X1    g0542(.A(G330), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n500), .A2(new_n511), .A3(new_n520), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n605), .A2(new_n544), .A3(KEYINPUT95), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n551), .B2(new_n608), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(G179), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n744), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT95), .B1(new_n605), .B2(new_n544), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n551), .A2(new_n608), .A3(new_n747), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n526), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(KEYINPUT30), .A3(G179), .A4(new_n629), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n608), .A2(G179), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n646), .A2(new_n526), .A3(new_n552), .A4(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT31), .B1(new_n758), .B2(new_n705), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n617), .A2(new_n661), .A3(new_n664), .A4(new_n708), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n743), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n687), .A2(new_n694), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n679), .A2(new_n617), .A3(new_n676), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n705), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT96), .B1(new_n766), .B2(KEYINPUT29), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT96), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n769), .C1(new_n695), .C2(new_n705), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n610), .B(KEYINPUT97), .Z(new_n772));
  NAND3_X1  g0572(.A1(new_n615), .A2(new_n684), .A3(KEYINPUT26), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n691), .A2(KEYINPUT98), .A3(KEYINPUT26), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n693), .A2(KEYINPUT26), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n772), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n661), .A2(new_n533), .A3(new_n616), .ZN(new_n780));
  OAI211_X1 g0580(.A(KEYINPUT29), .B(new_n708), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n763), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n742), .B1(new_n782), .B2(G1), .ZN(G364));
  AOI21_X1  g0583(.A(new_n223), .B1(G20), .B2(new_n393), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n211), .A2(new_n318), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n313), .A2(new_n464), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n464), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n211), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n343), .B1(new_n792), .B2(G77), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n785), .A2(new_n789), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n788), .B(new_n793), .C1(new_n453), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(KEYINPUT32), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(KEYINPUT32), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n211), .B1(new_n796), .B2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n800), .B(new_n801), .C1(G97), .C2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n211), .A2(new_n464), .A3(new_n534), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n806), .A2(G190), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n806), .A2(new_n318), .A3(new_n807), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n804), .B1(new_n202), .B2(new_n808), .C1(new_n428), .C2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n313), .A2(new_n464), .A3(new_n790), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n795), .B(new_n810), .C1(G107), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT33), .B(G317), .Z(new_n815));
  OAI22_X1  g0615(.A1(new_n814), .A2(new_n808), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G311), .A2(new_n792), .B1(new_n798), .B2(G329), .ZN(new_n817));
  INV_X1    g0617(.A(new_n794), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n288), .B1(new_n818), .B2(G322), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(new_n539), .C2(new_n802), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n811), .B1(new_n786), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n816), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n784), .B1(new_n813), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n274), .A2(G20), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n210), .B1(new_n826), .B2(G45), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n736), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n214), .A2(new_n288), .ZN(new_n831));
  INV_X1    g0631(.A(G355), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(G116), .B2(new_n214), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n215), .A2(new_n288), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n222), .B2(new_n490), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n250), .A2(new_n490), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n833), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(G13), .A2(G33), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(G20), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n784), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n830), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n843), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n825), .B(new_n845), .C1(new_n719), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n724), .A2(new_n829), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n719), .A2(G330), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(G396));
  NAND2_X1  g0652(.A1(new_n764), .A2(new_n765), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n396), .A2(new_n708), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n385), .A2(new_n391), .B1(new_n379), .B2(new_n708), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n395), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n394), .B(new_n708), .C1(G179), .C2(new_n384), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n856), .B1(new_n766), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n763), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n829), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n784), .A2(new_n841), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n830), .B1(new_n230), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n808), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n868), .A2(G303), .B1(G116), .B2(new_n792), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n821), .B2(new_n809), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT101), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n794), .A2(new_n539), .B1(new_n802), .B2(new_n205), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT102), .Z(new_n873));
  NAND2_X1  g0673(.A1(new_n812), .A2(G87), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n787), .A2(G107), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n288), .B1(new_n798), .B2(G311), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n818), .B1(new_n792), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n808), .B2(new_n880), .C1(new_n881), .C2(new_n809), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT34), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n812), .A2(G68), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n787), .A2(G50), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n803), .A2(new_n266), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n343), .B1(new_n798), .B2(G132), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n883), .B2(KEYINPUT34), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n871), .A2(new_n878), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n784), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n867), .B1(new_n861), .B2(new_n842), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n865), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(G384));
  XNOR2_X1  g0697(.A(new_n479), .B(KEYINPUT104), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT35), .ZN(new_n899));
  OAI211_X1 g0699(.A(G116), .B(new_n224), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n222), .B(G77), .C1(new_n428), .C2(new_n453), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n202), .A2(G68), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n210), .B(G13), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n366), .A2(new_n705), .ZN(new_n907));
  INV_X1    g0707(.A(new_n359), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n667), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n366), .B(new_n705), .C1(new_n365), .C2(new_n359), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n856), .B2(new_n859), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT16), .B1(new_n455), .B2(new_n446), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n421), .B1(new_n448), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(new_n421), .C1(new_n448), .C2(new_n914), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n471), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n707), .A3(new_n918), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n449), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n470), .A2(new_n471), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n470), .A2(new_n707), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n449), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n920), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n474), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n927), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n913), .A2(new_n934), .B1(new_n666), .B2(new_n703), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  AOI221_X4 g0736(.A(new_n931), .B1(new_n474), .B2(new_n928), .C1(new_n922), .C2(new_n926), .ZN(new_n937));
  INV_X1    g0737(.A(new_n449), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n458), .A2(new_n460), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n466), .B1(new_n939), .B2(new_n421), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n941), .A2(KEYINPUT106), .A3(new_n925), .A4(new_n924), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n926), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n923), .A2(new_n924), .A3(new_n449), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT37), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n474), .A2(new_n470), .A3(new_n707), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n936), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n667), .A2(new_n705), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n935), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n475), .A2(new_n781), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n767), .B2(new_n770), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n673), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n954), .B(new_n957), .Z(new_n958));
  INV_X1    g0758(.A(KEYINPUT107), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n759), .B2(new_n760), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n762), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n860), .B1(new_n909), .B2(new_n910), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n937), .C2(new_n949), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT40), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n758), .A2(new_n705), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT31), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT107), .B1(new_n969), .B2(new_n961), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n762), .A2(new_n962), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n964), .B(new_n966), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n965), .A2(KEYINPUT40), .B1(new_n934), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n475), .A3(new_n963), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n970), .A2(new_n971), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n974), .B1(new_n675), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(G330), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n958), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n210), .B2(new_n826), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n958), .A2(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n906), .B1(new_n981), .B2(new_n982), .ZN(G367));
  NAND2_X1  g0783(.A1(new_n834), .A2(new_n246), .ZN(new_n984));
  INV_X1    g0784(.A(new_n844), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n215), .B2(new_n587), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n830), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n595), .A2(new_n613), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n705), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n615), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n610), .B2(new_n989), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n786), .A2(new_n630), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G311), .A2(new_n868), .B1(new_n992), .B2(KEYINPUT46), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(KEYINPUT46), .B2(new_n992), .C1(new_n539), .C2(new_n809), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G303), .A2(new_n818), .B1(new_n798), .B2(G317), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n995), .B(new_n343), .C1(new_n821), .C2(new_n791), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n811), .A2(new_n205), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n802), .A2(new_n206), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n994), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT109), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1001), .A2(new_n808), .B1(new_n809), .B2(new_n433), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G150), .A2(new_n818), .B1(new_n798), .B2(G137), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n343), .B1(new_n792), .B2(G50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n428), .C2(new_n802), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n230), .A2(new_n811), .B1(new_n786), .B2(new_n453), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT47), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n784), .B1(new_n1008), .B2(KEYINPUT47), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n987), .B1(new_n846), .B2(new_n991), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n705), .A2(new_n489), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n525), .A2(new_n1012), .A3(new_n532), .A4(new_n529), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n684), .A2(new_n705), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n711), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n660), .B1(new_n1018), .B2(new_n586), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n649), .A2(new_n708), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n725), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1015), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(KEYINPUT44), .A3(new_n1022), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n713), .B2(new_n1015), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1016), .A2(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n728), .B2(new_n730), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n723), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT92), .B1(new_n719), .B2(G330), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n727), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n729), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1023), .A2(new_n1016), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n724), .A2(KEYINPUT93), .A3(new_n727), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT108), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n722), .A2(KEYINPUT108), .A3(new_n723), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n726), .A2(new_n1020), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n709), .A2(new_n712), .A3(new_n725), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  MUX2_X1   g0846(.A(new_n1040), .B(new_n1042), .S(new_n1046), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n782), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n736), .B(KEYINPUT41), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n828), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1022), .A2(new_n698), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n708), .B1(new_n1051), .B2(new_n682), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT42), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n727), .A2(new_n1053), .A3(new_n709), .A4(new_n1015), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT42), .B1(new_n1044), .B2(new_n1022), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n728), .A2(new_n730), .A3(new_n1022), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1011), .B1(new_n1050), .B2(new_n1062), .ZN(G387));
  AOI21_X1  g0863(.A(new_n1046), .B1(new_n724), .B2(new_n1039), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n828), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n831), .A2(new_n738), .B1(G107), .B2(new_n214), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n243), .A2(new_n490), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n738), .ZN(new_n1069));
  AOI211_X1 g0869(.A(G45), .B(new_n1069), .C1(G68), .C2(G77), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n375), .A2(new_n202), .ZN(new_n1071));
  XOR2_X1   g0871(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1072));
  XNOR2_X1  g0872(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n835), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1067), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n829), .B1(new_n1075), .B2(new_n985), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT111), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n868), .A2(G159), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT112), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n809), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n267), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n794), .A2(new_n202), .B1(new_n797), .B2(new_n881), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n288), .B1(new_n791), .B2(new_n428), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n802), .A2(new_n374), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n997), .B1(G77), .B2(new_n787), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1079), .A2(new_n1081), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n288), .B1(new_n798), .B2(G326), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G317), .A2(new_n818), .B1(new_n792), .B2(G303), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT113), .B(G322), .Z(new_n1090));
  INV_X1    g0890(.A(G311), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1089), .B1(new_n808), .B2(new_n1090), .C1(new_n1091), .C2(new_n809), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n787), .A2(G294), .B1(G283), .B2(new_n803), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT49), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1088), .B1(new_n630), .B2(new_n811), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1087), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT114), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n784), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1077), .B1(new_n727), .B2(new_n846), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1066), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n782), .A2(new_n1065), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(KEYINPUT115), .A3(new_n736), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n782), .A2(new_n1065), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT115), .B1(new_n1106), .B2(new_n736), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(G393));
  NOR2_X1   g0911(.A1(new_n1015), .A2(new_n846), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT116), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n844), .B1(new_n205), .B2(new_n214), .C1(new_n835), .C2(new_n253), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n829), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n868), .A2(G317), .B1(G311), .B2(new_n818), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT52), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G107), .A2(new_n812), .B1(new_n787), .B2(G283), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n791), .A2(new_n539), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n343), .B1(new_n1090), .B2(new_n797), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(G116), .C2(new_n803), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1121), .C1(new_n822), .C2(new_n809), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n808), .A2(new_n881), .B1(new_n433), .B2(new_n794), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT51), .Z(new_n1124));
  OAI221_X1 g0924(.A(new_n288), .B1(new_n797), .B2(new_n1001), .C1(new_n376), .C2(new_n791), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G77), .B2(new_n803), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G68), .A2(new_n787), .B1(new_n812), .B2(G87), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n202), .C2(new_n809), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1117), .A2(new_n1122), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1115), .B1(new_n1129), .B2(new_n784), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1113), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1038), .B2(new_n827), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n771), .A2(new_n781), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1133), .A2(new_n863), .A3(new_n1065), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1038), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n737), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1106), .A2(new_n1038), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1132), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G390));
  INV_X1    g0939(.A(new_n952), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n937), .B2(new_n949), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n708), .B(new_n858), .C1(new_n779), .C2(new_n780), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n912), .B1(new_n1142), .B2(new_n859), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n763), .A2(new_n861), .A3(new_n911), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n950), .A2(new_n951), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n856), .A2(new_n859), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n952), .B1(new_n1147), .B2(new_n911), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1144), .B(new_n1145), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n963), .A2(G330), .A3(new_n964), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n854), .B1(new_n764), .B2(new_n765), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n859), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n911), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n950), .A2(new_n951), .B1(new_n1154), .B2(new_n1140), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n827), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1146), .A2(new_n842), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n786), .A2(new_n881), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n808), .C1(new_n880), .C2(new_n809), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n791), .A2(new_n1165), .B1(new_n797), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n343), .B(new_n1167), .C1(G132), .C2(new_n818), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n202), .B2(new_n811), .C1(new_n433), .C2(new_n802), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n885), .B1(new_n539), .B2(new_n797), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT119), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G107), .A2(new_n1080), .B1(new_n868), .B2(G283), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n803), .A2(G77), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n343), .B1(new_n794), .B2(new_n630), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G97), .B2(new_n792), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n788), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1164), .A2(new_n1169), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1177), .A2(new_n784), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n830), .B(new_n1178), .C1(new_n268), .C2(new_n866), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1159), .B1(new_n1160), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(KEYINPUT118), .B(G330), .C1(new_n970), .C2(new_n971), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n861), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT118), .B1(new_n963), .B2(G330), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n912), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1145), .A2(new_n859), .A3(new_n1142), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n762), .A2(new_n962), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n743), .B1(new_n1187), .B2(new_n960), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n969), .A2(new_n961), .ZN(new_n1189));
  AND4_X1   g0989(.A1(new_n617), .A2(new_n661), .A3(new_n664), .A4(new_n708), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G330), .B(new_n861), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1188), .A2(new_n964), .B1(new_n1191), .B2(new_n912), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT117), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n912), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1150), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT117), .B1(new_n1197), .B2(new_n1147), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1186), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1188), .A2(new_n475), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n956), .A2(new_n673), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1158), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1199), .A2(new_n1149), .A3(new_n1157), .A4(new_n1202), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n736), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1180), .A2(new_n1206), .ZN(G378));
  AOI21_X1  g1007(.A(new_n830), .B1(new_n202), .B2(new_n866), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G128), .A2(new_n818), .B1(new_n792), .B2(G137), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n881), .B2(new_n802), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1165), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n787), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1080), .A2(G132), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n1166), .C2(new_n808), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n812), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G97), .A2(new_n1080), .B1(new_n868), .B2(G116), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n787), .A2(G77), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n732), .B(new_n343), .C1(new_n791), .C2(new_n374), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n794), .A2(new_n206), .B1(new_n797), .B2(new_n821), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G68), .C2(new_n803), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n812), .A2(new_n266), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT58), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G50), .B1(new_n255), .B2(new_n732), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n288), .B2(G41), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT120), .Z(new_n1232));
  AND4_X1   g1032(.A1(new_n1219), .A2(new_n1228), .A3(new_n1229), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n280), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(new_n703), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n322), .A2(new_n370), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n322), .B2(new_n370), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1208), .B1(new_n1103), .B2(new_n1233), .C1(new_n1244), .C2(new_n842), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT121), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1245), .B(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT122), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n974), .B2(new_n743), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n947), .A2(new_n948), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n931), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n933), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n963), .A2(new_n964), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n966), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n972), .B1(new_n933), .B2(new_n932), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT122), .B(G330), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1249), .A2(new_n1256), .A3(new_n1244), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n975), .A2(KEYINPUT122), .A3(G330), .A4(new_n1243), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n954), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n913), .A2(new_n934), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n666), .A2(new_n703), .ZN(new_n1263));
  AND4_X1   g1063(.A1(KEYINPUT123), .A2(new_n953), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT123), .B1(new_n935), .B2(new_n953), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1261), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1247), .B1(new_n1268), .B2(new_n828), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1205), .A2(new_n1202), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT57), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1205), .B2(new_n1202), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1257), .A2(new_n954), .A3(new_n1258), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n954), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n736), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1269), .B1(new_n1271), .B2(new_n1277), .ZN(G375));
  OAI21_X1  g1078(.A(KEYINPUT124), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1193), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1197), .A2(KEYINPUT117), .A3(new_n1147), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1280), .A2(new_n1281), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n957), .A2(new_n1200), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1279), .A2(new_n1285), .A3(new_n1049), .A4(new_n1203), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n912), .A2(new_n841), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(G107), .A2(new_n792), .B1(new_n798), .B2(G303), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1288), .B(new_n343), .C1(new_n821), .C2(new_n794), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n230), .A2(new_n811), .B1(new_n786), .B2(new_n205), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1084), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n630), .B2(new_n809), .C1(new_n539), .C2(new_n808), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(G132), .A2(new_n868), .B1(new_n1080), .B2(new_n1211), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n288), .B1(new_n794), .B2(new_n880), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n791), .A2(new_n881), .B1(new_n797), .B2(new_n1163), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1294), .B(new_n1295), .C1(G50), .C2(new_n803), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n787), .A2(G159), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1293), .A2(new_n1225), .A3(new_n1296), .A4(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1103), .B1(new_n1292), .B2(new_n1298), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n830), .B(new_n1299), .C1(new_n428), .C2(new_n866), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1282), .B2(new_n827), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1286), .A2(new_n1303), .ZN(G381));
  AND3_X1   g1104(.A1(new_n1266), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n828), .B1(new_n1305), .B2(new_n1275), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1247), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1270), .B1(new_n1305), .B2(new_n1275), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1272), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1257), .A2(new_n1258), .A3(new_n954), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1261), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n737), .B1(new_n1312), .B2(new_n1273), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1308), .B1(new_n1310), .B2(new_n1313), .ZN(new_n1314));
  NOR4_X1   g1114(.A1(G378), .A2(G381), .A3(G384), .A4(G390), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT115), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1134), .B2(new_n737), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1108), .A3(new_n1107), .ZN(new_n1318));
  INV_X1    g1118(.A(G396), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1105), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1320), .A2(G387), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1314), .A2(new_n1315), .A3(new_n1321), .ZN(G407));
  INV_X1    g1122(.A(G378), .ZN(new_n1323));
  INV_X1    g1123(.A(G213), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(G343), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1314), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G407), .A2(new_n1326), .A3(G213), .ZN(G409));
  OAI211_X1 g1127(.A(G378), .B(new_n1269), .C1(new_n1271), .C2(new_n1277), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1049), .B(new_n1270), .C1(new_n1305), .C2(new_n1275), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n828), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1307), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1323), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1328), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1325), .ZN(new_n1334));
  OAI21_X1  g1134(.A(KEYINPUT60), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1279), .A3(new_n1285), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n737), .B1(new_n1337), .B2(KEYINPUT60), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(G384), .B1(new_n1339), .B2(new_n1303), .ZN(new_n1340));
  AOI211_X1 g1140(.A(new_n896), .B(new_n1302), .C1(new_n1336), .C2(new_n1338), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1333), .A2(new_n1334), .A3(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT125), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1346), .B1(G387), .B2(new_n1138), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(G393), .A2(G396), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1319), .B1(new_n1318), .B2(new_n1105), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1347), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(G387), .B(new_n1138), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G393), .A2(G396), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1320), .ZN(new_n1354));
  OR2_X1    g1154(.A1(G387), .A2(new_n1138), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G387), .A2(new_n1138), .ZN(new_n1356));
  AOI22_X1  g1156(.A1(new_n1354), .A2(new_n1347), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1352), .A2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1325), .B1(new_n1328), .B2(new_n1332), .ZN(new_n1359));
  NOR3_X1   g1159(.A1(new_n1340), .A2(new_n1341), .A3(new_n1344), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1358), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1325), .A2(G2897), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1340), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1341), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1362), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1362), .ZN(new_n1366));
  NOR3_X1   g1166(.A1(new_n1340), .A2(new_n1341), .A3(new_n1366), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1365), .A2(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1247), .B1(new_n1312), .B2(new_n828), .ZN(new_n1369));
  AOI21_X1  g1169(.A(G378), .B1(new_n1369), .B2(new_n1329), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1370), .B1(new_n1314), .B2(G378), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1368), .B1(new_n1371), .B2(new_n1325), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT61), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1345), .A2(new_n1361), .A3(new_n1372), .A4(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(KEYINPUT126), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1342), .A2(new_n1362), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1366), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1373), .B1(new_n1359), .B2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT126), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1380), .A2(new_n1381), .A3(new_n1345), .A4(new_n1361), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1375), .A2(new_n1382), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1379), .A2(KEYINPUT127), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT127), .ZN(new_n1385));
  OAI211_X1 g1185(.A(new_n1385), .B(new_n1373), .C1(new_n1359), .C2(new_n1378), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1343), .A2(KEYINPUT62), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT62), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1359), .A2(new_n1388), .A3(new_n1342), .ZN(new_n1389));
  NAND4_X1  g1189(.A1(new_n1384), .A2(new_n1386), .A3(new_n1387), .A4(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1390), .A2(new_n1358), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1383), .A2(new_n1391), .ZN(G405));
  NOR2_X1   g1192(.A1(new_n1314), .A2(G378), .ZN(new_n1393));
  INV_X1    g1193(.A(new_n1328), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  INV_X1    g1195(.A(new_n1342), .ZN(new_n1396));
  XNOR2_X1  g1196(.A(new_n1395), .B(new_n1396), .ZN(new_n1397));
  XNOR2_X1  g1197(.A(new_n1397), .B(new_n1358), .ZN(G402));
endmodule


