//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  XOR2_X1   g000(.A(KEYINPUT26), .B(G101), .Z(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G134), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT11), .B1(new_n199), .B2(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n197), .A2(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n206), .A3(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(G128), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT64), .A3(G146), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT64), .B1(new_n209), .B2(G146), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n213), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n209), .A2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n213), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT68), .A3(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n201), .A2(KEYINPUT67), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n199), .B2(G137), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(G131), .C1(new_n201), .C2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n208), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT0), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n222), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n224), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n244), .B2(new_n213), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n222), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n200), .A2(new_n201), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT66), .A3(G131), .A4(new_n198), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n202), .B2(new_n203), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n205), .A2(new_n207), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n236), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G119), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G116), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT2), .B(G113), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n250), .A2(new_n252), .ZN(new_n265));
  INV_X1    g079(.A(new_n207), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n206), .B1(new_n202), .B2(new_n203), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n247), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n263), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n236), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n195), .B1(new_n264), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n195), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n194), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n254), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n269), .A2(KEYINPUT30), .A3(new_n236), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n263), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n271), .A3(new_n192), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT31), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n279), .A2(new_n282), .A3(new_n271), .A4(new_n192), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n194), .C1(new_n272), .C2(new_n273), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n275), .A2(new_n281), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(KEYINPUT73), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT32), .B1(new_n286), .B2(new_n289), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n254), .A2(new_n263), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n270), .B1(new_n269), .B2(new_n236), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT28), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n271), .A2(new_n195), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n192), .B(KEYINPUT71), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT74), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n279), .A2(new_n271), .ZN(new_n301));
  INV_X1    g115(.A(new_n192), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n296), .A2(new_n305), .A3(new_n297), .A4(new_n298), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n300), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n272), .A2(new_n273), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n302), .A2(new_n304), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n293), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n291), .A2(new_n292), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G953), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G221), .A3(G234), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT22), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(G137), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n255), .B2(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n222), .A2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G110), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n255), .A2(G128), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n321), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n222), .A2(G119), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n255), .A2(G128), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n326), .A2(new_n322), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n330), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n318), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n326), .A2(new_n322), .A3(new_n334), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n326), .B2(new_n322), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n329), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT79), .A3(new_n327), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n212), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  INV_X1    g160(.A(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G140), .ZN(new_n348));
  AND4_X1   g162(.A1(new_n342), .A2(new_n346), .A3(new_n348), .A4(new_n212), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT78), .B1(new_n346), .B2(KEYINPUT16), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT16), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n345), .A4(G125), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n351), .A2(G146), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n337), .A2(new_n341), .A3(new_n350), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT81), .ZN(new_n358));
  INV_X1    g172(.A(new_n356), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n340), .A2(new_n327), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(new_n318), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n341), .A4(new_n350), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n212), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n356), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n321), .A2(new_n326), .A3(new_n324), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G110), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n333), .A2(new_n330), .A3(new_n335), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT82), .B1(new_n364), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n374), .B(new_n371), .C1(new_n358), .C2(new_n363), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n317), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G902), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n364), .A2(new_n372), .A3(new_n316), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT25), .ZN(new_n380));
  INV_X1    g194(.A(G234), .ZN(new_n381));
  OAI21_X1  g195(.A(G217), .B1(new_n381), .B2(G902), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n382), .B(KEYINPUT75), .Z(new_n383));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n376), .A2(new_n384), .A3(new_n377), .A4(new_n378), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n380), .A2(KEYINPUT83), .A3(new_n383), .A4(new_n385), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n383), .A2(G902), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n378), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n312), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT68), .B1(new_n228), .B2(new_n223), .ZN(new_n396));
  AND4_X1   g210(.A1(KEYINPUT68), .A2(new_n223), .A3(new_n213), .A4(new_n224), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n210), .A2(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n237), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT85), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G104), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G107), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n403), .A2(G107), .ZN(new_n406));
  OAI21_X1  g220(.A(G101), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n403), .B2(G107), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n409));
  INV_X1    g223(.A(G107), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G104), .ZN(new_n411));
  INV_X1    g225(.A(G101), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n408), .A2(new_n411), .A3(new_n412), .A4(new_n404), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n402), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n221), .A2(new_n230), .A3(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n253), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT12), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT12), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n421), .B(new_n253), .C1(new_n416), .C2(new_n417), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n394), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(G110), .B(G140), .Z(new_n424));
  AND2_X1   g238(.A1(new_n313), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT10), .B1(new_n402), .B2(new_n415), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n408), .A2(new_n411), .A3(new_n404), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(G101), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(G101), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n413), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n247), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n231), .A2(KEYINPUT10), .A3(new_n415), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n428), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n427), .B1(new_n436), .B2(new_n253), .ZN(new_n437));
  INV_X1    g251(.A(new_n417), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n415), .B2(new_n402), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n421), .B1(new_n439), .B2(new_n253), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n418), .A2(KEYINPUT12), .A3(new_n419), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT86), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n423), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT87), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n436), .A2(new_n253), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n436), .A2(new_n253), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n427), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n423), .A2(new_n437), .A3(new_n442), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n377), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n377), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n446), .B1(new_n422), .B2(new_n420), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n427), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n445), .A2(new_n437), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G469), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT9), .B(G234), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT84), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n231), .A2(new_n347), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n248), .B2(new_n347), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n313), .A2(G224), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(G110), .B(G122), .Z(new_n472));
  NAND3_X1  g286(.A1(new_n433), .A2(new_n263), .A3(new_n431), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(G113), .C1(KEYINPUT5), .C2(new_n256), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n415), .A2(new_n261), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT89), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT89), .B1(new_n473), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n472), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n471), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n469), .A2(new_n470), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n414), .A2(KEYINPUT90), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n475), .A2(new_n261), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n487), .B(new_n488), .Z(new_n489));
  XOR2_X1   g303(.A(new_n472), .B(KEYINPUT8), .Z(new_n490));
  AOI21_X1  g304(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n469), .A2(KEYINPUT7), .A3(new_n470), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n483), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n494), .A3(new_n377), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n485), .A2(new_n494), .A3(new_n377), .A4(new_n496), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT91), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT88), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n495), .A2(new_n503), .A3(new_n497), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n313), .A2(G952), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(G237), .ZN(new_n506));
  NAND2_X1  g320(.A1(G234), .A2(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G902), .A3(G953), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n508), .B(KEYINPUT98), .Z(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT21), .B(G898), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n500), .A2(new_n502), .A3(new_n504), .A4(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n467), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G113), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(new_n403), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n188), .A2(G214), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(G143), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n209), .A2(KEYINPUT92), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n520), .A2(new_n521), .A3(G214), .A4(new_n188), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n203), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n522), .A3(G131), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n519), .A2(new_n522), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT17), .A3(G131), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(new_n356), .A3(new_n366), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n346), .A2(new_n348), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G146), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n344), .B2(new_n349), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT93), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(KEYINPUT18), .A3(G131), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(new_n532), .C1(new_n344), .C2(new_n349), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n523), .B1(new_n538), .B2(new_n203), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n535), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n516), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT95), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n530), .A2(new_n540), .A3(new_n516), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n542), .B(new_n377), .C1(new_n545), .C2(new_n541), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G475), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n524), .A2(new_n526), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n343), .B(KEYINPUT19), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n212), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n356), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n540), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n516), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n540), .A2(KEYINPUT94), .A3(new_n552), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G475), .B1(new_n558), .B2(new_n543), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n548), .B1(new_n559), .B2(new_n377), .ZN(new_n560));
  INV_X1    g374(.A(new_n543), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n516), .B1(new_n553), .B2(new_n554), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n557), .ZN(new_n563));
  NOR4_X1   g377(.A1(new_n563), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n547), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n222), .A2(G143), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT97), .ZN(new_n567));
  OAI21_X1  g381(.A(G134), .B1(new_n567), .B2(KEYINPUT13), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n566), .B(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n222), .B2(G143), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n568), .A2(new_n571), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n574));
  INV_X1    g388(.A(G122), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(G116), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n257), .A2(KEYINPUT96), .A3(G122), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n576), .A2(new_n577), .B1(G116), .B2(new_n575), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G107), .ZN(new_n579));
  INV_X1    g393(.A(new_n578), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n410), .ZN(new_n581));
  OAI22_X1  g395(.A1(new_n572), .A2(new_n573), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n571), .A2(new_n199), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT14), .B1(new_n576), .B2(new_n577), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n580), .B1(KEYINPUT14), .B2(new_n410), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n571), .A2(new_n199), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n462), .A2(G217), .A3(new_n313), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n582), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n582), .B2(new_n588), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n377), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n565), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n393), .A2(new_n514), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  NAND2_X1  g416(.A1(new_n286), .A2(new_n377), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n286), .A2(new_n289), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n392), .A2(new_n467), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n501), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n498), .B2(new_n499), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n512), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n594), .A2(new_n595), .ZN(new_n611));
  INV_X1    g425(.A(new_n593), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n592), .B2(new_n593), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n377), .A2(G478), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n565), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n607), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT99), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT34), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G104), .ZN(G6));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n560), .B2(new_n564), .ZN(new_n626));
  INV_X1    g440(.A(G475), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n540), .A2(KEYINPUT94), .A3(new_n552), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT94), .B1(new_n540), .B2(new_n552), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n629), .A3(new_n516), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n627), .B(new_n377), .C1(new_n630), .C2(new_n561), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT20), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n559), .A2(new_n548), .A3(new_n377), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(KEYINPUT100), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n597), .A2(new_n598), .B1(G475), .B2(new_n546), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n610), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n607), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  INV_X1    g456(.A(new_n606), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n514), .A2(new_n600), .A3(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n373), .A2(new_n375), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n317), .A2(KEYINPUT36), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT101), .Z(new_n647));
  OR2_X1    g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n390), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n388), .A2(new_n389), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT37), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G110), .ZN(G12));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n506), .B1(new_n509), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n632), .A2(KEYINPUT100), .A3(new_n633), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT100), .B1(new_n632), .B2(new_n633), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n637), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n635), .A2(KEYINPUT102), .A3(new_n637), .A4(new_n658), .ZN(new_n664));
  AND4_X1   g478(.A1(new_n466), .A2(new_n663), .A3(new_n461), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n307), .A2(new_n310), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT32), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n605), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n669), .A3(new_n290), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n651), .A2(new_n670), .A3(new_n609), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  INV_X1    g487(.A(new_n467), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n657), .B(KEYINPUT39), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n674), .A2(KEYINPUT40), .A3(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n632), .A2(new_n633), .B1(G475), .B2(new_n546), .ZN(new_n682));
  INV_X1    g496(.A(new_n599), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n651), .A2(new_n608), .A3(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT103), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n264), .A2(new_n271), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n280), .B1(new_n689), .B2(new_n298), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n293), .B1(new_n690), .B2(new_n377), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n291), .A2(new_n292), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n686), .B2(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n500), .A2(new_n504), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n681), .A2(new_n687), .A3(new_n693), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  NAND3_X1  g512(.A1(new_n565), .A2(new_n618), .A3(new_n658), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n565), .A2(new_n701), .A3(new_n618), .A4(new_n658), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n466), .A2(new_n700), .A3(new_n461), .A4(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n670), .A3(new_n609), .A4(new_n651), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  NAND2_X1  g519(.A1(new_n451), .A2(new_n377), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(KEYINPUT105), .A3(G469), .ZN(new_n707));
  NAND2_X1  g521(.A1(KEYINPUT105), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n451), .A2(new_n377), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n707), .A2(new_n466), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n393), .A2(new_n620), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND3_X1  g527(.A1(new_n393), .A2(new_n639), .A3(new_n710), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AND4_X1   g529(.A1(new_n466), .A2(new_n707), .A3(new_n609), .A4(new_n709), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n512), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n651), .A2(new_n670), .A3(new_n600), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n255), .ZN(G21));
  NAND2_X1  g534(.A1(new_n684), .A2(new_n609), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n511), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n274), .A2(new_n283), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n288), .B1(new_n723), .B2(new_n281), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT106), .B(G472), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n724), .B1(new_n603), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n388), .A3(new_n389), .A4(new_n391), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n710), .B(new_n722), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n710), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n726), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT108), .B1(new_n738), .B2(new_n722), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT109), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n575), .ZN(G24));
  NAND2_X1  g556(.A1(new_n700), .A2(new_n702), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n716), .A2(new_n744), .A3(new_n651), .A4(new_n726), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n694), .A2(new_n501), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n734), .A3(new_n670), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n744), .A2(new_n674), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n393), .A2(new_n703), .A3(KEYINPUT42), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  INV_X1    g569(.A(new_n750), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n665), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND2_X1  g572(.A1(new_n682), .A2(new_n618), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT112), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n682), .A2(KEYINPUT43), .A3(new_n618), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n759), .A2(new_n764), .A3(new_n760), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n643), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT113), .A4(new_n765), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n651), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n453), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n459), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n457), .A2(KEYINPUT45), .A3(new_n458), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n459), .A2(KEYINPUT45), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(G469), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n455), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n773), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n452), .B1(new_n774), .B2(new_n777), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n454), .B1(new_n784), .B2(new_n779), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n465), .B(new_n675), .C1(new_n783), .C2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n768), .A2(KEYINPUT44), .A3(new_n651), .A4(new_n769), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n772), .A2(new_n749), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  INV_X1    g604(.A(new_n786), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n453), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n466), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT47), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n734), .A2(new_n670), .A3(new_n743), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n796), .B(new_n466), .C1(new_n791), .C2(new_n792), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n749), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NOR2_X1   g613(.A1(new_n651), .A2(new_n657), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n291), .A2(new_n292), .ZN(new_n801));
  INV_X1    g615(.A(new_n691), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n721), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n803), .A3(new_n674), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n672), .A2(new_n704), .A3(new_n745), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n651), .A2(new_n726), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n743), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n810), .A2(new_n716), .B1(new_n665), .B2(new_n671), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n704), .A4(new_n804), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n805), .A2(new_n814), .A3(new_n806), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n711), .B(new_n714), .C1(new_n717), .C2(new_n718), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n732), .B2(new_n739), .ZN(new_n820));
  INV_X1    g634(.A(new_n644), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n637), .B1(new_n560), .B2(new_n564), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n513), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n821), .A2(new_n651), .B1(new_n607), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n392), .A2(new_n467), .ZN(new_n825));
  INV_X1    g639(.A(new_n513), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n619), .B(KEYINPUT114), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n643), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n828), .A2(new_n601), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n828), .B2(new_n601), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n674), .A2(new_n683), .A3(new_n547), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n748), .A2(new_n636), .A3(new_n657), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n670), .A3(new_n651), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n703), .A2(new_n651), .A3(new_n726), .A4(new_n749), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n754), .A2(new_n757), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n820), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n817), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n607), .A2(new_n823), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n652), .B2(new_n644), .ZN(new_n842));
  INV_X1    g656(.A(new_n831), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n828), .A2(new_n601), .A3(new_n829), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n754), .A2(new_n757), .A3(new_n835), .A4(new_n836), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n812), .A2(new_n807), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n730), .A2(new_n731), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n722), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n818), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n840), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n814), .B1(new_n805), .B2(new_n806), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n805), .A2(new_n806), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n815), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n846), .A2(new_n845), .A3(new_n850), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT53), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n838), .A2(new_n839), .A3(new_n847), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT54), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT117), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n733), .A2(new_n748), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n734), .A3(new_n506), .A4(new_n692), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(new_n619), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n853), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n865), .A2(new_n565), .A3(new_n618), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n794), .A2(new_n797), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n707), .A2(new_n709), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n465), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n748), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n766), .A2(new_n506), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n729), .B2(new_n728), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n869), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n864), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n809), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT119), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n738), .A2(new_n608), .A3(new_n695), .A4(new_n874), .ZN(new_n881));
  NOR2_X1   g695(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n877), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n877), .A2(KEYINPUT51), .A3(new_n880), .A4(new_n883), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n734), .A2(new_n670), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT48), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n505), .B(new_n890), .C1(new_n716), .C2(new_n876), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n863), .A2(new_n866), .A3(new_n868), .A4(new_n892), .ZN(new_n893));
  OR2_X1    g707(.A1(G952), .A2(G953), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n502), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n696), .A2(new_n465), .A3(new_n896), .A4(new_n759), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n871), .B(KEYINPUT49), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n734), .A3(new_n692), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(G75));
  XOR2_X1   g714(.A(new_n471), .B(KEYINPUT55), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n860), .A2(new_n861), .A3(G210), .A4(G902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n481), .A2(new_n484), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT120), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  INV_X1    g725(.A(new_n906), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n901), .A3(new_n907), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n313), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(G51));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n839), .B1(new_n817), .B2(new_n838), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n860), .A2(KEYINPUT54), .A3(new_n861), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n454), .B(KEYINPUT57), .Z(new_n924));
  OAI21_X1  g738(.A(new_n451), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n919), .A2(new_n920), .A3(new_n377), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n779), .A3(new_n784), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n915), .B1(new_n925), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n563), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT58), .A4(G902), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n563), .B1(new_n931), .B2(new_n627), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n932), .A3(new_n916), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n930), .A2(new_n932), .A3(KEYINPUT121), .A4(new_n916), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G60));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  AOI211_X1 g753(.A(new_n616), .B(new_n939), .C1(new_n921), .C2(new_n922), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n867), .B1(new_n921), .B2(new_n853), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n853), .A2(new_n867), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n915), .B(new_n940), .C1(new_n944), .C2(new_n616), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n860), .A2(new_n861), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n376), .A2(new_n378), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n915), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT61), .B1(new_n951), .B2(KEYINPUT122), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n919), .A2(new_n920), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(new_n648), .A3(new_n649), .A4(new_n948), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n952), .B(new_n955), .ZN(G66));
  INV_X1    g770(.A(G224), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n510), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n820), .A2(new_n832), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n906), .B1(G898), .B2(new_n313), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  AOI21_X1  g776(.A(new_n313), .B1(G227), .B2(G900), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  INV_X1    g778(.A(new_n963), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n789), .A2(new_n798), .ZN(new_n968));
  INV_X1    g782(.A(new_n677), .ZN(new_n969));
  INV_X1    g783(.A(new_n822), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n756), .B(new_n969), .C1(new_n970), .C2(new_n827), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n672), .A2(new_n704), .A3(new_n745), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT62), .B1(new_n697), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n697), .A2(new_n972), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n968), .B(new_n971), .C1(new_n973), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n277), .A2(new_n278), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n550), .B(KEYINPUT123), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n974), .B(new_n975), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(new_n984), .A3(new_n968), .A4(new_n971), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n978), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n793), .A2(new_n888), .A3(new_n675), .A4(new_n721), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT126), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n798), .A2(new_n754), .A3(new_n757), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n789), .A2(KEYINPUT125), .A3(new_n972), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT125), .B1(new_n789), .B2(new_n972), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n981), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n986), .A2(new_n313), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n981), .A2(G900), .A3(G953), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n964), .B(new_n967), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  AND4_X1   g810(.A1(new_n966), .A2(new_n994), .A3(new_n965), .A4(new_n995), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n992), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n959), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1003), .A2(new_n301), .A3(new_n192), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n301), .A2(new_n192), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n978), .A2(new_n959), .A3(new_n985), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n840), .A2(new_n852), .A3(new_n1005), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n301), .A2(new_n192), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1008), .A2(new_n1009), .A3(new_n1001), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n1004), .A2(new_n1007), .A3(new_n915), .A4(new_n1010), .ZN(G57));
endmodule


