//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT68), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT70), .Z(new_n462));
  NOR2_X1   g037(.A1(new_n460), .A2(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n468), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(new_n473), .ZN(G160));
  NAND3_X1  g049(.A1(new_n466), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(new_n465), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n468), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT72), .Z(new_n482));
  INV_X1    g057(.A(G2104), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n477), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n482), .A2(new_n485), .B1(new_n486), .B2(G136), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n477), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n468), .C1(new_n464), .C2(new_n465), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(new_n468), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n477), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI211_X1 g083(.A(G50), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT74), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT73), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n515), .B2(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n513), .A2(new_n514), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n505), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT6), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n508), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n510), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  OAI211_X1 g106(.A(G51), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT7), .Z(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n527), .B2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  OAI21_X1  g116(.A(new_n526), .B1(new_n511), .B2(new_n502), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(G52), .A3(G543), .ZN(new_n543));
  OAI211_X1 g118(.A(G90), .B(new_n515), .C1(new_n507), .C2(new_n508), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n513), .B2(new_n514), .ZN(new_n546));
  AND2_X1   g121(.A1(G77), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n512), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n543), .A2(new_n544), .A3(new_n548), .ZN(G171));
  OAI211_X1 g124(.A(G43), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n550));
  OAI211_X1 g125(.A(G81), .B(new_n515), .C1(new_n507), .C2(new_n508), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n513), .B2(new_n514), .ZN(new_n553));
  AND2_X1   g128(.A1(G68), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n512), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT77), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n550), .A2(new_n551), .A3(new_n558), .A4(new_n555), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND3_X1  g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n542), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g147(.A(G91), .B(new_n515), .C1(new_n507), .C2(new_n508), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n513), .B2(new_n514), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(KEYINPUT78), .A2(G78), .A3(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n572), .A2(new_n583), .ZN(G299));
  NAND3_X1  g159(.A1(new_n543), .A2(new_n544), .A3(new_n548), .ZN(G301));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND2_X1  g161(.A1(G166), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n520), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(new_n517), .A3(new_n518), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(new_n512), .B1(G88), .B2(new_n527), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n509), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n587), .A2(new_n594), .ZN(G303));
  OAI211_X1 g170(.A(G49), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n515), .B1(new_n507), .B2(new_n508), .ZN(new_n598));
  INV_X1    g173(.A(G87), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(new_n527), .A2(G86), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n542), .A2(G48), .A3(G543), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n515), .A2(G61), .ZN(new_n603));
  AND2_X1   g178(.A1(G73), .A2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n512), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(G305));
  OAI211_X1 g181(.A(G47), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n513), .B2(new_n514), .ZN(new_n609));
  AND2_X1   g184(.A1(G72), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n512), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n607), .B(new_n611), .C1(new_n598), .C2(new_n612), .ZN(G290));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(G301), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g190(.A(G54), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n513), .B2(new_n514), .ZN(new_n618));
  AND2_X1   g193(.A1(G79), .A2(G543), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n542), .A2(new_n623), .A3(G92), .A4(new_n515), .ZN(new_n624));
  OAI211_X1 g199(.A(G92), .B(new_n515), .C1(new_n507), .C2(new_n508), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n622), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n621), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n615), .B1(new_n627), .B2(new_n614), .ZN(G321));
  XNOR2_X1  g203(.A(G321), .B(KEYINPUT81), .ZN(G284));
  MUX2_X1   g204(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g205(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n627), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n557), .A2(new_n559), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n626), .A2(new_n624), .ZN(new_n636));
  INV_X1    g211(.A(new_n621), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n638), .A2(G559), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n635), .B1(G868), .B2(new_n639), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n486), .A2(G2104), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n486), .A2(G135), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT82), .ZN(new_n647));
  MUX2_X1   g222(.A(G99), .B(G111), .S(G2105), .Z(new_n648));
  AOI22_X1  g223(.A1(new_n479), .A2(G123), .B1(G2104), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(G156));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  INV_X1    g230(.A(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2427), .ZN(new_n658));
  INV_X1    g233(.A(G2430), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT17), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n672), .A3(new_n674), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n674), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n672), .A2(new_n674), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(new_n676), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n679), .A2(new_n651), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n651), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G2100), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n686), .B2(new_n687), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1956), .B(G2474), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1961), .B(G1966), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(KEYINPUT85), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT19), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n693), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(new_n697), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n701), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G1991), .B(G1996), .Z(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n711), .B(new_n714), .ZN(G229));
  NOR2_X1   g290(.A1(G16), .A2(G23), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT87), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(G288), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT33), .B(G1976), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(G166), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G16), .B2(G22), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G6), .A2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G305), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT32), .B(G1981), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n725), .B(new_n730), .C1(new_n724), .C2(new_n723), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT34), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(G25), .A2(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n479), .A2(G119), .ZN(new_n738));
  MUX2_X1   g313(.A(G95), .B(G107), .S(G2105), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G2104), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n486), .A2(G131), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n737), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n744));
  XOR2_X1   g319(.A(new_n743), .B(new_n744), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n718), .A2(G24), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT86), .Z(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G290), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G1986), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n745), .A2(KEYINPUT89), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n735), .A2(new_n736), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G171), .A2(new_n718), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G5), .B2(new_n718), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G160), .A2(G29), .ZN(new_n760));
  NOR2_X1   g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n760), .A2(G2084), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT31), .B(G11), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT30), .B(G28), .Z(new_n768));
  OAI211_X1 g343(.A(new_n766), .B(new_n767), .C1(G29), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(G2084), .B1(new_n760), .B2(new_n765), .ZN(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n650), .A2(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n759), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n479), .A2(G129), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT26), .Z(new_n776));
  NAND3_X1  g351(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n777));
  INV_X1    g352(.A(G141), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n776), .B(new_n777), .C1(new_n471), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n771), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n771), .B2(G32), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n771), .A2(G27), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n500), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT97), .B(G2078), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n771), .A2(G26), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT28), .Z(new_n794));
  MUX2_X1   g369(.A(G104), .B(G116), .S(G2105), .Z(new_n795));
  AOI22_X1  g370(.A1(new_n486), .A2(G140), .B1(G2104), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n479), .ZN(new_n797));
  INV_X1    g372(.A(G128), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n794), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(G2067), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n758), .B2(new_n757), .ZN(new_n803));
  NOR2_X1   g378(.A1(G29), .A2(G33), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT91), .Z(new_n805));
  AOI22_X1  g380(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n468), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT25), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n486), .A2(G139), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n805), .B1(new_n815), .B2(new_n771), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2072), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n773), .A2(new_n792), .A3(new_n803), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n771), .A2(G35), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT98), .Z(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G162), .B2(new_n771), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G2090), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n627), .A2(G16), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G4), .B2(G16), .ZN(new_n827));
  INV_X1    g402(.A(G1348), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n827), .A2(new_n828), .ZN(new_n832));
  NOR4_X1   g407(.A1(new_n818), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n718), .A2(G19), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n560), .B2(new_n718), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT90), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1341), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n782), .A2(new_n785), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT94), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n718), .A2(G21), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G168), .B2(new_n718), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT95), .B(G1966), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n841), .B(new_n842), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n718), .A2(G20), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT23), .Z(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G299), .B2(G16), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT100), .B(G1956), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n839), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n833), .A2(new_n837), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n753), .B2(new_n754), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n755), .A2(new_n851), .ZN(G311));
  OR2_X1    g427(.A1(new_n755), .A2(new_n851), .ZN(G150));
  NAND2_X1  g428(.A1(new_n627), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n511), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(G55), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n859));
  OAI211_X1 g434(.A(G93), .B(new_n515), .C1(new_n507), .C2(new_n508), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n556), .B(new_n858), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n864), .B1(new_n868), .B2(new_n634), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n855), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n872));
  AOI21_X1  g447(.A(G860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(G145));
  XNOR2_X1  g453(.A(new_n650), .B(new_n488), .ZN(new_n879));
  XOR2_X1   g454(.A(G160), .B(KEYINPUT102), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G142), .ZN(new_n882));
  AND2_X1   g457(.A1(G118), .A2(G2105), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(G106), .B2(new_n468), .ZN(new_n884));
  OAI22_X1  g459(.A1(new_n471), .A2(new_n882), .B1(new_n483), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G130), .B2(new_n479), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n643), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n643), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n888), .B(new_n889), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n742), .A2(KEYINPUT103), .ZN(new_n896));
  INV_X1    g471(.A(new_n889), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n896), .B(new_n892), .C1(new_n897), .C2(new_n887), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT104), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n815), .B1(new_n774), .B2(new_n779), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n780), .A2(new_n814), .A3(new_n812), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n799), .A2(new_n500), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n799), .A2(new_n500), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n901), .A2(new_n904), .A3(new_n905), .A4(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n895), .B2(new_n898), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n900), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n900), .B2(new_n911), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n914), .A2(new_n913), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n881), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n900), .A2(new_n909), .A3(new_n911), .ZN(new_n919));
  INV_X1    g494(.A(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT106), .B1(new_n920), .B2(new_n899), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n909), .A2(new_n922), .A3(new_n895), .A4(new_n898), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n919), .A2(new_n921), .A3(new_n881), .A4(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n918), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g504(.A1(new_n868), .A2(new_n614), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n639), .B(KEYINPUT107), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(new_n870), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n582), .B1(new_n569), .B2(new_n571), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n638), .A2(KEYINPUT109), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G299), .B2(new_n627), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n638), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT108), .B1(G299), .B2(new_n627), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n935), .B(new_n937), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(G290), .A2(G288), .ZN(new_n944));
  NOR2_X1   g519(.A1(G290), .A2(G288), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(G305), .B1(new_n510), .B2(new_n529), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n727), .A2(new_n590), .A3(new_n592), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n947), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n946), .A2(new_n948), .A3(new_n947), .A4(KEYINPUT110), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n938), .B1(new_n638), .B2(new_n934), .ZN(new_n958));
  NAND3_X1  g533(.A1(G299), .A2(KEYINPUT108), .A3(new_n627), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT41), .A3(new_n935), .A4(new_n937), .ZN(new_n961));
  NAND2_X1  g536(.A1(G299), .A2(new_n627), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n937), .A2(new_n935), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT41), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n933), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n943), .A2(new_n957), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n957), .B1(new_n943), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n955), .A2(new_n956), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n931), .B1(new_n972), .B2(G868), .ZN(G295));
  AOI21_X1  g548(.A(new_n931), .B1(new_n972), .B2(G868), .ZN(G331));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n527), .A2(G89), .ZN(new_n976));
  INV_X1    g551(.A(new_n538), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n536), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G301), .B1(new_n978), .B2(new_n534), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n535), .A2(G171), .A3(new_n536), .A4(new_n539), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n869), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n942), .B1(new_n982), .B2(new_n964), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n869), .A2(new_n979), .A3(new_n980), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n560), .A2(new_n875), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n986), .A3(new_n864), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT41), .A3(new_n963), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n983), .A2(new_n984), .A3(new_n954), .A4(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n941), .A2(new_n985), .A3(new_n987), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n954), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n966), .A2(new_n988), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n990), .A2(new_n925), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n964), .B1(new_n985), .B2(new_n987), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n954), .B1(new_n997), .B2(new_n941), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n988), .A2(KEYINPUT41), .A3(new_n963), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT112), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n961), .A2(new_n965), .B1(new_n985), .B2(new_n987), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n991), .ZN(new_n1004));
  AOI21_X1  g579(.A(G37), .B1(new_n1004), .B2(new_n993), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n954), .B1(new_n1003), .B2(new_n991), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n975), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n996), .A2(new_n1011), .A3(new_n1006), .A4(new_n1000), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1005), .A2(new_n1000), .A3(new_n1006), .A4(new_n990), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1009), .B1(new_n975), .B2(new_n1015), .ZN(G397));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n500), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT114), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n495), .B2(new_n499), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1024));
  INV_X1    g599(.A(G40), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n469), .A2(new_n473), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1018), .B2(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1020), .A2(KEYINPUT117), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1956), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1020), .A2(KEYINPUT45), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1034), .A2(new_n1026), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1018), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT56), .B(G2072), .Z(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1033), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n934), .B(KEYINPUT57), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1042), .B(KEYINPUT119), .Z(new_n1044));
  INV_X1    g619(.A(new_n1033), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1040), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(KEYINPUT118), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT50), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1018), .A2(new_n1030), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1026), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n828), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1019), .A2(new_n1026), .A3(new_n1022), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n801), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n638), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1043), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1043), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(KEYINPUT60), .A3(new_n1057), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n627), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1055), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1996), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1037), .A2(new_n1072), .A3(new_n1026), .A4(new_n1034), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT120), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT120), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n560), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1078), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n560), .B(new_n1080), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1041), .A2(new_n1060), .A3(new_n1042), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1054), .A2(KEYINPUT60), .A3(new_n638), .A4(new_n1057), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1059), .B1(new_n1068), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G286), .A2(G8), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT122), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1053), .ZN(new_n1088));
  INV_X1    g663(.A(G2084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1023), .A2(new_n1036), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1035), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1088), .A2(new_n1089), .B1(new_n1091), .B2(new_n842), .ZN(new_n1092));
  INV_X1    g667(.A(G8), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT51), .B(new_n1087), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1092), .A2(new_n1087), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n842), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1089), .B(new_n1026), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1087), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1095), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1038), .A2(new_n724), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1024), .A2(new_n1032), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(G2090), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G8), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n587), .A2(new_n594), .A3(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT55), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n587), .A2(new_n594), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1053), .A2(new_n758), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1038), .B2(G2078), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(G301), .B(KEYINPUT54), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1038), .ZN(new_n1118));
  INV_X1    g693(.A(G2078), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1119), .A2(KEYINPUT123), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(KEYINPUT123), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1114), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1090), .A2(new_n1035), .A3(KEYINPUT53), .A4(new_n1119), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1113), .A2(new_n1115), .A3(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1116), .A2(new_n1123), .B1(new_n1125), .B2(new_n1117), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1056), .A2(new_n1093), .ZN(new_n1127));
  INV_X1    g702(.A(G1976), .ZN(new_n1128));
  OR2_X1    g703(.A1(G288), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(G288), .B2(new_n1128), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1055), .A2(G8), .A3(new_n1129), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT52), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G305), .B(G1981), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT49), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT116), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1055), .B(G8), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1131), .B(new_n1133), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1103), .B1(new_n1053), .B2(G2090), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1109), .A2(KEYINPUT115), .A3(new_n1110), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT115), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1141), .B(G8), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  AND4_X1   g719(.A1(new_n1112), .A2(new_n1126), .A3(new_n1140), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1085), .A2(new_n1102), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1140), .A2(new_n1144), .A3(new_n1112), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1099), .A2(G168), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1141), .A2(G8), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1111), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1151), .A2(new_n1153), .A3(new_n1144), .A4(new_n1140), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1125), .A2(G171), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1094), .A2(new_n1095), .A3(new_n1101), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1144), .A2(new_n1139), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G288), .A2(G1976), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(G1981), .B2(G305), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1127), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1146), .A2(new_n1155), .A3(new_n1161), .A4(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n780), .B(G1996), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n799), .B(new_n801), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n742), .B(new_n744), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G290), .B(new_n749), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1037), .A2(new_n1027), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1167), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1072), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT46), .Z(new_n1179));
  INV_X1    g754(.A(new_n1175), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n780), .B2(new_n1169), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1183));
  XNOR2_X1  g758(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n742), .A2(new_n744), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT124), .Z(new_n1186));
  OAI22_X1  g761(.A1(new_n1186), .A2(new_n1170), .B1(G2067), .B2(new_n799), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1175), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT48), .ZN(new_n1190));
  OR3_X1    g765(.A1(new_n1180), .A2(G1986), .A3(G290), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1184), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1177), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g770(.A(new_n1010), .ZN(new_n1197));
  AND2_X1   g771(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g774(.A(new_n714), .ZN(new_n1201));
  XNOR2_X1  g775(.A(new_n711), .B(new_n1201), .ZN(new_n1202));
  AND2_X1   g776(.A1(new_n670), .A2(G319), .ZN(new_n1203));
  NAND4_X1  g777(.A1(new_n1202), .A2(new_n1203), .A3(new_n691), .A4(KEYINPUT126), .ZN(new_n1204));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1205));
  NAND4_X1  g779(.A1(new_n670), .A2(new_n689), .A3(G319), .A4(new_n690), .ZN(new_n1206));
  OAI21_X1  g780(.A(new_n1205), .B1(G229), .B2(new_n1206), .ZN(new_n1207));
  AND2_X1   g781(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1208), .B1(new_n917), .B2(new_n926), .ZN(new_n1209));
  INV_X1    g783(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n1200), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1212));
  NOR3_X1   g786(.A1(new_n1015), .A2(new_n1212), .A3(new_n1209), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1213), .ZN(G308));
  NAND3_X1  g788(.A1(new_n1200), .A2(new_n1210), .A3(KEYINPUT127), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n1212), .B1(new_n1015), .B2(new_n1209), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1216), .ZN(G225));
endmodule


