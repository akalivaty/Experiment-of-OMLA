

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  NOR2_X1 U323 ( .A1(n506), .A2(n452), .ZN(n568) );
  AND2_X1 U324 ( .A1(n391), .A2(n390), .ZN(n392) );
  NOR2_X1 U325 ( .A1(n558), .A2(n387), .ZN(n388) );
  INV_X1 U326 ( .A(G78GAT), .ZN(n304) );
  XNOR2_X1 U327 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U328 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U329 ( .A(KEYINPUT36), .B(n567), .Z(n588) );
  INV_X1 U330 ( .A(G183GAT), .ZN(n454) );
  XNOR2_X1 U331 ( .A(KEYINPUT114), .B(n460), .ZN(n545) );
  XNOR2_X1 U332 ( .A(n454), .B(KEYINPUT124), .ZN(n455) );
  XNOR2_X1 U333 ( .A(n463), .B(KEYINPUT50), .ZN(n464) );
  XNOR2_X1 U334 ( .A(n456), .B(n455), .ZN(G1350GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n292) );
  XNOR2_X1 U336 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n309) );
  XNOR2_X1 U338 ( .A(G71GAT), .B(G57GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n293), .B(KEYINPUT13), .ZN(n382) );
  XOR2_X1 U340 ( .A(G127GAT), .B(G155GAT), .Z(n433) );
  XNOR2_X1 U341 ( .A(n382), .B(n433), .ZN(n294) );
  AND2_X1 U342 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  NAND2_X1 U343 ( .A1(n294), .A2(n295), .ZN(n299) );
  INV_X1 U344 ( .A(n294), .ZN(n297) );
  INV_X1 U345 ( .A(n295), .ZN(n296) );
  NAND2_X1 U346 ( .A1(n297), .A2(n296), .ZN(n298) );
  NAND2_X1 U347 ( .A1(n299), .A2(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n300), .B(KEYINPUT83), .Z(n303) );
  XNOR2_X1 U349 ( .A(G8GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n301), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U351 ( .A(n400), .B(KEYINPUT82), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G1GAT), .Z(n341) );
  XNOR2_X1 U354 ( .A(G22GAT), .B(n341), .ZN(n305) );
  XOR2_X1 U355 ( .A(n309), .B(n308), .Z(n494) );
  INV_X1 U356 ( .A(n494), .ZN(n584) );
  XNOR2_X1 U357 ( .A(KEYINPUT111), .B(n584), .ZN(n462) );
  XOR2_X1 U358 ( .A(G120GAT), .B(KEYINPUT0), .Z(n311) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n442) );
  XOR2_X1 U361 ( .A(n442), .B(G71GAT), .Z(n313) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n331) );
  XOR2_X1 U364 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT17), .B(KEYINPUT88), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(n316), .B(KEYINPUT87), .Z(n318) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(KEYINPUT89), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n398) );
  XOR2_X1 U370 ( .A(KEYINPUT86), .B(G190GAT), .Z(n320) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(G99GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U373 ( .A(G127GAT), .B(G176GAT), .Z(n322) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G183GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U376 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n324) );
  XNOR2_X1 U377 ( .A(KEYINPUT64), .B(KEYINPUT90), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U379 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U381 ( .A(n398), .B(n329), .Z(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n506) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n332), .B(G29GAT), .ZN(n333) );
  XOR2_X1 U385 ( .A(n333), .B(KEYINPUT7), .Z(n335) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(G50GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n361) );
  XOR2_X1 U388 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n337) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G8GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n361), .B(n338), .ZN(n349) );
  XOR2_X1 U392 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n340) );
  XNOR2_X1 U393 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U395 ( .A(G113GAT), .B(G197GAT), .Z(n343) );
  XOR2_X1 U396 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XNOR2_X1 U397 ( .A(n420), .B(n341), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U399 ( .A(n345), .B(n344), .Z(n347) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n575) );
  XNOR2_X1 U403 ( .A(n575), .B(KEYINPUT72), .ZN(n558) );
  XOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n351) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(G92GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n365) );
  XOR2_X1 U407 ( .A(KEYINPUT81), .B(KEYINPUT9), .Z(n353) );
  XNOR2_X1 U408 ( .A(KEYINPUT65), .B(KEYINPUT67), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n354), .B(KEYINPUT80), .Z(n356) );
  XOR2_X1 U411 ( .A(G190GAT), .B(G218GAT), .Z(n399) );
  XNOR2_X1 U412 ( .A(G134GAT), .B(n399), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U414 ( .A(G99GAT), .B(G85GAT), .Z(n373) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(n373), .Z(n358) );
  NAND2_X1 U416 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U418 ( .A(n360), .B(n359), .Z(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT79), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U420 ( .A(n361), .B(n426), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X2 U422 ( .A(n365), .B(n364), .Z(n567) );
  NOR2_X1 U423 ( .A1(n494), .A2(n588), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n366), .B(KEYINPUT45), .ZN(n386) );
  XOR2_X1 U425 ( .A(G92GAT), .B(G64GAT), .Z(n368) );
  XNOR2_X1 U426 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U428 ( .A(G176GAT), .B(n369), .Z(n397) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n371) );
  XNOR2_X1 U430 ( .A(G120GAT), .B(KEYINPUT77), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U432 ( .A(n373), .B(n372), .Z(n375) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U435 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n377) );
  XNOR2_X1 U436 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U439 ( .A(G78GAT), .B(G148GAT), .Z(n381) );
  XNOR2_X1 U440 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n412) );
  XNOR2_X1 U442 ( .A(n412), .B(n382), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n397), .B(n385), .ZN(n580) );
  NAND2_X1 U445 ( .A1(n386), .A2(n580), .ZN(n387) );
  XOR2_X1 U446 ( .A(KEYINPUT112), .B(n388), .Z(n395) );
  XNOR2_X1 U447 ( .A(KEYINPUT41), .B(n580), .ZN(n564) );
  NAND2_X1 U448 ( .A1(n575), .A2(n564), .ZN(n389) );
  XNOR2_X1 U449 ( .A(KEYINPUT46), .B(n389), .ZN(n391) );
  INV_X1 U450 ( .A(n567), .ZN(n390) );
  AND2_X1 U451 ( .A1(n462), .A2(n392), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(KEYINPUT47), .ZN(n394) );
  NAND2_X1 U453 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U454 ( .A(KEYINPUT48), .B(n396), .ZN(n457) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n406) );
  XOR2_X1 U456 ( .A(G197GAT), .B(KEYINPUT21), .Z(n425) );
  XNOR2_X1 U457 ( .A(n425), .B(n399), .ZN(n404) );
  XOR2_X1 U458 ( .A(G36GAT), .B(n400), .Z(n402) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n529) );
  NAND2_X1 U463 ( .A1(n457), .A2(n529), .ZN(n409) );
  XNOR2_X1 U464 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n407), .B(KEYINPUT54), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n572) );
  XOR2_X1 U467 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n411) );
  XNOR2_X1 U468 ( .A(G211GAT), .B(KEYINPUT22), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n416) );
  XOR2_X1 U470 ( .A(G204GAT), .B(n412), .Z(n414) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n430) );
  XOR2_X1 U474 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n418) );
  XNOR2_X1 U475 ( .A(G155GAT), .B(KEYINPUT91), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n419), .B(G218GAT), .Z(n422) );
  XNOR2_X1 U478 ( .A(G50GAT), .B(n420), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n423), .B(KEYINPUT2), .ZN(n441) );
  XOR2_X1 U482 ( .A(n424), .B(n441), .Z(n428) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n474) );
  XOR2_X1 U486 ( .A(G57GAT), .B(G85GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G141GAT), .B(G148GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U489 ( .A(n434), .B(n433), .Z(n436) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(G162GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n438) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n446) );
  NAND2_X1 U499 ( .A1(G225GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT6), .B(n447), .Z(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n571) );
  INV_X1 U503 ( .A(n571), .ZN(n527) );
  NOR2_X1 U504 ( .A1(n474), .A2(n527), .ZN(n450) );
  AND2_X1 U505 ( .A1(n572), .A2(n450), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  INV_X1 U507 ( .A(n568), .ZN(n453) );
  NOR2_X1 U508 ( .A1(n462), .A2(n453), .ZN(n456) );
  XOR2_X1 U509 ( .A(n529), .B(KEYINPUT27), .Z(n476) );
  NOR2_X1 U510 ( .A1(n476), .A2(n571), .ZN(n468) );
  NAND2_X1 U511 ( .A1(n457), .A2(n468), .ZN(n548) );
  NOR2_X1 U512 ( .A1(n506), .A2(n548), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT113), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n474), .B(KEYINPUT28), .ZN(n535) );
  NOR2_X1 U515 ( .A1(n459), .A2(n535), .ZN(n460) );
  INV_X1 U516 ( .A(n545), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n465) );
  INV_X1 U518 ( .A(G127GAT), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n465), .B(n464), .ZN(G1342GAT) );
  NAND2_X1 U520 ( .A1(n558), .A2(n580), .ZN(n497) );
  XOR2_X1 U521 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n467) );
  OR2_X1 U522 ( .A1(n494), .A2(n567), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n467), .B(n466), .ZN(n483) );
  NAND2_X1 U524 ( .A1(n506), .A2(n468), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n535), .A2(n469), .ZN(n481) );
  INV_X1 U526 ( .A(n506), .ZN(n532) );
  NAND2_X1 U527 ( .A1(n529), .A2(n532), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT97), .B(n470), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n474), .A2(n471), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT98), .B(n472), .Z(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT25), .B(n473), .ZN(n478) );
  NAND2_X1 U532 ( .A1(n474), .A2(n506), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT26), .ZN(n574) );
  NOR2_X1 U534 ( .A1(n476), .A2(n574), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n478), .A2(n477), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n527), .A2(n479), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n493) );
  INV_X1 U538 ( .A(n493), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n483), .A2(n482), .ZN(n515) );
  NOR2_X1 U540 ( .A1(n497), .A2(n515), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(n484), .Z(n491) );
  NAND2_X1 U542 ( .A1(n527), .A2(n491), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(n485), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n491), .A2(n529), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT100), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n491), .A2(n532), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n535), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U553 ( .A1(n588), .A2(n493), .ZN(n495) );
  NAND2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n496) );
  XOR2_X1 U555 ( .A(KEYINPUT37), .B(n496), .Z(n526) );
  NOR2_X1 U556 ( .A1(n526), .A2(n497), .ZN(n499) );
  XNOR2_X1 U557 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n510) );
  NOR2_X1 U559 ( .A1(n510), .A2(n571), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  INV_X1 U563 ( .A(n529), .ZN(n503) );
  NOR2_X1 U564 ( .A1(n510), .A2(n503), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  XNOR2_X1 U567 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n508) );
  NOR2_X1 U568 ( .A1(n506), .A2(n510), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U570 ( .A(G43GAT), .B(n509), .Z(G1330GAT) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n513) );
  INV_X1 U572 ( .A(n535), .ZN(n511) );
  NOR2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n517) );
  INV_X1 U576 ( .A(n575), .ZN(n514) );
  NAND2_X1 U577 ( .A1(n564), .A2(n514), .ZN(n525) );
  NOR2_X1 U578 ( .A1(n525), .A2(n515), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n522), .A2(n527), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n518), .Z(G1332GAT) );
  XOR2_X1 U582 ( .A(G64GAT), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U583 ( .A1(n522), .A2(n529), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n532), .A2(n522), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U588 ( .A1(n522), .A2(n535), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n527), .A2(n536), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT108), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  XOR2_X1 U596 ( .A(G99GAT), .B(KEYINPUT109), .Z(n534) );
  NAND2_X1 U597 ( .A1(n536), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n538) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U602 ( .A(G106GAT), .B(n539), .Z(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT115), .Z(n541) );
  NAND2_X1 U604 ( .A1(n545), .A2(n558), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U607 ( .A1(n564), .A2(n545), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U611 ( .A1(n567), .A2(n545), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n574), .A2(n548), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n575), .A2(n556), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n551) );
  NAND2_X1 U617 ( .A1(n556), .A2(n564), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT117), .Z(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n584), .A2(n556), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n556), .A2(n567), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .Z(n560) );
  NAND2_X1 U627 ( .A1(n568), .A2(n558), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n562) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(n563), .Z(n566) );
  NAND2_X1 U633 ( .A1(n568), .A2(n564), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .Z(n577) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n583), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n583), .ZN(n587) );
  OR2_X1 U647 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

