//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  XNOR2_X1  g000(.A(KEYINPUT99), .B(G952), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT21), .B(G898), .Z(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G214), .B1(G237), .B2(G902), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n194), .B(KEYINPUT88), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G116), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(G113), .C1(KEYINPUT5), .C2(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT2), .B(G113), .Z(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n198), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G104), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n213), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n213), .B1(new_n206), .B2(new_n208), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n215), .B1(new_n214), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n222), .B(G101), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n213), .A3(new_n216), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n222), .B1(new_n228), .B2(G101), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT80), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n223), .B2(new_n225), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT79), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .A4(new_n226), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n203), .B(new_n198), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n239));
  OAI211_X1 g053(.A(G101), .B(new_n239), .C1(new_n223), .C2(new_n225), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n228), .A2(KEYINPUT82), .A3(G101), .A4(new_n239), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n221), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n197), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n245), .B2(KEYINPUT89), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n243), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n237), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n235), .B2(new_n230), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n252), .A2(new_n253), .A3(new_n221), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n247), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT90), .B(G224), .Z(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G953), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(KEYINPUT64), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n262), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n261), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n265), .A2(G146), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT65), .B(G143), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n260), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n261), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT0), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT64), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n263), .A2(G143), .ZN(new_n280));
  AOI21_X1  g094(.A(G146), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n275), .B(new_n278), .C1(new_n281), .C2(new_n268), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n258), .B1(new_n274), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n269), .B1(new_n272), .B2(G146), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n285));
  OAI21_X1  g099(.A(G128), .B1(new_n271), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n280), .A3(G146), .ZN(new_n287));
  INV_X1    g101(.A(new_n271), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n277), .A2(KEYINPUT1), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n287), .A2(new_n292), .A3(new_n288), .A4(new_n289), .ZN(new_n293));
  AOI221_X4 g107(.A(G125), .B1(new_n284), .B2(new_n286), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n257), .B1(new_n283), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n275), .B1(new_n281), .B2(new_n268), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n287), .A2(new_n288), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n259), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n282), .ZN(new_n299));
  OAI21_X1  g113(.A(G125), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n291), .A2(new_n293), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n284), .A2(new_n286), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n258), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n257), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n253), .B1(new_n252), .B2(new_n221), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n245), .A2(KEYINPUT89), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n197), .A4(new_n248), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n255), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n221), .B(new_n248), .C1(new_n236), .C2(new_n244), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT7), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n283), .B2(new_n294), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n300), .A2(new_n303), .A3(KEYINPUT7), .A4(new_n304), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n205), .A2(KEYINPUT91), .A3(new_n217), .A4(new_n219), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT91), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n204), .B(new_n202), .C1(new_n220), .C2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n246), .B(KEYINPUT8), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AND4_X1   g133(.A1(new_n295), .A2(new_n313), .A3(new_n314), .A4(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT92), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n311), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n295), .A2(new_n313), .A3(new_n314), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT92), .ZN(new_n324));
  AOI21_X1  g138(.A(G902), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n310), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n310), .B2(new_n325), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n193), .B(new_n196), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT9), .B(G234), .ZN(new_n330));
  INV_X1    g144(.A(G217), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n330), .A2(new_n331), .A3(G953), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n272), .A2(G128), .ZN(new_n333));
  INV_X1    g147(.A(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n277), .A2(G143), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G116), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n207), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n333), .A2(KEYINPUT13), .A3(new_n335), .ZN(new_n339));
  OAI21_X1  g153(.A(G134), .B1(new_n333), .B2(KEYINPUT13), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n336), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G122), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G116), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n207), .B1(new_n343), .B2(KEYINPUT14), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(new_n336), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n332), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(new_n348), .A3(new_n332), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT98), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G478), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT15), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n357), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G475), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n354), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT96), .ZN(new_n364));
  XNOR2_X1  g178(.A(G113), .B(G122), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n212), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT74), .B1(new_n258), .B2(G140), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n258), .A2(G140), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT19), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n258), .A2(G140), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT19), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n262), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT95), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(KEYINPUT16), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT16), .B1(new_n369), .B2(G125), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n262), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  INV_X1    g199(.A(G953), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n272), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n385), .A2(new_n386), .A3(G143), .A4(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G131), .ZN(new_n391));
  INV_X1    g205(.A(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n394), .B2(KEYINPUT94), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n380), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n390), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT93), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n372), .B2(G146), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n372), .A2(new_n401), .A3(G146), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n375), .A2(new_n371), .A3(new_n262), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n400), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n366), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  AOI211_X1 g221(.A(G146), .B(new_n382), .C1(new_n372), .C2(KEYINPUT16), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n384), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n392), .B1(new_n388), .B2(new_n389), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT17), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n409), .B(new_n411), .C1(KEYINPUT17), .C2(new_n394), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n366), .A3(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n364), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n416));
  INV_X1    g230(.A(new_n393), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT94), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  INV_X1    g232(.A(new_n384), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n397), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n378), .B(KEYINPUT95), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n406), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n366), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n416), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n415), .B1(new_n425), .B2(KEYINPUT20), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n413), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n427), .A2(new_n416), .A3(new_n428), .A4(new_n364), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n412), .A2(new_n406), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n423), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n413), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n354), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G475), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n329), .A2(new_n361), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n334), .B2(G137), .ZN(new_n439));
  INV_X1    g253(.A(G137), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT11), .A3(G134), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n334), .A2(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT66), .A2(G131), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n443), .B(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n273), .B1(new_n284), .B2(new_n275), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n446), .B(new_n282), .C1(new_n447), .C2(new_n259), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n291), .A2(new_n293), .B1(new_n284), .B2(new_n286), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n392), .B1(G134), .B2(new_n440), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n443), .A2(new_n392), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n237), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n443), .B(new_n444), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n298), .A2(new_n454), .A3(new_n299), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n301), .B2(new_n302), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT30), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n448), .B(new_n458), .C1(new_n449), .C2(new_n451), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n453), .B1(new_n460), .B2(new_n237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n385), .A2(new_n386), .A3(G210), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n462), .B(KEYINPUT27), .Z(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G101), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(KEYINPUT29), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n237), .B1(new_n452), .B2(KEYINPUT68), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n455), .A2(new_n456), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT28), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n238), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n237), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n473), .A2(new_n477), .A3(new_n465), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n354), .B1(new_n468), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n473), .A2(KEYINPUT70), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT70), .B1(new_n473), .B2(new_n477), .ZN(new_n481));
  AND4_X1   g295(.A1(KEYINPUT29), .A2(new_n480), .A3(new_n466), .A4(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G472), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(G472), .A2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n465), .B1(new_n473), .B2(new_n477), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT31), .B1(new_n461), .B2(new_n466), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n238), .B1(new_n457), .B2(new_n459), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  NOR4_X1   g303(.A1(new_n488), .A2(new_n453), .A3(new_n489), .A4(new_n465), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n486), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n486), .B(KEYINPUT69), .C1(new_n487), .C2(new_n490), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n485), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT32), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI211_X1 g311(.A(KEYINPUT32), .B(new_n485), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n483), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G221), .ZN(new_n500));
  INV_X1    g314(.A(new_n330), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n354), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT76), .Z(new_n503));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n292), .B1(new_n273), .B2(new_n289), .ZN(new_n508));
  INV_X1    g322(.A(new_n293), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n220), .B(new_n302), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G128), .B1(new_n281), .B2(new_n285), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n291), .A2(new_n293), .B1(new_n511), .B2(new_n297), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n220), .B2(new_n512), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n505), .B(new_n507), .C1(new_n513), .C2(new_n446), .ZN(new_n514));
  AND4_X1   g328(.A1(KEYINPUT85), .A2(new_n513), .A3(new_n504), .A4(new_n446), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n297), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n220), .B1(new_n301), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n217), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n518), .A2(new_n519), .B1(new_n449), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n298), .A2(new_n299), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n250), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n236), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n454), .B(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n386), .A2(G227), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT77), .ZN(new_n528));
  XNOR2_X1  g342(.A(G110), .B(G140), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n516), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n236), .A2(new_n523), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n449), .A2(new_n520), .ZN(new_n534));
  INV_X1    g348(.A(new_n518), .ZN(new_n535));
  INV_X1    g349(.A(new_n519), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n533), .A2(new_n537), .A3(new_n525), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT86), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n524), .B2(new_n454), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n537), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT86), .A3(new_n446), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n532), .B1(new_n543), .B2(new_n531), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n354), .ZN(new_n546));
  NAND2_X1  g360(.A1(G469), .A2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT86), .B1(new_n541), .B2(new_n446), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n539), .B(new_n454), .C1(new_n533), .C2(new_n537), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n526), .B(new_n531), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n505), .B1(new_n513), .B2(new_n446), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n506), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n513), .A2(KEYINPUT85), .A3(new_n504), .A4(new_n446), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n530), .B1(new_n557), .B2(new_n538), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n552), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n552), .B2(new_n558), .ZN(new_n560));
  OAI21_X1  g374(.A(G469), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n503), .B1(new_n549), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n331), .B1(G234), .B2(new_n354), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n200), .B2(G128), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT73), .B1(new_n200), .B2(G128), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G110), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT71), .B1(new_n200), .B2(G128), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT71), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n277), .A3(G119), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n200), .A2(G128), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT72), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n570), .A2(new_n572), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G110), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n569), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n409), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n382), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n404), .B1(new_n582), .B2(new_n262), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n566), .A2(new_n567), .ZN(new_n584));
  INV_X1    g398(.A(G110), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n566), .A2(new_n567), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n578), .A2(new_n579), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n564), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n587), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(new_n419), .A3(new_n404), .ZN(new_n592));
  OAI221_X1 g406(.A(new_n569), .B1(new_n578), .B2(new_n579), .C1(new_n384), .C2(new_n408), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT75), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n386), .A2(G221), .A3(G234), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n590), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n592), .A2(new_n593), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n564), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT25), .B1(new_n602), .B2(new_n354), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT25), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n604), .B(G902), .C1(new_n598), .C2(new_n601), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n563), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n563), .A2(G902), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n437), .A2(new_n499), .A3(new_n562), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AND2_X1   g426(.A1(new_n562), .A2(new_n610), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n350), .A2(new_n351), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n352), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n616), .A2(G478), .A3(new_n354), .A4(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n356), .B1(new_n614), .B2(G902), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT101), .B1(new_n436), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n362), .B1(new_n433), .B2(new_n354), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n426), .B2(new_n429), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n626), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n329), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n493), .A2(new_n494), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n354), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n495), .B1(new_n632), .B2(G472), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n613), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR2_X1   g450(.A1(new_n415), .A2(KEYINPUT20), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n428), .B1(new_n427), .B2(new_n364), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n435), .B(new_n361), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n329), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n613), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT102), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  OAI21_X1  g458(.A(new_n599), .B1(KEYINPUT36), .B2(new_n597), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n592), .A2(new_n593), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n608), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT103), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n606), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n437), .A2(new_n562), .A3(new_n633), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  OAI21_X1  g467(.A(new_n190), .B1(G900), .B2(new_n192), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n639), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(new_n196), .C1(new_n327), .C2(new_n328), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n310), .A2(new_n325), .ZN(new_n659));
  INV_X1    g473(.A(new_n326), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n310), .A2(new_n325), .A3(new_n326), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n196), .A4(new_n656), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(new_n499), .A3(new_n562), .A4(new_n650), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  AOI21_X1  g482(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT105), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n461), .A2(new_n466), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n354), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n497), .B2(new_n498), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT38), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n663), .B(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n361), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n626), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n606), .A3(new_n196), .A4(new_n649), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n676), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n654), .B(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n562), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n562), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n682), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(new_n272), .Z(G45));
  NOR3_X1   g504(.A1(new_n626), .A2(new_n622), .A3(new_n655), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n663), .A2(new_n196), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n499), .A2(new_n562), .A3(new_n693), .A4(new_n650), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NOR3_X1   g509(.A1(new_n557), .A2(new_n538), .A3(new_n530), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n526), .B1(new_n550), .B2(new_n551), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n696), .B1(new_n697), .B2(new_n530), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n698), .B2(G902), .ZN(new_n699));
  INV_X1    g513(.A(new_n502), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n699), .A2(new_n546), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n499), .A2(new_n630), .A3(new_n610), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n499), .A2(new_n610), .A3(new_n640), .A4(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AND3_X1   g520(.A1(new_n626), .A2(new_n193), .A3(new_n679), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n499), .A2(new_n650), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n196), .B1(new_n327), .B2(new_n328), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n701), .A2(new_n710), .A3(KEYINPUT107), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n699), .A2(new_n546), .A3(new_n700), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n709), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  OAI211_X1 g531(.A(new_n196), .B(new_n680), .C1(new_n327), .C2(new_n328), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n663), .A2(new_n720), .A3(new_n196), .A4(new_n680), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n466), .B1(new_n480), .B2(new_n481), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n487), .A2(new_n490), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n484), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n493), .B2(new_n494), .ZN(new_n726));
  INV_X1    g540(.A(G472), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n610), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n699), .A2(new_n546), .A3(new_n700), .A4(new_n193), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  OAI211_X1 g546(.A(new_n650), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n733));
  INV_X1    g547(.A(new_n691), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT107), .B1(new_n701), .B2(new_n710), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n713), .A2(new_n709), .A3(new_n712), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n552), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n531), .B1(new_n516), .B2(new_n526), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n543), .B2(new_n531), .ZN(new_n743));
  OAI211_X1 g557(.A(G469), .B(new_n741), .C1(new_n743), .C2(new_n740), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n546), .A3(new_n547), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n327), .A2(new_n328), .A3(new_n195), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n745), .A2(new_n746), .A3(new_n700), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n499), .A3(new_n610), .A4(new_n691), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT111), .ZN(new_n751));
  INV_X1    g565(.A(new_n610), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n495), .B(new_n496), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(new_n483), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n691), .A4(new_n747), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n748), .A2(new_n756), .A3(new_n749), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n656), .A3(new_n747), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n623), .A2(new_n626), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n623), .A2(new_n765), .A3(new_n626), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n650), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n633), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT112), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n633), .A2(new_n767), .A3(new_n762), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n771), .B(new_n762), .C1(new_n633), .C2(new_n767), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n746), .A4(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n741), .C1(new_n743), .C2(new_n740), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(G469), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT45), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n547), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT46), .B(new_n547), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n546), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n700), .A3(new_n685), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n440), .ZN(G39));
  XNOR2_X1  g598(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n781), .A2(new_n700), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n746), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n499), .A2(new_n610), .A3(new_n788), .A4(new_n734), .ZN(new_n789));
  INV_X1    g603(.A(new_n546), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n777), .B2(new_n778), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n502), .B1(new_n791), .B2(new_n780), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(KEYINPUT47), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n787), .B(new_n789), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  OR3_X1    g610(.A1(new_n752), .A2(new_n503), .A3(new_n195), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n699), .A2(new_n546), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n763), .B(new_n797), .C1(new_n799), .C2(KEYINPUT49), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n676), .A3(new_n678), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n606), .A2(new_n649), .A3(new_n654), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n606), .A2(new_n649), .A3(new_n805), .A4(new_n654), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n807), .A2(new_n745), .A3(new_n700), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n722), .A3(new_n675), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n738), .A2(new_n667), .A3(new_n809), .A4(new_n694), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n811));
  INV_X1    g625(.A(new_n694), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n738), .A2(new_n667), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n738), .A2(new_n667), .A3(KEYINPUT116), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n809), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n811), .B1(new_n817), .B2(KEYINPUT52), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n626), .A2(new_n361), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n329), .A2(KEYINPUT115), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT115), .B1(new_n329), .B2(new_n820), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n613), .A2(new_n633), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n436), .A2(new_n623), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n329), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n562), .A2(new_n826), .A3(new_n610), .A4(new_n633), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(new_n611), .A3(new_n651), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n736), .A2(new_n737), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n499), .A2(new_n650), .A3(new_n707), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n705), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n702), .A2(new_n731), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n702), .A2(new_n731), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n716), .A4(new_n705), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n828), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n435), .B1(new_n637), .B2(new_n638), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n788), .A2(new_n361), .A3(new_n838), .A4(new_n655), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n499), .A3(new_n562), .A4(new_n650), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n735), .A2(new_n747), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n760), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n757), .A2(new_n755), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n843), .B2(new_n751), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n818), .A2(new_n819), .A3(new_n837), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n810), .B(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n837), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n849), .A3(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n819), .ZN(new_n851));
  INV_X1    g665(.A(new_n842), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n758), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n832), .A2(new_n833), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n611), .A2(new_n651), .A3(new_n827), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(KEYINPUT53), .A3(new_n824), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n818), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n850), .B1(KEYINPUT54), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n728), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n189), .A2(new_n764), .A3(new_n188), .A4(new_n766), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n195), .A3(new_n678), .A4(new_n701), .ZN(new_n864));
  OR2_X1    g678(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n701), .A3(new_n746), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n733), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n788), .A2(new_n713), .A3(new_n752), .A4(new_n190), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n676), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n436), .A3(new_n623), .ZN(new_n873));
  OR4_X1    g687(.A1(new_n866), .A2(new_n868), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n863), .A2(new_n746), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n787), .B1(new_n792), .B2(new_n794), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n798), .A2(new_n503), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n875), .B1(new_n874), .B2(new_n879), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n499), .A2(new_n610), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n869), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT48), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n872), .A2(new_n629), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n863), .A2(new_n715), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n188), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n860), .A2(new_n880), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n802), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n386), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n859), .A2(G210), .A3(G902), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n255), .A2(new_n309), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT119), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n306), .B(KEYINPUT55), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n894), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n859), .A2(G210), .A3(G902), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n859), .A2(new_n905), .A3(G210), .A4(G902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n901), .B1(new_n907), .B2(new_n899), .ZN(G51));
  XOR2_X1   g722(.A(new_n547), .B(KEYINPUT57), .Z(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n851), .A2(new_n910), .A3(new_n858), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n851), .B2(new_n858), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n544), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n859), .A2(G902), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n915), .A2(new_n776), .A3(new_n775), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n893), .B1(new_n914), .B2(new_n916), .ZN(G54));
  AOI22_X1  g731(.A1(new_n819), .A2(new_n848), .B1(new_n857), .B2(new_n818), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n354), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT121), .B1(new_n920), .B2(new_n427), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n893), .B1(new_n920), .B2(new_n427), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n923));
  INV_X1    g737(.A(new_n427), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n923), .B(new_n924), .C1(new_n915), .C2(new_n919), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(G60));
  NAND2_X1  g740(.A1(new_n616), .A2(new_n619), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT59), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n928), .B(new_n930), .C1(new_n911), .C2(new_n912), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n894), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n860), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n859), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n602), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n893), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n645), .A2(new_n647), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n859), .A2(new_n941), .A3(new_n937), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n940), .B(new_n942), .C1(KEYINPUT123), .C2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n918), .B2(new_n936), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n942), .A3(new_n894), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n936), .B1(new_n851), .B2(new_n858), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT123), .B(new_n894), .C1(new_n947), .C2(new_n602), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n943), .A2(new_n949), .ZN(G66));
  INV_X1    g764(.A(new_n256), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n386), .B1(new_n951), .B2(new_n191), .ZN(new_n952));
  INV_X1    g766(.A(new_n837), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n386), .ZN(new_n954));
  INV_X1    g768(.A(G898), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n897), .B1(new_n955), .B2(G953), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n758), .A2(new_n795), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n719), .A2(new_n721), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n882), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n700), .A3(new_n781), .A4(new_n685), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n760), .C1(new_n773), .C2(new_n782), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n813), .A2(new_n814), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n694), .A3(new_n816), .ZN(new_n964));
  NOR4_X1   g778(.A1(new_n958), .A2(new_n962), .A3(new_n964), .A4(G953), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n373), .A2(new_n377), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n460), .B(new_n967), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n965), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n758), .A2(new_n795), .ZN(new_n973));
  INV_X1    g787(.A(new_n962), .ZN(new_n974));
  INV_X1    g788(.A(new_n964), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n973), .A2(new_n974), .A3(new_n386), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT127), .B1(new_n976), .B2(new_n970), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n963), .A2(new_n689), .A3(new_n694), .A4(new_n816), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n815), .A2(new_n981), .A3(new_n689), .A4(new_n816), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n825), .A2(new_n820), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n562), .A2(new_n685), .A3(new_n746), .A4(new_n983), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n984), .A2(new_n882), .A3(KEYINPUT124), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT124), .B1(new_n984), .B2(new_n882), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n783), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n980), .A2(new_n982), .A3(new_n795), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n386), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n969), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT125), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n990), .A2(new_n993), .A3(new_n969), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n978), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n386), .B1(G227), .B2(G900), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n990), .B2(new_n969), .ZN(new_n998));
  AOI211_X1 g812(.A(KEYINPUT125), .B(new_n968), .C1(new_n989), .C2(new_n386), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n996), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n965), .B2(new_n971), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT126), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n998), .A2(new_n999), .A3(new_n1005), .A4(new_n1002), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n997), .B1(new_n1004), .B2(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND3_X1  g823(.A1(new_n973), .A2(new_n975), .A3(new_n974), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n953), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n465), .A3(new_n461), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n672), .A2(new_n467), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n845), .A2(new_n849), .A3(new_n1009), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1012), .A2(new_n894), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1009), .B1(new_n989), .B2(new_n953), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n461), .A2(new_n465), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(G57));
endmodule


