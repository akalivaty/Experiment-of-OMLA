//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n204), .A2(new_n205), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n203), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n210), .A2(new_n204), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n203), .A2(new_n213), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n225), .A3(KEYINPUT89), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT89), .B1(new_n223), .B2(new_n225), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n215), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G1gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT91), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(KEYINPUT90), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT16), .B1(new_n236), .B2(G1gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n230), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n233), .B1(new_n232), .B2(new_n238), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n229), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT92), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n238), .B(new_n248), .C1(G1gat), .C2(new_n230), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G8gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n239), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n223), .A2(new_n225), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n214), .B1(new_n256), .B2(new_n226), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT17), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n245), .B1(new_n260), .B2(KEYINPUT93), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n257), .A2(new_n258), .ZN(new_n263));
  AOI211_X1 g062(.A(KEYINPUT17), .B(new_n214), .C1(new_n256), .C2(new_n226), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(new_n252), .ZN(new_n266));
  NAND2_X1  g065(.A1(G229gat), .A2(G233gat), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n261), .A2(new_n266), .A3(KEYINPUT18), .A4(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT94), .B1(new_n229), .B2(new_n243), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(new_n244), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n267), .B(KEYINPUT13), .Z(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G113gat), .B(G141gat), .ZN(new_n273));
  INV_X1    g072(.A(G197gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT11), .B(G169gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT12), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n268), .A2(new_n272), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n261), .A2(new_n267), .A3(new_n266), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT18), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT95), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT95), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n281), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n272), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n278), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G1gat), .B(G29gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  AND2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n302));
  OR2_X1    g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(KEYINPUT75), .A3(new_n304), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n298), .A2(new_n299), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n302), .B(new_n310), .C1(new_n311), .C2(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n312), .A3(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G127gat), .ZN(new_n319));
  INV_X1    g118(.A(G127gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT69), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n325), .A3(G113gat), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n329), .A4(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT1), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n329), .A2(new_n337), .A3(new_n331), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n322), .B1(new_n342), .B2(KEYINPUT1), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n322), .B(new_n345), .C1(new_n342), .C2(KEYINPUT1), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n332), .A2(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n317), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n341), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n315), .A4(new_n316), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n349), .A2(new_n313), .A3(new_n350), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(KEYINPUT4), .B2(new_n357), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n356), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n355), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n313), .B1(new_n349), .B2(new_n350), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n367), .B(new_n363), .C1(new_n357), .C2(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n339), .A2(new_n340), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n339), .A2(new_n340), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n350), .B(new_n313), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n358), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n347), .A2(new_n374), .A3(new_n313), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT78), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n377), .A3(new_n358), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n354), .A2(new_n376), .A3(new_n378), .A4(new_n355), .ZN(new_n379));
  AND4_X1   g178(.A1(KEYINPUT80), .A2(new_n369), .A3(KEYINPUT5), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n366), .B2(new_n368), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT80), .B1(new_n382), .B2(new_n379), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n297), .B(new_n362), .C1(new_n380), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n297), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n379), .A3(KEYINPUT5), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n382), .A2(KEYINPUT80), .A3(new_n379), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n361), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n388), .B1(new_n393), .B2(KEYINPUT85), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n395), .B(new_n361), .C1(new_n391), .C2(new_n392), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n394), .A2(KEYINPUT86), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n362), .B1(new_n380), .B2(new_n383), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n297), .B1(new_n399), .B2(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(KEYINPUT85), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n387), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT38), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT74), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(G183gat), .A3(G190gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G183gat), .B(G190gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n407), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G169gat), .ZN(new_n413));
  INV_X1    g212(.A(G176gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(KEYINPUT23), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n418), .B(KEYINPUT25), .C1(G176gat), .C2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT64), .B(G176gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n421), .B2(new_n419), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n410), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n412), .A2(new_n420), .B1(KEYINPUT25), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n415), .A2(KEYINPUT26), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n415), .B1(new_n416), .B2(KEYINPUT26), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT67), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n427), .B2(new_n426), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT27), .B(G183gat), .ZN(new_n430));
  INV_X1    g229(.A(G190gat), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(KEYINPUT28), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n432), .A2(KEYINPUT28), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n434), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n429), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n424), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n438), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(new_n440), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n406), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G197gat), .B(G204gat), .ZN(new_n445));
  INV_X1    g244(.A(G211gat), .ZN(new_n446));
  INV_X1    g245(.A(G218gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n445), .B1(KEYINPUT22), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G211gat), .B(G218gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT74), .B1(new_n439), .B2(new_n440), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n444), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n441), .A2(new_n443), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n451), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G8gat), .B(G36gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(G64gat), .B(G92gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(KEYINPUT37), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n405), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n454), .A2(new_n456), .A3(new_n460), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n461), .B1(new_n457), .B2(KEYINPUT37), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n444), .A2(new_n451), .A3(new_n453), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n455), .A2(new_n452), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT37), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n405), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n403), .A2(new_n404), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT3), .B1(new_n307), .B2(new_n312), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n451), .B1(new_n476), .B2(KEYINPUT29), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT3), .B1(new_n452), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n313), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n477), .A2(new_n482), .B1(G228gat), .B2(G233gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n481), .B(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(G78gat), .B(G106gat), .Z(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G50gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n487), .B(KEYINPUT84), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT86), .B1(new_n394), .B2(new_n396), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n400), .A2(new_n398), .A3(new_n401), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n457), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n500));
  INV_X1    g299(.A(new_n354), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n360), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n355), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n388), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n357), .A2(new_n364), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT39), .B1(new_n506), .B2(new_n363), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n462), .A2(KEYINPUT30), .A3(new_n467), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n505), .B(KEYINPUT40), .C1(new_n503), .C2(new_n507), .ZN(new_n512));
  AND4_X1   g311(.A1(new_n500), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n496), .B1(new_n499), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n475), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n391), .A2(new_n392), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n297), .B1(new_n516), .B2(new_n362), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n404), .B1(new_n386), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n511), .A2(new_n500), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT82), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT82), .B1(new_n518), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n496), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G43gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n442), .B(new_n351), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(G227gat), .A3(G233gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(KEYINPUT32), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n527), .B(KEYINPUT32), .C1(new_n528), .C2(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n442), .B(new_n347), .ZN(new_n534));
  NAND2_X1  g333(.A1(G227gat), .A2(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT72), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n536), .A2(KEYINPUT34), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n534), .B2(new_n535), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n531), .A2(new_n541), .A3(new_n532), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(KEYINPUT36), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT73), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT73), .B1(new_n533), .B2(new_n542), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n549), .B2(KEYINPUT36), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n515), .A2(new_n522), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n495), .A2(new_n544), .A3(new_n543), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n520), .A2(new_n521), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT35), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n549), .A2(new_n519), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n386), .B1(new_n497), .B2(new_n498), .ZN(new_n557));
  INV_X1    g356(.A(new_n404), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n553), .A2(new_n554), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n292), .B1(new_n551), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G57gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT97), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT98), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n562), .A3(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n565), .A3(G57gat), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n564), .A2(new_n567), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  OR2_X1    g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n573), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n563), .A2(new_n566), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n575), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n575), .B1(new_n563), .B2(new_n566), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT96), .B1(new_n583), .B2(new_n578), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n577), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  AND2_X1   g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G127gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n577), .A2(new_n582), .A3(new_n584), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT99), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n243), .B1(new_n592), .B2(KEYINPUT21), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G155gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n594), .B(new_n598), .Z(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  OAI211_X1 g401(.A(KEYINPUT100), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT7), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n610), .A3(G85gat), .A4(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(G99gat), .ZN(new_n612));
  INV_X1    g411(.A(G106gat), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT8), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n605), .A2(new_n607), .A3(new_n611), .A4(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n603), .A2(new_n614), .A3(new_n604), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n606), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n265), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n257), .B2(new_n619), .ZN(new_n625));
  OR3_X1    g424(.A1(new_n621), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n622), .B1(new_n621), .B2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n626), .A2(new_n631), .A3(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n620), .B2(new_n585), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n618), .A2(new_n638), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n639), .A2(new_n585), .A3(new_n615), .A4(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n619), .A2(new_n590), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n637), .A2(new_n641), .A3(new_n642), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT103), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n641), .A3(new_n644), .ZN(new_n654));
  INV_X1    g453(.A(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n649), .A2(new_n656), .A3(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n599), .A2(new_n636), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n561), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n518), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n234), .ZN(G1324gat));
  INV_X1    g467(.A(new_n666), .ZN(new_n669));
  INV_X1    g468(.A(new_n519), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AND3_X1   g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n233), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT42), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(G1325gat));
  NAND2_X1  g479(.A1(new_n550), .A2(KEYINPUT105), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n682), .B(new_n545), .C1(new_n549), .C2(KEYINPUT36), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n666), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n549), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n666), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT106), .Z(G1326gat));
  NOR2_X1   g488(.A1(new_n666), .A2(new_n495), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n664), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n599), .A2(new_n636), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT107), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n561), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n518), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n208), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n522), .A2(KEYINPUT108), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n701), .B(new_n496), .C1(new_n520), .C2(new_n521), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n468), .A2(new_n472), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n468), .B1(KEYINPUT37), .B2(new_n457), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n467), .B(new_n704), .C1(new_n705), .C2(new_n405), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n557), .A2(new_n706), .A3(new_n558), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n499), .A2(new_n513), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n495), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n550), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n560), .B1(new_n703), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n636), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n551), .A2(new_n560), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n635), .A2(new_n713), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717));
  INV_X1    g516(.A(new_n599), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(new_n292), .A3(new_n664), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n716), .A2(new_n717), .A3(new_n697), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n714), .A2(new_n715), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n700), .A2(new_n515), .A3(new_n550), .A4(new_n702), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n635), .B1(new_n722), .B2(new_n560), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n721), .B(new_n719), .C1(new_n723), .C2(KEYINPUT44), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT109), .B1(new_n724), .B2(new_n518), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n725), .A3(G29gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n699), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT110), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n699), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1328gat));
  NAND3_X1  g530(.A1(new_n696), .A2(new_n209), .A3(new_n670), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT46), .Z(new_n733));
  OAI21_X1  g532(.A(G36gat), .B1(new_n724), .B2(new_n519), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1329gat));
  OAI21_X1  g534(.A(G43gat), .B1(new_n724), .B2(new_n550), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n696), .A2(new_n216), .A3(new_n549), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT47), .ZN(new_n738));
  OAI21_X1  g537(.A(G43gat), .B1(new_n724), .B2(new_n684), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g540(.A(new_n696), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n217), .B1(new_n742), .B2(new_n495), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n496), .A2(G50gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n724), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g545(.A1(new_n599), .A2(new_n636), .A3(new_n693), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n711), .A2(new_n292), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n518), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(new_n562), .ZN(G1332gat));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n519), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n748), .A2(new_n756), .A3(new_n684), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT111), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n748), .B2(new_n686), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT50), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1334gat));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n495), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g565(.A1(new_n718), .A2(new_n291), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n693), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n716), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n518), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n636), .A4(new_n767), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n635), .B(new_n768), .C1(new_n722), .C2(new_n560), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT113), .B1(new_n775), .B2(KEYINPUT51), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n711), .A2(new_n636), .A3(new_n767), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n697), .A2(new_n601), .A3(new_n664), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n771), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  NAND3_X1  g583(.A1(new_n716), .A2(new_n670), .A3(new_n769), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n693), .A2(new_n519), .A3(G92gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n788));
  INV_X1    g587(.A(new_n772), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n785), .B2(G92gat), .ZN(new_n793));
  INV_X1    g592(.A(new_n787), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n774), .B2(new_n781), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(KEYINPUT114), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n797), .B(new_n794), .C1(new_n774), .C2(new_n781), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n792), .B1(new_n796), .B2(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n770), .B2(new_n684), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n549), .A2(new_n612), .A3(new_n664), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT115), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n782), .B2(new_n802), .ZN(G1338gat));
  OR2_X1    g602(.A1(new_n788), .A2(new_n789), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n495), .A2(new_n693), .A3(G106gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n716), .A2(new_n496), .A3(new_n769), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(G106gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n808), .ZN(new_n810));
  INV_X1    g609(.A(new_n805), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n774), .B2(new_n781), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n807), .A2(new_n808), .B1(new_n810), .B2(new_n812), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n650), .A2(new_n814), .A3(new_n652), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n647), .B2(new_n648), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n645), .A2(new_n646), .A3(new_n655), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n660), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n663), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n291), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n261), .A2(new_n266), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n825), .A2(new_n267), .B1(new_n271), .B2(new_n270), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n277), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n287), .A2(new_n664), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n636), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n285), .B1(new_n281), .B2(new_n282), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n832), .A2(new_n280), .B1(new_n277), .B2(new_n826), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n635), .A2(new_n819), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n823), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n599), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n665), .A2(new_n292), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n496), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n686), .A2(new_n518), .A3(new_n670), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n327), .B1(new_n841), .B2(new_n291), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n518), .B1(new_n837), .B2(new_n838), .ZN(new_n843));
  INV_X1    g642(.A(new_n552), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n670), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n292), .A2(G113gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT116), .Z(G1340gat));
  AOI21_X1  g648(.A(G120gat), .B1(new_n846), .B2(new_n664), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n693), .A2(new_n325), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n841), .B2(new_n851), .ZN(G1341gat));
  INV_X1    g651(.A(new_n841), .ZN(new_n853));
  OAI21_X1  g652(.A(G127gat), .B1(new_n853), .B2(new_n599), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n846), .A2(new_n320), .A3(new_n718), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1342gat));
  OR4_X1    g655(.A1(G134gat), .A2(new_n845), .A3(new_n670), .A4(new_n635), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n853), .B2(new_n635), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1343gat));
  AOI21_X1  g660(.A(new_n495), .B1(new_n681), .B2(new_n683), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n843), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n670), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n292), .A2(G141gat), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n665), .A2(new_n292), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n822), .B1(new_n287), .B2(new_n290), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n815), .A2(new_n818), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n870), .A2(new_n873), .B1(new_n833), .B2(new_n664), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n835), .B1(new_n874), .B2(new_n636), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n875), .B2(new_n599), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n495), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n819), .B(new_n822), .C1(new_n287), .C2(new_n290), .ZN(new_n879));
  INV_X1    g678(.A(new_n828), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n635), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n718), .B1(new_n881), .B2(new_n835), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n878), .B(new_n496), .C1(new_n882), .C2(new_n869), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n550), .A2(new_n697), .A3(new_n519), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n877), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885), .B2(new_n292), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n291), .A2(new_n823), .A3(new_n873), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n636), .B1(new_n889), .B2(new_n828), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n599), .B1(new_n890), .B2(new_n836), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n838), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n878), .B1(new_n892), .B2(new_n496), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT118), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n895), .A3(new_n883), .A4(new_n884), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n291), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n867), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT119), .B1(new_n899), .B2(KEYINPUT58), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n866), .B1(new_n897), .B2(G141gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n868), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n887), .B1(new_n900), .B2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n864), .A2(new_n905), .A3(new_n664), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n878), .B1(new_n876), .B2(new_n495), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT120), .B(new_n878), .C1(new_n876), .C2(new_n495), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT57), .B(new_n496), .C1(new_n882), .C2(new_n869), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n664), .A3(new_n884), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n664), .A3(new_n896), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(new_n907), .A3(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n906), .B1(new_n915), .B2(new_n917), .ZN(G1345gat));
  INV_X1    g717(.A(G155gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n864), .A2(new_n919), .A3(new_n718), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n894), .A2(new_n718), .A3(new_n896), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(G1346gat));
  AND3_X1   g721(.A1(new_n894), .A2(new_n636), .A3(new_n896), .ZN(new_n923));
  INV_X1    g722(.A(G162gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n636), .A2(new_n924), .A3(new_n519), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n923), .A2(new_n924), .B1(new_n863), .B2(new_n925), .ZN(G1347gat));
  NAND2_X1  g725(.A1(new_n670), .A2(new_n518), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n686), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n839), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n413), .A3(new_n292), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n697), .B1(new_n837), .B2(new_n838), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n552), .A2(new_n519), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n291), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n930), .B1(new_n413), .B2(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(new_n414), .B1(new_n933), .B2(new_n693), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT121), .ZN(new_n938));
  INV_X1    g737(.A(new_n929), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n664), .A2(new_n421), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1349gat));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n430), .A3(new_n718), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n929), .A2(new_n943), .A3(new_n599), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n929), .B2(new_n599), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G183gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n929), .B2(new_n635), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n431), .A3(new_n636), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1351gat));
  AND2_X1   g751(.A1(new_n862), .A2(new_n670), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n931), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(KEYINPUT123), .A3(new_n931), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n291), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n927), .B1(new_n681), .B2(new_n683), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n913), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(new_n274), .A3(new_n292), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n959), .A2(new_n962), .ZN(G1352gat));
  OAI21_X1  g762(.A(G204gat), .B1(new_n961), .B2(new_n693), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n693), .A2(G204gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n953), .A2(new_n931), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n964), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  NAND4_X1  g771(.A1(new_n956), .A2(new_n446), .A3(new_n718), .A4(new_n957), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT125), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n913), .A2(new_n718), .A3(new_n960), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n974), .B(new_n978), .C1(new_n980), .C2(new_n976), .ZN(G1354gat));
  NAND3_X1  g780(.A1(new_n958), .A2(new_n447), .A3(new_n636), .ZN(new_n982));
  OAI21_X1  g781(.A(G218gat), .B1(new_n961), .B2(new_n635), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


