//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933;
  OR2_X1    g000(.A1(KEYINPUT70), .A2(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT70), .A2(G237), .ZN(new_n188));
  AOI21_X1  g002(.A(G953), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G214), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT91), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT18), .B1(new_n192), .B2(KEYINPUT91), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT65), .B(G146), .ZN(new_n197));
  XNOR2_X1  g011(.A(G125), .B(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(new_n198), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n192), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(G131), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n192), .A2(KEYINPUT17), .A3(G131), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n207), .B(G146), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n192), .A2(G131), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n190), .B(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n195), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n204), .B(new_n209), .C1(new_n213), .C2(KEYINPUT17), .ZN(new_n214));
  XNOR2_X1  g028(.A(G113), .B(G122), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT93), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n203), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(KEYINPUT92), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n198), .B(KEYINPUT19), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n197), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n210), .A2(new_n212), .A3(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(new_n221), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n226), .A2(new_n203), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n219), .B1(new_n227), .B2(new_n217), .ZN(new_n228));
  INV_X1    g042(.A(G475), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n228), .A2(KEYINPUT20), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n219), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n217), .B1(new_n226), .B2(new_n203), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n229), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT20), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n217), .B1(new_n203), .B2(new_n214), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n230), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G475), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n231), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT15), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G478), .ZN(new_n242));
  XOR2_X1   g056(.A(KEYINPUT9), .B(G234), .Z(new_n243));
  INV_X1    g057(.A(G953), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(G217), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G122), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G116), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G107), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(G116), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT14), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT94), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(KEYINPUT14), .B2(new_n249), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(G107), .ZN(new_n257));
  XNOR2_X1  g071(.A(G128), .B(G143), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(KEYINPUT13), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n191), .A2(G128), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n262), .B(G134), .C1(KEYINPUT13), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n259), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n252), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n246), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n261), .A2(new_n267), .A3(new_n246), .ZN(new_n270));
  AOI21_X1  g084(.A(G902), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT95), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n242), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n272), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n242), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n274), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n244), .A2(G952), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(G234), .B2(G237), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT21), .B(G898), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI211_X1 g095(.A(new_n230), .B(new_n244), .C1(G234), .C2(G237), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR3_X1    g097(.A1(new_n240), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  AOI22_X1  g099(.A1(KEYINPUT66), .A2(new_n285), .B1(new_n259), .B2(G137), .ZN(new_n286));
  OAI22_X1  g100(.A1(KEYINPUT66), .A2(new_n285), .B1(new_n259), .B2(G137), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  INV_X1    g102(.A(G137), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT11), .A4(G134), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT67), .A4(new_n290), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(G131), .A3(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n286), .A2(new_n287), .A3(new_n195), .A4(new_n290), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n293), .A2(new_n300), .A3(G131), .A4(new_n294), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n298), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n197), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n191), .A2(G146), .ZN(new_n306));
  INV_X1    g120(.A(G128), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT1), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n305), .B2(KEYINPUT1), .ZN(new_n310));
  MUX2_X1   g124(.A(G146), .B(new_n197), .S(new_n191), .Z(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n216), .A2(G107), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n216), .A2(G107), .ZN(new_n315));
  OAI21_X1  g129(.A(G101), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n250), .A3(G104), .ZN(new_n319));
  INV_X1    g133(.A(G101), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n317), .A2(new_n319), .A3(new_n320), .A4(new_n313), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n312), .A2(KEYINPUT10), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n312), .A2(KEYINPUT84), .A3(KEYINPUT10), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n305), .A2(new_n306), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n309), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n323), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n322), .B1(new_n332), .B2(new_n309), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(KEYINPUT10), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT0), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n307), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n311), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n307), .ZN(new_n344));
  INV_X1    g158(.A(new_n329), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n343), .A2(new_n344), .B1(new_n345), .B2(new_n342), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n317), .A2(new_n319), .A3(new_n313), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G101), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n350), .A3(G101), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(KEYINPUT4), .ZN(new_n352));
  INV_X1    g166(.A(new_n321), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(KEYINPUT81), .B2(new_n348), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n352), .A2(new_n354), .A3(KEYINPUT82), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT82), .B1(new_n352), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n346), .B(new_n349), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n304), .A2(new_n328), .A3(new_n340), .A4(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n244), .A2(G227), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n328), .A2(new_n340), .A3(new_n357), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n298), .A2(new_n301), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(KEYINPUT85), .A3(new_n361), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n364), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n334), .B1(new_n312), .B2(new_n323), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT12), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  AND4_X1   g188(.A1(KEYINPUT12), .A2(new_n373), .A3(new_n298), .A4(new_n301), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n358), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n361), .B(KEYINPUT80), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(G469), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n374), .A2(new_n375), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n362), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n361), .B1(new_n370), .B2(new_n358), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n380), .B(new_n230), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n380), .A2(new_n230), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n243), .ZN(new_n388));
  OAI21_X1  g202(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT78), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT79), .Z(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G214), .B1(G237), .B2(G902), .ZN(new_n393));
  XOR2_X1   g207(.A(new_n393), .B(KEYINPUT86), .Z(new_n394));
  XOR2_X1   g208(.A(G116), .B(G119), .Z(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT2), .B(G113), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(new_n349), .C1(new_n355), .C2(new_n356), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n399));
  INV_X1    g213(.A(G119), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G116), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n401), .B(KEYINPUT87), .Z(new_n402));
  OAI21_X1  g216(.A(G113), .B1(new_n395), .B2(new_n399), .ZN(new_n403));
  OAI22_X1  g217(.A1(new_n402), .A2(new_n403), .B1(new_n395), .B2(new_n396), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n404), .A2(new_n322), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(G110), .B(G122), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n407), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n411), .A3(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT88), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n398), .A2(new_n414), .A3(new_n411), .A4(new_n405), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n413), .A2(new_n415), .B1(new_n407), .B2(new_n406), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n410), .B1(new_n416), .B2(new_n409), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n346), .A2(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n312), .A2(new_n205), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT89), .B(G224), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n244), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n244), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n423), .A3(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G210), .B1(G237), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n422), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n418), .A2(new_n429), .A3(new_n423), .A4(new_n419), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n407), .B(KEYINPUT8), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n404), .A2(new_n322), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n405), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n413), .B2(new_n415), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n427), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n428), .B1(new_n427), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n394), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT90), .ZN(new_n443));
  INV_X1    g257(.A(new_n410), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n413), .A2(new_n415), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n408), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n446), .B2(KEYINPUT6), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n438), .B1(new_n447), .B2(new_n425), .ZN(new_n448));
  INV_X1    g262(.A(new_n428), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n439), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n394), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n284), .B(new_n392), .C1(new_n443), .C2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT72), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n289), .A2(G134), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n259), .A2(G137), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n312), .A2(new_n296), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n346), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n366), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n397), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n463));
  INV_X1    g277(.A(new_n459), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n369), .B2(new_n346), .ZN(new_n465));
  INV_X1    g279(.A(new_n397), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n346), .B1(new_n302), .B2(new_n303), .ZN(new_n468));
  AND4_X1   g282(.A1(new_n463), .A2(new_n468), .A3(new_n466), .A4(new_n459), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n462), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(G101), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n189), .A2(G210), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n459), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n461), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n397), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n465), .A2(new_n466), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n474), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT31), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT31), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n480), .A2(new_n484), .A3(new_n481), .A4(new_n474), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n476), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n487));
  NOR2_X1   g301(.A1(G472), .A2(G902), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G472), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n481), .A2(KEYINPUT28), .ZN(new_n493));
  INV_X1    g307(.A(new_n469), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n468), .A2(new_n459), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n397), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n474), .A2(KEYINPUT29), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT71), .B1(new_n470), .B2(new_n475), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT71), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n495), .A2(new_n502), .A3(new_n462), .A4(new_n474), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n480), .A2(new_n481), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n504), .B2(new_n475), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n492), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n455), .B1(new_n491), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n486), .A2(new_n488), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n500), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G472), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT72), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT76), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n400), .A2(G128), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT23), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(KEYINPUT23), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(G119), .C2(new_n307), .ZN(new_n521));
  XNOR2_X1  g335(.A(G119), .B(G128), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  OAI22_X1  g337(.A1(new_n521), .A2(G110), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n221), .A3(new_n199), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(G110), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n522), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n208), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n244), .A2(G221), .A3(G234), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n517), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT76), .A4(new_n534), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n529), .A2(new_n535), .A3(KEYINPUT75), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT75), .B1(new_n529), .B2(new_n535), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G217), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(G234), .B2(new_n230), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n540), .A2(G902), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n543), .A2(KEYINPUT77), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT25), .B1(new_n540), .B2(G902), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n538), .A2(new_n539), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n536), .A2(new_n537), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n230), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n549), .A3(new_n542), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n543), .A2(KEYINPUT77), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n454), .A2(new_n516), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  NAND2_X1  g369(.A1(new_n486), .A2(new_n230), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G472), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n509), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n558), .A2(new_n552), .A3(new_n392), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n440), .A2(new_n441), .ZN(new_n560));
  INV_X1    g374(.A(new_n393), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT96), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n563), .A2(KEYINPUT96), .ZN(new_n565));
  INV_X1    g379(.A(new_n270), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n268), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n269), .A2(KEYINPUT96), .A3(new_n563), .A4(new_n270), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(G478), .A3(new_n230), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n569), .A2(KEYINPUT97), .A3(G478), .A4(new_n230), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n573), .C1(G478), .C2(new_n271), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n240), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n283), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n559), .A2(new_n562), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT34), .B(G104), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G6));
  INV_X1    g393(.A(new_n240), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n277), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n283), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n559), .A2(new_n562), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT98), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G107), .Z(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G9));
  NAND2_X1  g400(.A1(new_n443), .A2(new_n453), .ZN(new_n587));
  INV_X1    g401(.A(new_n284), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n558), .A2(new_n392), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(new_n529), .Z(new_n591));
  OAI211_X1 g405(.A(new_n591), .B(new_n230), .C1(new_n541), .C2(G234), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n550), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT37), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G110), .ZN(G12));
  NOR2_X1   g413(.A1(new_n595), .A2(new_n392), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n508), .A2(new_n515), .A3(new_n562), .A4(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G900), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n279), .B1(new_n282), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n580), .A2(new_n277), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n307), .ZN(G30));
  XNOR2_X1  g421(.A(new_n451), .B(KEYINPUT38), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n481), .A2(new_n497), .A3(new_n475), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT100), .B1(new_n614), .B2(new_n609), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n615), .A3(new_n230), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n616), .A2(new_n617), .A3(G472), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n616), .B2(G472), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n512), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n608), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n603), .B(KEYINPUT39), .Z(new_n622));
  NAND3_X1  g436(.A1(new_n387), .A2(new_n391), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT40), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n593), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n240), .A2(new_n277), .A3(new_n393), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n621), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT102), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G143), .ZN(G45));
  AND3_X1   g444(.A1(new_n508), .A2(new_n515), .A3(new_n562), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n575), .A2(new_n603), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n600), .A4(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT103), .B1(new_n601), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G146), .ZN(G48));
  OR2_X1    g452(.A1(new_n382), .A2(new_n383), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n230), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(KEYINPUT104), .A3(G469), .ZN(new_n641));
  INV_X1    g455(.A(new_n390), .ZN(new_n642));
  NAND2_X1  g456(.A1(KEYINPUT104), .A2(G469), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n230), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n560), .A2(new_n645), .A3(new_n561), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n508), .A2(new_n646), .A3(new_n515), .A4(new_n553), .ZN(new_n647));
  INV_X1    g461(.A(new_n576), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT41), .B(G113), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G15));
  NAND4_X1  g465(.A1(new_n516), .A2(new_n553), .A3(new_n582), .A4(new_n646), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT105), .B(G116), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G18));
  INV_X1    g468(.A(new_n645), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n508), .A2(new_n515), .A3(new_n562), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n588), .A2(new_n596), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n400), .ZN(G21));
  NAND2_X1  g473(.A1(new_n627), .A2(new_n451), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n283), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n498), .A2(new_n474), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n483), .A2(new_n485), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n488), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n557), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n552), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n661), .A2(new_n655), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  AND3_X1   g482(.A1(new_n664), .A2(new_n557), .A3(new_n593), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n646), .A2(new_n669), .A3(new_n633), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT106), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G125), .ZN(G27));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n450), .A2(new_n439), .A3(new_n393), .ZN(new_n674));
  INV_X1    g488(.A(new_n387), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n674), .A2(new_n390), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n508), .A2(new_n515), .A3(new_n553), .A4(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n673), .B1(new_n677), .B2(new_n635), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n552), .B1(new_n512), .B2(new_n514), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(KEYINPUT42), .A3(new_n676), .A4(new_n633), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT107), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n678), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G131), .ZN(G33));
  OR2_X1    g500(.A1(new_n677), .A2(new_n605), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G134), .ZN(G36));
  NAND2_X1  g502(.A1(new_n574), .A2(new_n580), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n574), .A2(KEYINPUT43), .A3(new_n580), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n558), .B(new_n593), .C1(new_n693), .C2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n698));
  OR3_X1    g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n674), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n372), .A2(new_n378), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n702), .B(G469), .C1(new_n704), .C2(G902), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n384), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(KEYINPUT46), .A3(new_n386), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n390), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n709), .A2(new_n622), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n699), .A2(new_n700), .A3(new_n701), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT109), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n289), .ZN(G39));
  XOR2_X1   g527(.A(new_n709), .B(KEYINPUT47), .Z(new_n714));
  OR2_X1    g528(.A1(new_n516), .A2(new_n674), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n552), .A3(new_n633), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G140), .ZN(G42));
  NAND2_X1  g532(.A1(new_n641), .A2(new_n644), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT49), .ZN(new_n720));
  INV_X1    g534(.A(new_n394), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n552), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n391), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n608), .A2(new_n723), .A3(new_n689), .ZN(new_n724));
  INV_X1    g538(.A(new_n620), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n693), .A2(new_n279), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n666), .ZN(new_n728));
  INV_X1    g542(.A(new_n719), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n723), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n714), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n700), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n608), .A2(new_n393), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n727), .A2(new_n655), .A3(new_n666), .A4(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT50), .Z(new_n735));
  NAND2_X1  g549(.A1(new_n725), .A2(new_n553), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n700), .A2(new_n729), .A3(new_n279), .A4(new_n642), .ZN(new_n737));
  OR4_X1    g551(.A1(new_n240), .A2(new_n736), .A3(new_n574), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n694), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n669), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n732), .A2(new_n735), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n278), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n727), .A2(new_n646), .A3(new_n666), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n452), .B1(new_n451), .B2(new_n394), .ZN(new_n747));
  AOI211_X1 g561(.A(KEYINPUT90), .B(new_n721), .C1(new_n450), .C2(new_n439), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n576), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n587), .A2(KEYINPUT110), .A3(new_n576), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n559), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n652), .A2(new_n753), .A3(new_n554), .ZN(new_n754));
  OAI221_X1 g568(.A(new_n667), .B1(new_n656), .B2(new_n657), .C1(new_n648), .C2(new_n647), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n587), .A2(new_n559), .A3(new_n582), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n597), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n597), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n240), .A2(new_n277), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n674), .A2(new_n595), .A3(new_n392), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n508), .A2(new_n764), .A3(new_n515), .A4(new_n604), .ZN(new_n765));
  OAI22_X1  g579(.A1(new_n763), .A2(new_n765), .B1(new_n677), .B2(new_n605), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n676), .A2(new_n633), .A3(new_n669), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n685), .A2(new_n756), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n660), .A2(new_n390), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n603), .B(KEYINPUT113), .Z(new_n771));
  NOR3_X1   g585(.A1(new_n675), .A2(new_n593), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n620), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n670), .B(new_n773), .C1(new_n601), .C2(new_n605), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n637), .A2(KEYINPUT52), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(new_n637), .B2(new_n775), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n769), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n652), .A2(new_n753), .A3(new_n554), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n667), .B1(new_n647), .B2(new_n648), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n658), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n762), .A3(new_n768), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n684), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n683), .B1(new_n678), .B2(new_n680), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n777), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n670), .B1(new_n601), .B2(new_n605), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT112), .B(new_n670), .C1(new_n601), .C2(new_n605), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n637), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n781), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n637), .A2(KEYINPUT52), .A3(new_n775), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n790), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n779), .B1(new_n789), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n793), .A2(new_n794), .B1(new_n634), .B2(new_n636), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n637), .A2(new_n775), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n804), .A2(new_n796), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n681), .A2(KEYINPUT53), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n785), .A3(new_n808), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n803), .A2(new_n809), .A3(KEYINPUT54), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n745), .A2(new_n746), .A3(new_n800), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n736), .A2(new_n575), .A3(new_n737), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n739), .A2(new_n679), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(KEYINPUT48), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n813), .B(new_n815), .Z(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n814), .B2(KEYINPUT48), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(G952), .A2(G953), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n726), .B1(new_n818), .B2(new_n819), .ZN(G75));
  XNOR2_X1  g634(.A(new_n425), .B(KEYINPUT55), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(G210), .B(G902), .C1(new_n803), .C2(new_n809), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n447), .B(KEYINPUT116), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT117), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n823), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n823), .B2(new_n824), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n822), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(G210), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n780), .B1(new_n769), .B2(new_n778), .ZN(new_n832));
  INV_X1    g646(.A(new_n785), .ZN(new_n833));
  INV_X1    g647(.A(new_n808), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n798), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n831), .B(new_n230), .C1(new_n832), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n826), .B1(new_n836), .B2(KEYINPUT56), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n823), .A2(new_n824), .A3(new_n827), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n244), .A2(G952), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n830), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT118), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n830), .A2(new_n839), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(G51));
  NAND2_X1  g660(.A1(new_n832), .A2(new_n835), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n810), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n385), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n386), .A2(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n639), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n230), .B1(new_n832), .B2(new_n835), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(G469), .A3(new_n704), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n840), .B1(new_n853), .B2(new_n855), .ZN(G54));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n229), .ZN(new_n859));
  NAND3_X1  g673(.A1(KEYINPUT119), .A2(KEYINPUT58), .A3(G475), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n228), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n841), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT120), .ZN(G60));
  NAND2_X1  g680(.A1(G478), .A2(G902), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT59), .Z(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n810), .B2(new_n800), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n849), .A2(new_n569), .ZN(new_n870));
  OAI221_X1 g684(.A(new_n841), .B1(new_n869), .B2(new_n569), .C1(new_n870), .C2(new_n868), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(G63));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n873));
  NAND2_X1  g687(.A1(G217), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT60), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n832), .B2(new_n835), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n540), .B(KEYINPUT122), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n873), .B(new_n841), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n876), .A2(new_n591), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n841), .B1(new_n876), .B2(new_n878), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n884), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n886), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n882), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(G66));
  AOI21_X1  g705(.A(new_n244), .B1(new_n280), .B2(new_n421), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n756), .A2(new_n762), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(new_n244), .ZN(new_n894));
  INV_X1    g708(.A(G898), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n825), .B1(new_n895), .B2(G953), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n894), .B(new_n896), .ZN(G69));
  NAND2_X1  g711(.A1(new_n477), .A2(new_n479), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n222), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n602), .B2(G953), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n717), .A2(new_n711), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n685), .A2(new_n687), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n710), .A2(new_n451), .A3(new_n627), .A4(new_n679), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n804), .A2(new_n901), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(G953), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n244), .B1(G227), .B2(G900), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT124), .Z(new_n907));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n628), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n804), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT62), .Z(new_n912));
  NOR2_X1   g726(.A1(new_n674), .A2(new_n623), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n575), .A2(new_n581), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n516), .A2(new_n553), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n901), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n244), .A3(new_n899), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n905), .A2(new_n909), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n907), .A2(new_n908), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n918), .B(new_n919), .Z(G72));
  NAND2_X1  g734(.A1(G472), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT63), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n893), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n904), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n480), .A2(new_n481), .A3(new_n475), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT126), .Z(new_n927));
  OAI21_X1  g741(.A(new_n841), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n916), .A2(new_n893), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n610), .B1(new_n929), .B2(new_n922), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n781), .A2(new_n799), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n610), .A2(new_n922), .A3(new_n926), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n928), .A2(new_n930), .A3(new_n933), .ZN(G57));
endmodule


