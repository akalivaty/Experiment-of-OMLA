//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT91), .Z(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT13), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n206), .B1(new_n209), .B2(new_n205), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT89), .B1(new_n210), .B2(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT87), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G29gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n217), .A3(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n212), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n213), .B1(new_n220), .B2(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(new_n206), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT88), .B(G43gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G50gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n205), .A2(G43gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT86), .B1(new_n230), .B2(new_n206), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT86), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT15), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n213), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT87), .B(G29gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n212), .B1(new_n237), .B2(G36gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT14), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(new_n234), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G22gat), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n244), .A2(G1gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT16), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n246), .B2(G1gat), .ZN(new_n247));
  INV_X1    g046(.A(G8gat), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n248), .A2(KEYINPUT90), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(KEYINPUT90), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(KEYINPUT90), .A3(new_n248), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n243), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n241), .B1(new_n228), .B2(new_n234), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n253), .A3(new_n252), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n204), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n254), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n235), .A2(new_n259), .A3(new_n242), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n203), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT18), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n243), .A2(KEYINPUT17), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(new_n259), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n254), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT18), .A3(new_n203), .A4(new_n257), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G169gat), .B(G197gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G141gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT12), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n264), .A2(new_n275), .A3(new_n268), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G230gat), .ZN(new_n280));
  INV_X1    g079(.A(G233gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G99gat), .A2(G106gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT95), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT95), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(G99gat), .A3(G106gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT8), .ZN(new_n287));
  XNOR2_X1  g086(.A(G99gat), .B(G106gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G85gat), .A2(G92gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT96), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n295), .A2(new_n290), .A3(new_n291), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT96), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n288), .A4(new_n287), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n288), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT8), .ZN(new_n301));
  INV_X1    g100(.A(new_n290), .ZN(new_n302));
  INV_X1    g101(.A(new_n291), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n289), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT97), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(new_n287), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT97), .A3(new_n300), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G57gat), .B(G64gat), .Z(new_n311));
  NAND2_X1  g110(.A1(G71gat), .A2(G78gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT9), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT94), .ZN(new_n315));
  XNOR2_X1  g114(.A(G71gat), .B(G78gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n317), .A3(new_n313), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n311), .A2(new_n315), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n311), .A2(new_n318), .A3(new_n315), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(KEYINPUT92), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT92), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(G71gat), .A3(G78gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR3_X1   g124(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n321), .B(new_n323), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n319), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n299), .A3(new_n305), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT99), .B(KEYINPUT10), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n310), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT10), .A3(new_n330), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n282), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n282), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n329), .B2(new_n331), .ZN(new_n339));
  XNOR2_X1  g138(.A(G120gat), .B(G148gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n337), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n337), .B2(new_n339), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n279), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n265), .A2(new_n266), .A3(new_n310), .ZN(new_n349));
  AND2_X1   g148(.A1(G232gat), .A2(G233gat), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n335), .A2(new_n256), .B1(KEYINPUT41), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G134gat), .B(G162gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G190gat), .B(G218gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT98), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n350), .A2(KEYINPUT41), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  AND2_X1   g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n354), .A2(new_n358), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT21), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n328), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G127gat), .B(G155gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G231gat), .A2(G233gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(G183gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G211gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n366), .B(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n254), .B1(new_n363), .B2(new_n328), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n370), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n362), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT65), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n387), .B(new_n388), .C1(G183gat), .C2(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT27), .B(G183gat), .ZN(new_n391));
  INV_X1    g190(.A(G190gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n394), .A2(new_n395), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n378), .B(KEYINPUT26), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n398));
  AOI22_X1  g197(.A1(new_n383), .A2(new_n397), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n390), .A2(KEYINPUT25), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT64), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n389), .B(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n380), .B(new_n383), .C1(KEYINPUT66), .C2(KEYINPUT25), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n403), .C1(KEYINPUT66), .C2(new_n384), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n400), .B2(new_n404), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n409), .B2(new_n406), .ZN(new_n410));
  XOR2_X1   g209(.A(G211gat), .B(G218gat), .Z(new_n411));
  XOR2_X1   g210(.A(G197gat), .B(G204gat), .Z(new_n412));
  AOI21_X1  g211(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n411), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT70), .B(new_n417), .C1(new_n413), .C2(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n419), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n400), .B2(new_n404), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n407), .B(new_n421), .C1(new_n406), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT72), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  AOI21_X1  g227(.A(new_n377), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n424), .A2(new_n428), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G113gat), .ZN(new_n432));
  INV_X1    g231(.A(G120gat), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT1), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n432), .B2(new_n433), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT68), .ZN(new_n436));
  XNOR2_X1  g235(.A(G127gat), .B(G134gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT69), .B1(new_n405), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G227gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n281), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n405), .A2(new_n438), .ZN(new_n443));
  INV_X1    g242(.A(new_n438), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT69), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n400), .A2(new_n444), .A3(new_n404), .A4(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n439), .A2(new_n442), .A3(new_n443), .A4(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND3_X1  g249(.A1(new_n439), .A2(new_n443), .A3(new_n446), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n451), .A2(new_n441), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n447), .B(new_n450), .C1(new_n452), .C2(KEYINPUT33), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT34), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n447), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT33), .B1(new_n451), .B2(new_n441), .ZN(new_n457));
  INV_X1    g256(.A(new_n450), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n451), .A2(new_n441), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT32), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n453), .A2(new_n455), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n457), .A2(new_n456), .A3(new_n458), .ZN(new_n464));
  AOI211_X1 g263(.A(new_n441), .B(new_n451), .C1(KEYINPUT33), .C2(new_n450), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n460), .B2(KEYINPUT32), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n454), .B(KEYINPUT34), .C1(new_n451), .C2(new_n441), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G22gat), .B(G50gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G155gat), .ZN(new_n472));
  INV_X1    g271(.A(G162gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT2), .ZN(new_n475));
  NOR2_X1   g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G141gat), .B(G148gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n476), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n474), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n481), .B(new_n482), .C1(new_n478), .C2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT75), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n478), .A2(new_n483), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(KEYINPUT75), .A3(new_n481), .A4(new_n482), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n479), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n408), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n491), .A2(KEYINPUT79), .A3(new_n421), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT79), .B1(new_n491), .B2(new_n421), .ZN(new_n493));
  AND2_X1   g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n414), .A2(KEYINPUT78), .A3(new_n417), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n417), .B2(new_n414), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT78), .B1(new_n414), .B2(new_n417), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n490), .B1(new_n498), .B2(new_n408), .ZN(new_n499));
  INV_X1    g298(.A(new_n489), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(new_n493), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n491), .A2(new_n421), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n421), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n489), .B1(new_n506), .B2(new_n490), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n494), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n503), .B1(new_n502), .B2(new_n508), .ZN(new_n511));
  XOR2_X1   g310(.A(G78gat), .B(G106gat), .Z(new_n512));
  NOR3_X1   g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n508), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT31), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n514), .B1(new_n516), .B2(new_n509), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n471), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n509), .A3(new_n514), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n470), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n431), .B(new_n469), .C1(new_n518), .C2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n489), .A2(new_n444), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT4), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n489), .A2(new_n444), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT77), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(KEYINPUT77), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n500), .A2(KEYINPUT3), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n444), .B1(new_n489), .B2(new_n490), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT5), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n533), .A2(new_n534), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n524), .B2(new_n527), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT4), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n524), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n489), .B(new_n444), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n535), .A2(new_n538), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G1gat), .B(G29gat), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT0), .B(G57gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT6), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT80), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n542), .A2(new_n545), .ZN(new_n556));
  INV_X1    g355(.A(new_n532), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT77), .B1(new_n525), .B2(new_n528), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n539), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n538), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT80), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n553), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(KEYINPUT6), .A3(new_n551), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n523), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n522), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n518), .A2(new_n521), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT6), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n561), .B2(new_n551), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n546), .A2(new_n552), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n463), .A2(new_n468), .ZN(new_n572));
  INV_X1    g371(.A(new_n431), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n567), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT35), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n519), .A2(new_n520), .A3(new_n470), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n470), .B1(new_n519), .B2(new_n520), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n571), .A2(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n469), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT83), .ZN(new_n585));
  INV_X1    g384(.A(new_n424), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n585), .B(new_n428), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n420), .B2(new_n423), .ZN(new_n589));
  INV_X1    g388(.A(new_n428), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT83), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n587), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n590), .B(new_n594), .C1(new_n586), .C2(new_n587), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n407), .B1(new_n422), .B2(new_n406), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n419), .ZN(new_n598));
  OAI22_X1  g397(.A1(new_n598), .A2(KEYINPUT81), .B1(new_n419), .B2(new_n410), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT37), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n430), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n563), .A2(new_n595), .A3(new_n602), .A4(new_n564), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n552), .B1(new_n561), .B2(KEYINPUT80), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(KEYINPUT80), .B2(new_n561), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n559), .A2(new_n607), .A3(new_n537), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n608), .A2(new_n552), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n544), .A2(new_n537), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT39), .B(new_n610), .C1(new_n535), .C2(new_n536), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n606), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AND4_X1   g411(.A1(new_n606), .A2(new_n611), .A3(new_n608), .A4(new_n552), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n605), .B(new_n431), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n603), .A2(new_n614), .A3(new_n567), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n615), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n348), .B(new_n376), .C1(new_n576), .C2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n571), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g419(.A1(new_n617), .A2(new_n431), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT16), .B(G8gat), .Z(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT42), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT100), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT42), .B1(new_n621), .B2(new_n248), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n622), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(G1325gat));
  AOI21_X1  g427(.A(G15gat), .B1(new_n617), .B2(new_n572), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n581), .A2(new_n583), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(G15gat), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n617), .B2(new_n632), .ZN(G1326gat));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n579), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT101), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT43), .B(G22gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1327gat));
  AND3_X1   g436(.A1(new_n584), .A2(new_n615), .A3(KEYINPUT102), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT102), .B1(new_n584), .B2(new_n615), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n522), .A2(new_n565), .B1(new_n574), .B2(KEYINPUT35), .ZN(new_n640));
  OAI22_X1  g439(.A1(new_n638), .A2(new_n639), .B1(new_n640), .B2(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(KEYINPUT103), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n361), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n348), .A2(new_n375), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n362), .B1(new_n576), .B2(new_n616), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n237), .B1(new_n650), .B2(new_n571), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n648), .A2(new_n647), .ZN(new_n652));
  INV_X1    g451(.A(new_n237), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n618), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT45), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(G1328gat));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n647), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(G36gat), .A3(new_n573), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT104), .ZN(new_n661));
  OAI21_X1  g460(.A(G36gat), .B1(new_n650), .B2(new_n573), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(KEYINPUT104), .A3(new_n659), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .A4(new_n664), .ZN(G1329gat));
  NAND3_X1  g464(.A1(new_n652), .A2(new_n572), .A3(new_n223), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n630), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(new_n223), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(KEYINPUT47), .B(new_n666), .C1(new_n667), .C2(new_n223), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1330gat));
  NAND3_X1  g471(.A1(new_n652), .A2(new_n205), .A3(new_n579), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n650), .A2(new_n567), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(new_n205), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT48), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT48), .B(new_n673), .C1(new_n674), .C2(new_n205), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1331gat));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n576), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n681), .B(new_n642), .C1(new_n639), .C2(new_n638), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n262), .A2(new_n263), .ZN(new_n684));
  INV_X1    g483(.A(new_n258), .ZN(new_n685));
  AND4_X1   g484(.A1(new_n275), .A2(new_n684), .A3(new_n268), .A4(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n275), .B1(new_n264), .B2(new_n268), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n362), .A2(new_n688), .A3(new_n346), .A4(new_n375), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n618), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n431), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT49), .B(G64gat), .Z(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(G1333gat));
  NAND2_X1  g495(.A1(new_n690), .A2(new_n572), .ZN(new_n697));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n630), .A2(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n697), .A2(new_n698), .B1(new_n690), .B2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g500(.A1(new_n690), .A2(new_n579), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g502(.A1(new_n279), .A2(new_n375), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n346), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n646), .A2(new_n649), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G85gat), .B1(new_n707), .B2(new_n571), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n361), .B(new_n704), .C1(new_n641), .C2(new_n643), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n682), .A2(KEYINPUT51), .A3(new_n361), .A4(new_n704), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(new_n548), .A3(new_n618), .A4(new_n346), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n708), .A2(new_n714), .ZN(G1336gat));
  OAI21_X1  g514(.A(G92gat), .B1(new_n707), .B2(new_n573), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n573), .A2(G92gat), .A3(new_n347), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT105), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g520(.A(G99gat), .B1(new_n707), .B2(new_n630), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n469), .A2(G99gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n713), .A2(new_n346), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1338gat));
  NOR2_X1   g524(.A1(new_n567), .A2(G106gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n347), .B(new_n727), .C1(new_n711), .C2(new_n712), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT107), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n346), .A3(new_n726), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n646), .A2(new_n579), .A3(new_n649), .A4(new_n706), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT53), .B1(new_n733), .B2(G106gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(KEYINPUT106), .A3(G106gat), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n733), .B2(G106gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n736), .A2(new_n737), .A3(new_n728), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(G1339gat));
  AOI21_X1  g539(.A(new_n203), .B1(new_n267), .B2(new_n257), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n255), .A2(new_n257), .A3(new_n204), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n274), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n346), .A2(new_n278), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT97), .B1(new_n308), .B2(new_n300), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n306), .B(new_n288), .C1(new_n296), .C2(new_n287), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n330), .B1(new_n748), .B2(new_n299), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n311), .A2(new_n315), .A3(new_n318), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n325), .A2(new_n326), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n321), .A2(new_n323), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n319), .A3(new_n305), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n294), .B2(new_n298), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n749), .A2(new_n755), .A3(new_n332), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT10), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n310), .A2(new_n757), .A3(new_n328), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n338), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n334), .A2(new_n282), .A3(new_n336), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n342), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n337), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n764), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n343), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n761), .A2(new_n764), .A3(KEYINPUT108), .A4(KEYINPUT55), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n766), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n769), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n745), .B1(new_n775), .B2(new_n688), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n362), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n769), .A2(new_n774), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n772), .A2(new_n773), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n278), .A2(new_n743), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n778), .A2(new_n779), .A3(new_n361), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n375), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n361), .A2(new_n279), .A3(new_n346), .A4(new_n374), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n522), .A2(new_n618), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n432), .A3(new_n279), .ZN(new_n788));
  INV_X1    g587(.A(new_n786), .ZN(new_n789));
  OAI21_X1  g588(.A(G113gat), .B1(new_n789), .B2(new_n688), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1340gat));
  NAND2_X1  g590(.A1(new_n346), .A2(new_n433), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G120gat), .B1(new_n789), .B2(new_n347), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1341gat));
  NAND2_X1  g595(.A1(new_n786), .A2(new_n375), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT112), .B(G127gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1342gat));
  NAND2_X1  g598(.A1(new_n786), .A2(new_n361), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(G134gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT56), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(G134gat), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n804), .B(new_n805), .C1(KEYINPUT56), .C2(new_n801), .ZN(G1343gat));
  NOR3_X1   g605(.A1(new_n631), .A2(new_n571), .A3(new_n431), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n784), .A2(new_n579), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n781), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n765), .B2(new_n766), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n765), .A2(new_n814), .A3(new_n766), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n279), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n772), .A2(new_n773), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n745), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n362), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n813), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(KEYINPUT116), .A3(new_n362), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n375), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT57), .B(new_n579), .C1(new_n825), .C2(new_n783), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n808), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n279), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n809), .A2(new_n808), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n688), .A2(G141gat), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n828), .A2(G141gat), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g631(.A(G148gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n833), .A3(new_n346), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  AOI211_X1 g634(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n761), .C2(new_n764), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n688), .A2(new_n815), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n744), .B1(new_n837), .B2(new_n779), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n781), .B1(new_n838), .B2(new_n361), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n783), .B1(new_n839), .B2(new_n374), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT117), .B(new_n835), .C1(new_n840), .C2(new_n567), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n579), .B(new_n810), .C1(new_n782), .C2(new_n783), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n375), .B1(new_n821), .B2(new_n781), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n579), .B1(new_n844), .B2(new_n783), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT117), .B1(new_n845), .B2(new_n835), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n346), .B(new_n807), .C1(new_n843), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G148gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n812), .A2(new_n826), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n346), .A3(new_n807), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n833), .A2(KEYINPUT59), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT118), .B1(new_n848), .B2(KEYINPUT59), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n834), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT119), .B(new_n834), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1345gat));
  AOI21_X1  g659(.A(G155gat), .B1(new_n829), .B2(new_n375), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n374), .A2(new_n472), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n827), .B2(new_n862), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n829), .B2(new_n361), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n362), .A2(new_n473), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n827), .B2(new_n865), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n579), .A2(new_n469), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n431), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n784), .A2(new_n571), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n688), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n784), .A2(new_n571), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n688), .A2(G169gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(G1348gat));
  INV_X1    g677(.A(G176gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n870), .A2(new_n879), .A3(new_n347), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n346), .A3(new_n869), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n879), .ZN(G1349gat));
  NOR2_X1   g681(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n875), .A2(new_n391), .A3(new_n375), .A4(new_n869), .ZN(new_n884));
  OAI21_X1  g683(.A(G183gat), .B1(new_n870), .B2(new_n374), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT122), .Z(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n886), .B(new_n889), .ZN(G1350gat));
  NOR2_X1   g689(.A1(new_n362), .A2(G190gat), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n869), .B(new_n891), .C1(new_n873), .C2(new_n874), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G190gat), .B1(new_n870), .B2(new_n362), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT61), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT124), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1351gat));
  INV_X1    g700(.A(new_n843), .ZN(new_n902));
  INV_X1    g701(.A(new_n846), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n630), .A2(new_n431), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n571), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n688), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n905), .A2(new_n567), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n875), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n873), .B2(new_n874), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT125), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n688), .A2(G197gat), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n910), .B(new_n911), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n914), .B2(new_n916), .ZN(new_n920));
  INV_X1    g719(.A(new_n910), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT126), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(G1352gat));
  OR2_X1    g722(.A1(new_n347), .A2(G204gat), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n915), .A2(KEYINPUT62), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n346), .A3(new_n908), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G204gat), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT62), .B1(new_n915), .B2(new_n924), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(G1353gat));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n916), .ZN(new_n930));
  INV_X1    g729(.A(G211gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n375), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n904), .A2(new_n375), .A3(new_n908), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(KEYINPUT63), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  INV_X1    g738(.A(G218gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n909), .A2(new_n940), .A3(new_n362), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n930), .A2(new_n361), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n940), .ZN(G1355gat));
endmodule


