//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT79), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n204), .B(new_n206), .Z(new_n207));
  XOR2_X1   g006(.A(G155gat), .B(G162gat), .Z(new_n208));
  XNOR2_X1  g007(.A(G141gat), .B(G148gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(KEYINPUT2), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G141gat), .B(G148gat), .Z(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT2), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G204gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G197gat), .ZN(new_n219));
  INV_X1    g018(.A(G197gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G204gat), .ZN(new_n221));
  INV_X1    g020(.A(G211gat), .ZN(new_n222));
  INV_X1    g021(.A(G218gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n219), .B(new_n221), .C1(new_n224), .C2(KEYINPUT22), .ZN(new_n225));
  XOR2_X1   g024(.A(G211gat), .B(G218gat), .Z(new_n226));
  OR2_X1    g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT29), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n217), .B1(new_n229), .B2(KEYINPUT3), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n210), .A2(new_n216), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n227), .A2(new_n228), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n230), .A2(KEYINPUT80), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n239), .B(new_n217), .C1(new_n229), .C2(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n229), .A2(new_n244), .ZN(new_n245));
  AOI211_X1 g044(.A(KEYINPUT81), .B(KEYINPUT29), .C1(new_n227), .C2(new_n228), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n232), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n217), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n236), .B(KEYINPUT71), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n242), .B1(new_n249), .B2(new_n235), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n207), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n241), .A2(new_n242), .B1(new_n248), .B2(new_n250), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n255), .A2(KEYINPUT82), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n255), .B2(KEYINPUT82), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(G22gat), .B1(new_n252), .B2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(new_n207), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n255), .B2(KEYINPUT82), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(KEYINPUT82), .A3(new_n256), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n269), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n272), .A4(new_n271), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n274), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G183gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT27), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT28), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT67), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n294), .B2(KEYINPUT28), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n281), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT23), .B1(new_n278), .B2(KEYINPUT64), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n299), .B(new_n300), .C1(G169gat), .C2(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n301), .A3(new_n272), .ZN(new_n302));
  AND3_X1   g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n297), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(KEYINPUT65), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n316), .C1(new_n308), .C2(new_n291), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n298), .A2(KEYINPUT25), .A3(new_n301), .A4(new_n272), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n307), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n296), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n291), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n289), .ZN(new_n326));
  INV_X1    g125(.A(new_n319), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT66), .B1(new_n282), .B2(new_n286), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(new_n303), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(new_n314), .A3(new_n311), .A4(new_n312), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n326), .A2(new_n281), .B1(new_n331), .B2(new_n307), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n322), .B(KEYINPUT72), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n321), .A2(new_n323), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n267), .B1(new_n335), .B2(new_n237), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n322), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n296), .B2(new_n320), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT73), .A4(new_n236), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G8gat), .B(G36gat), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT75), .ZN(new_n343));
  XOR2_X1   g142(.A(G64gat), .B(G92gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n236), .B(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n334), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n296), .A2(new_n320), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n323), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n341), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  AOI211_X1 g156(.A(new_n345), .B(new_n352), .C1(new_n336), .C2(new_n340), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT30), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(KEYINPUT77), .A3(new_n355), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n341), .B2(new_n353), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT74), .B(new_n352), .C1(new_n336), .C2(new_n340), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n366), .B2(new_n345), .ZN(new_n367));
  NOR4_X1   g166(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT76), .A4(new_n346), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(KEYINPUT1), .ZN(new_n371));
  XOR2_X1   g170(.A(G127gat), .B(G134gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n231), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR3_X1    g175(.A1(new_n372), .A2(KEYINPUT1), .A3(new_n370), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(KEYINPUT1), .B2(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n233), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n376), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n217), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n374), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n381), .A3(new_n383), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT39), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n389), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n399), .A2(new_n389), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT39), .B1(new_n388), .B2(new_n389), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n401), .B(new_n396), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT40), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n405), .B2(new_n404), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n266), .B1(new_n369), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n396), .B1(new_n386), .B2(new_n391), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n398), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n392), .A2(KEYINPUT6), .A3(new_n397), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT87), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n414), .A3(KEYINPUT6), .A4(new_n397), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n411), .A2(new_n413), .A3(new_n415), .A4(new_n354), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n349), .A2(new_n351), .A3(new_n348), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n236), .B1(new_n337), .B2(new_n339), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n350), .A2(new_n234), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n338), .B1(new_n421), .B2(new_n322), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n236), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT84), .B(KEYINPUT37), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n352), .B1(new_n336), .B2(new_n340), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT37), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n346), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT83), .B1(new_n422), .B2(new_n236), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n418), .A2(new_n419), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n417), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT84), .B1(new_n434), .B2(KEYINPUT37), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT86), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(KEYINPUT37), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  INV_X1    g239(.A(new_n430), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n425), .B2(new_n426), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n424), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n416), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT73), .B1(new_n422), .B2(new_n236), .ZN(new_n445));
  INV_X1    g244(.A(new_n340), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n353), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT74), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n363), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT37), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n346), .B1(new_n425), .B2(new_n426), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT88), .B1(new_n452), .B2(new_n429), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n454), .B(new_n428), .C1(new_n450), .C2(new_n451), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n444), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n408), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT32), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT70), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n350), .B2(new_n379), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n350), .A2(new_n379), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n350), .A2(new_n459), .A3(new_n379), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n458), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT33), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n462), .A2(new_n465), .A3(new_n463), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n332), .A2(KEYINPUT70), .A3(new_n373), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n461), .B2(new_n460), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT32), .B1(new_n478), .B2(new_n465), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n478), .B2(new_n465), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n481), .A3(new_n471), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n476), .B1(new_n473), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT36), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n482), .ZN(new_n486));
  INV_X1    g285(.A(new_n476), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n411), .A2(new_n412), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n361), .B(new_n493), .C1(new_n367), .C2(new_n368), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n494), .B2(new_n266), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n457), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n369), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n265), .A2(new_n488), .A3(new_n490), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n411), .A2(new_n415), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT35), .B1(new_n499), .B2(new_n413), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n483), .A2(new_n484), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n265), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT35), .B1(new_n494), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G183gat), .B(G211gat), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G78gat), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT97), .ZN(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(KEYINPUT97), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n513), .A2(new_n509), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT21), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G231gat), .A2(G233gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n517), .B(new_n518), .Z(new_n519));
  XNOR2_X1  g318(.A(G127gat), .B(G155gat), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n508), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n525), .A3(new_n507), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  AOI21_X1  g331(.A(G1gat), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n531), .B(new_n534), .C1(new_n532), .C2(G1gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G8gat), .ZN(new_n539));
  INV_X1    g338(.A(G8gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n515), .A2(new_n516), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT98), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n544), .B2(KEYINPUT21), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT99), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n528), .A2(new_n530), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n528), .B2(new_n530), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G134gat), .B(G162gat), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT41), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555));
  NOR2_X1   g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT14), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(KEYINPUT14), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT91), .B(G36gat), .ZN(new_n559));
  INV_X1    g358(.A(G29gat), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G43gat), .B(G50gat), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT90), .ZN(new_n563));
  XNOR2_X1  g362(.A(G43gat), .B(G50gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n561), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n563), .B2(new_n566), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT92), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT92), .B1(new_n569), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n555), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT17), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT100), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT7), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n580), .B2(KEYINPUT101), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n590), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n579), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n574), .ZN(new_n598));
  INV_X1    g397(.A(new_n594), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n598), .A2(new_n599), .B1(KEYINPUT41), .B2(new_n553), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n595), .B2(new_n600), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n554), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  INV_X1    g406(.A(new_n554), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n603), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n552), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n552), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n550), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G169gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT89), .B(G197gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  INV_X1    g420(.A(new_n579), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n598), .B2(new_n555), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n542), .B(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n623), .A2(new_n625), .B1(new_n542), .B2(new_n598), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT95), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT18), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n577), .A2(new_n625), .A3(new_n579), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n598), .A2(new_n542), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n632), .A2(KEYINPUT18), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT96), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n630), .A3(new_n633), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n598), .B(new_n542), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n629), .B(KEYINPUT13), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n621), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n636), .A2(new_n641), .A3(new_n621), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G230gat), .ZN(new_n650));
  INV_X1    g449(.A(G233gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n594), .A2(new_n515), .A3(new_n516), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n592), .A2(new_n543), .A3(new_n593), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT102), .B(KEYINPUT10), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n544), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n652), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n652), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n649), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n544), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n663));
  INV_X1    g462(.A(new_n656), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n653), .B2(new_n654), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n649), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n666), .B(new_n667), .C1(new_n655), .C2(new_n660), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n615), .A2(new_n646), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n506), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n493), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT103), .B(G1gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1324gat));
  NOR2_X1   g473(.A1(new_n671), .A2(new_n497), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n676), .A2(KEYINPUT105), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n676), .A2(KEYINPUT105), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n680), .A2(new_n681), .B1(G8gat), .B2(new_n678), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(KEYINPUT42), .A3(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n502), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n671), .A2(G15gat), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n492), .A2(KEYINPUT106), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n492), .A2(KEYINPUT106), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n671), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(G1326gat));
  NAND3_X1  g490(.A1(new_n506), .A2(new_n266), .A3(new_n670), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT108), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  NOR3_X1   g497(.A1(new_n550), .A2(new_n646), .A3(new_n669), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n457), .A2(new_n495), .B1(new_n501), .B2(new_n504), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n614), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT109), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n705), .B(KEYINPUT44), .C1(new_n701), .C2(new_n614), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n506), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n701), .A2(KEYINPUT110), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n703), .A3(new_n613), .A4(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n700), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n493), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n494), .A2(new_n266), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n485), .A2(new_n491), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n456), .B2(new_n408), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n501), .A2(new_n504), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n613), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n700), .ZN(new_n721));
  INV_X1    g520(.A(new_n493), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n560), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n724), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n369), .A3(new_n559), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT111), .Z(new_n728));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n497), .ZN(new_n729));
  OAI221_X1 g528(.A(new_n728), .B1(KEYINPUT46), .B2(new_n726), .C1(new_n559), .C2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n705), .B1(new_n720), .B2(KEYINPUT44), .ZN(new_n732));
  INV_X1    g531(.A(new_n706), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n711), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n492), .A3(new_n699), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n685), .A2(G43gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n702), .A2(new_n699), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT112), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n731), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT112), .B1(new_n721), .B2(new_n737), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n731), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n689), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n712), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT113), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n745), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n689), .B(new_n700), .C1(new_n707), .C2(new_n711), .ZN(new_n751));
  INV_X1    g550(.A(G43gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n739), .B1(new_n735), .B2(G43gat), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n753), .B(new_n754), .C1(new_n731), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n749), .A2(new_n756), .ZN(G1330gat));
  AOI21_X1  g556(.A(new_n203), .B1(new_n712), .B2(new_n266), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n720), .A2(G50gat), .A3(new_n265), .A4(new_n700), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n760), .B(new_n763), .ZN(G1331gat));
  INV_X1    g563(.A(new_n669), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n615), .A2(new_n645), .A3(new_n765), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n709), .A2(new_n710), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n722), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g568(.A(new_n497), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n771), .B(new_n772), .Z(G1333gat));
  AOI21_X1  g572(.A(G71gat), .B1(new_n767), .B2(new_n502), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n746), .A2(G71gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n767), .A2(new_n266), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n550), .A2(new_n645), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n702), .A2(KEYINPUT51), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT51), .B1(new_n702), .B2(new_n781), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n669), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n586), .A3(new_n722), .ZN(new_n786));
  INV_X1    g585(.A(new_n734), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n669), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n787), .A2(new_n493), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  NOR4_X1   g592(.A1(new_n787), .A2(new_n587), .A3(new_n497), .A4(new_n788), .ZN(new_n794));
  AOI21_X1  g593(.A(G92gat), .B1(new_n785), .B2(new_n369), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1337gat));
  AOI21_X1  g598(.A(G99gat), .B1(new_n785), .B2(new_n502), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n787), .A2(new_n788), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n746), .A2(G99gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(G1338gat));
  INV_X1    g602(.A(G106gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n784), .B2(new_n265), .ZN(new_n805));
  INV_X1    g604(.A(new_n788), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n734), .A2(G106gat), .A3(new_n266), .A4(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n810), .B(new_n811), .Z(G1339gat));
  NAND3_X1  g611(.A1(new_n657), .A2(new_n658), .A3(new_n652), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n666), .A3(KEYINPUT54), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n659), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n814), .A2(new_n816), .A3(KEYINPUT55), .A4(new_n649), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n668), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n667), .B1(new_n659), .B2(new_n815), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n819), .B2(new_n814), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n636), .A2(new_n641), .A3(new_n621), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n642), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n626), .A2(new_n630), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n639), .A2(new_n640), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n620), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n644), .A2(new_n669), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n613), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n612), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n821), .B1(new_n829), .B2(new_n610), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n644), .A2(new_n826), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n549), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n550), .A2(new_n614), .A3(new_n646), .A4(new_n765), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n722), .A3(new_n498), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n497), .ZN(new_n839));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n645), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n497), .A2(new_n722), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n835), .B2(new_n265), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT118), .B(new_n266), .C1(new_n833), .C2(new_n834), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n685), .B(new_n841), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n645), .A2(G113gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  AOI21_X1  g648(.A(G120gat), .B1(new_n839), .B2(new_n669), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n669), .A2(G120gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n847), .B2(new_n851), .ZN(G1341gat));
  NAND3_X1  g651(.A1(new_n847), .A2(G127gat), .A3(new_n550), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n838), .A2(new_n497), .A3(new_n550), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(G127gat), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(G1342gat));
  NAND2_X1  g656(.A1(new_n847), .A2(new_n613), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G134gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n497), .A2(new_n613), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(G134gat), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n838), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n838), .A2(KEYINPUT56), .A3(new_n861), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G1343gat));
  AND2_X1   g663(.A1(new_n820), .A2(KEYINPUT121), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n820), .A2(KEYINPUT121), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n865), .A2(new_n866), .A3(new_n818), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n645), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n613), .B1(new_n868), .B2(new_n827), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n549), .B1(new_n869), .B2(new_n832), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n834), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n265), .ZN(new_n873));
  INV_X1    g672(.A(new_n835), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n265), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n841), .A2(new_n492), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n645), .A2(G141gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n689), .A2(new_n266), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n874), .A2(new_n493), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n497), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n646), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n879), .A2(new_n880), .B1(new_n885), .B2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1344gat));
  NOR2_X1   g687(.A1(new_n879), .A2(new_n765), .ZN(new_n889));
  INV_X1    g688(.A(G148gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n889), .A2(KEYINPUT59), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n871), .B2(new_n266), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n874), .A2(new_n876), .A3(new_n265), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n669), .A3(new_n878), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n669), .A2(new_n890), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n891), .A2(new_n897), .B1(new_n884), .B2(new_n898), .ZN(G1345gat));
  OAI21_X1  g698(.A(G155gat), .B1(new_n879), .B2(new_n549), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n550), .A2(new_n213), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n884), .B2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n879), .B2(new_n614), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n860), .A2(G162gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n883), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1347gat));
  NOR4_X1   g705(.A1(new_n874), .A2(new_n722), .A3(new_n497), .A4(new_n503), .ZN(new_n907));
  AOI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n645), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n497), .A2(new_n722), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n502), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n843), .B2(new_n845), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT124), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n914), .B(new_n911), .C1(new_n843), .C2(new_n845), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n645), .A2(G169gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  INV_X1    g717(.A(G176gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n907), .A2(new_n919), .A3(new_n669), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(new_n669), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(G1349gat));
  AND3_X1   g721(.A1(new_n907), .A2(new_n293), .A3(new_n550), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n913), .A2(new_n550), .A3(new_n915), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(G183gat), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n925), .B(new_n927), .ZN(G1350gat));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n613), .A3(new_n915), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(G190gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n930), .B2(G190gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(G190gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT126), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n931), .A3(G190gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(KEYINPUT61), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n907), .A2(new_n286), .A3(new_n613), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(G1351gat));
  NAND2_X1  g739(.A1(new_n689), .A2(new_n909), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n895), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n220), .A3(new_n646), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n875), .A2(new_n942), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n645), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n944), .A2(new_n947), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n945), .A2(G204gat), .A3(new_n765), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n895), .A2(new_n669), .A3(new_n942), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n953), .B(new_n955), .C1(new_n950), .C2(new_n949), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n946), .A2(new_n222), .A3(new_n550), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n895), .A2(new_n550), .A3(new_n942), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n943), .B2(new_n614), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n223), .A3(new_n613), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


