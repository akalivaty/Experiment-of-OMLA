//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1155,
    new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT65), .Z(new_n462));
  INV_X1    g037(.A(G2106), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(new_n455), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(KEYINPUT67), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G137), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n478), .A2(new_n483), .ZN(G160));
  AOI21_X1  g059(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  AOI22_X1  g060(.A1(G124), .A2(new_n485), .B1(new_n479), .B2(G136), .ZN(new_n486));
  INV_X1    g061(.A(G100), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n487), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT68), .B1(new_n487), .B2(new_n466), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G112), .B2(new_n466), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT69), .Z(G162));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n469), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n470), .A2(new_n475), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n512), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n510), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND3_X1  g097(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n518), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n516), .A2(new_n517), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT70), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n512), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n527), .B1(new_n534), .B2(G51), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n515), .A2(new_n514), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n518), .ZN(new_n540));
  AOI22_X1  g115(.A1(G651), .A2(new_n539), .B1(new_n540), .B2(G90), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n531), .A2(new_n533), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n534), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n537), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(G651), .A2(new_n549), .B1(new_n540), .B2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT71), .Z(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n537), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n540), .A2(G91), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n530), .B2(G53), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  OR2_X1    g145(.A1(new_n507), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n530), .B2(G49), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n540), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n507), .A2(new_n511), .A3(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT72), .ZN(new_n576));
  OAI211_X1 g151(.A(G48), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n505), .B2(new_n506), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n507), .A2(new_n511), .A3(new_n583), .A4(G86), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n576), .A2(new_n577), .A3(new_n582), .A4(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n537), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(G651), .A2(new_n588), .B1(new_n540), .B2(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n542), .B2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n537), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n593), .A2(new_n596), .B1(G651), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT73), .ZN(new_n602));
  OAI21_X1  g177(.A(G54), .B1(new_n534), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n592), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n592), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g192(.A1(new_n470), .A2(new_n475), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n481), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n479), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n485), .A2(G123), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n624), .A3(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n635), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT75), .Z(new_n649));
  NOR2_X1   g224(.A1(G2072), .A2(G2078), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n444), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n647), .B(new_n648), .C1(new_n444), .C2(new_n650), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n649), .A3(new_n647), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT76), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT20), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n669), .A2(new_n666), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT77), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n669), .A3(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT78), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G22), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G166), .B2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(G1971), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n681), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT81), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT32), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n692), .A2(KEYINPUT34), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT34), .B1(new_n692), .B2(new_n695), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n681), .A2(G24), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G290), .B2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n479), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n485), .A2(G119), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n466), .A2(G107), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n704), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT79), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n703), .B2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n696), .A2(new_n697), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT36), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n710), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n710), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT29), .ZN(new_n723));
  INV_X1    g298(.A(G2090), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n618), .A2(G127), .ZN(new_n726));
  INV_X1    g301(.A(G115), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n472), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n466), .B1(new_n728), .B2(KEYINPUT86), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT86), .B2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n731));
  NAND2_X1  g306(.A1(G103), .A2(G2104), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n479), .A2(G139), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n710), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n710), .B2(G33), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(new_n442), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n681), .A2(G4), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n605), .B2(new_n681), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT82), .B(G1348), .Z(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT83), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n725), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G171), .A2(new_n681), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G5), .B2(new_n681), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(G1961), .ZN(new_n748));
  NAND2_X1  g323(.A1(G164), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G27), .B2(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(new_n443), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n443), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n747), .A2(G1961), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n748), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n710), .A2(G32), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n481), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n485), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT26), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT87), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(KEYINPUT87), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(new_n710), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n681), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(G1956), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G11), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT30), .B(G28), .Z(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G29), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n629), .A2(new_n710), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n681), .A2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G168), .B2(new_n681), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n779), .B1(new_n781), .B2(G1966), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n767), .A2(new_n772), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n552), .B2(G16), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G1966), .B2(new_n781), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n754), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n737), .A2(new_n442), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n710), .A2(G26), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT28), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n479), .A2(G140), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT84), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n485), .A2(G128), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n466), .A2(G116), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT85), .B(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n710), .B1(new_n801), .B2(G34), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n801), .B2(G34), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G160), .B2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G2084), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n788), .A2(new_n789), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n720), .A2(new_n744), .A3(new_n807), .ZN(G311));
  INV_X1    g383(.A(G311), .ZN(G150));
  NAND2_X1  g384(.A1(new_n605), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT38), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  INV_X1    g387(.A(G67), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n537), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n509), .B1(new_n814), .B2(KEYINPUT90), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(KEYINPUT90), .B2(new_n814), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT91), .B(G93), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n534), .A2(G55), .B1(new_n540), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n552), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n816), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(new_n551), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n811), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(G860), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n820), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT92), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(G145));
  NAND2_X1  g405(.A1(new_n730), .A2(new_n735), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n797), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n479), .A2(G142), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT93), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n485), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n466), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n708), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n832), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n501), .A2(new_n503), .ZN(new_n841));
  INV_X1    g416(.A(new_n498), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n763), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n621), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(G160), .B(new_n629), .Z(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G162), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  INV_X1    g427(.A(new_n850), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n846), .A2(new_n853), .A3(new_n847), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g431(.A1(new_n820), .A2(new_n608), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT96), .ZN(new_n858));
  XOR2_X1   g433(.A(G290), .B(G305), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n687), .B(G303), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n859), .B(new_n860), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n859), .B(new_n860), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(KEYINPUT95), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT95), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n614), .B(new_n822), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n601), .A2(new_n603), .ZN(new_n870));
  NAND2_X1  g445(.A1(G299), .A2(KEYINPUT94), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n564), .B(new_n872), .C1(new_n566), .C2(new_n568), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n870), .A2(new_n600), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n604), .A2(KEYINPUT94), .A3(G299), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(KEYINPUT41), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n869), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n868), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n869), .A2(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n869), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n866), .B(KEYINPUT95), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n867), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n858), .B1(new_n885), .B2(G868), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n884), .A2(KEYINPUT96), .A3(new_n608), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(G295));
  NOR2_X1   g463(.A1(new_n886), .A2(new_n887), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n890));
  INV_X1    g465(.A(new_n876), .ZN(new_n891));
  AOI21_X1  g466(.A(G301), .B1(new_n819), .B2(new_n821), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n819), .A2(G301), .A3(new_n821), .ZN(new_n894));
  AOI21_X1  g469(.A(G168), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n896), .A2(new_n892), .A3(G286), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n891), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n899));
  OAI21_X1  g474(.A(G286), .B1(new_n896), .B2(new_n892), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n893), .A2(G168), .A3(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n876), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT98), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(KEYINPUT98), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(new_n861), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n904), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n908), .B2(new_n861), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n904), .A2(KEYINPUT98), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n863), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n861), .B1(new_n905), .B2(new_n906), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT97), .B(KEYINPUT43), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n852), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n890), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n917), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n907), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n916), .A3(new_n852), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n909), .A2(new_n921), .B1(new_n922), .B2(new_n920), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n919), .B1(new_n923), .B2(new_n890), .ZN(G397));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n797), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n764), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n763), .A2(G1996), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G40), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n478), .A2(new_n931), .A3(new_n483), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(G164), .B2(G1384), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI211_X1 g510(.A(new_n715), .B(new_n708), .C1(new_n930), .C2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n797), .A2(G2067), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n936), .A2(KEYINPUT125), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT125), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n938), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n935), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n941), .A2(G1986), .A3(G290), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT48), .Z(new_n943));
  XNOR2_X1  g518(.A(new_n708), .B(new_n715), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n935), .B1(new_n930), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n935), .A2(new_n927), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT46), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n926), .A2(new_n764), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n941), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n950), .B(new_n951), .Z(new_n952));
  INV_X1    g527(.A(KEYINPUT127), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n940), .B(new_n954), .C1(new_n953), .C2(new_n952), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT102), .B(G8), .Z(new_n957));
  NOR3_X1   g532(.A1(new_n478), .A2(new_n931), .A3(new_n483), .ZN(new_n958));
  NOR2_X1   g533(.A1(G164), .A2(G1384), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n962));
  INV_X1    g537(.A(G86), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n577), .B1(new_n518), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(G61), .B1(new_n515), .B2(new_n514), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n509), .B1(new_n965), .B2(new_n580), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n962), .B(G1981), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G305), .B2(G1981), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n582), .A2(new_n575), .A3(new_n577), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n962), .B1(new_n969), .B2(G1981), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n961), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n582), .A2(new_n584), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n576), .A4(new_n577), .ZN(new_n974));
  OAI21_X1  g549(.A(G1981), .B1(new_n964), .B2(new_n966), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT104), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT49), .A4(new_n967), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(new_n977), .A3(new_n960), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n971), .A2(new_n977), .A3(KEYINPUT105), .A4(new_n960), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(G288), .A2(G1976), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT107), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n974), .B(KEYINPUT106), .Z(new_n986));
  OAI21_X1  g561(.A(new_n960), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G303), .A2(G8), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT100), .B(KEYINPUT55), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n988), .B(new_n989), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT101), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n958), .A3(new_n934), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n684), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n843), .A2(new_n996), .A3(new_n992), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n958), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n995), .B1(G2090), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n988), .B(new_n989), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT101), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n991), .A2(G8), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n958), .A2(new_n959), .ZN(new_n1005));
  INV_X1    g580(.A(new_n957), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n572), .A2(G1976), .A3(new_n573), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(KEYINPUT103), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1008), .A2(new_n1011), .B1(G288), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n960), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n982), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1004), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n987), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n982), .A2(KEYINPUT110), .A3(new_n1015), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT110), .B1(new_n982), .B2(new_n1015), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1004), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n999), .A2(KEYINPUT108), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n997), .A2(new_n958), .A3(new_n998), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n724), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n957), .B1(new_n1026), .B2(new_n995), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT109), .B1(new_n1027), .B2(new_n1001), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n1029));
  AOI21_X1  g604(.A(G2090), .B1(new_n999), .B2(KEYINPUT108), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1030), .A2(new_n1025), .B1(new_n684), .B2(new_n994), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1029), .B(new_n990), .C1(new_n1031), .C2(new_n957), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1022), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1966), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n994), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n997), .A2(new_n958), .A3(new_n998), .A4(new_n805), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n957), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1038), .A2(G168), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT63), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1004), .A2(KEYINPUT63), .A3(new_n1039), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1001), .B1(new_n1000), .B2(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1043), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1045), .A2(KEYINPUT111), .A3(new_n982), .A4(new_n1015), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1041), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n956), .B(new_n1019), .C1(new_n1040), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1016), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n982), .A2(KEYINPUT110), .A3(new_n1015), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1039), .A3(new_n1053), .A4(new_n1004), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1047), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT112), .B1(new_n1056), .B2(new_n1018), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G168), .A2(new_n957), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT119), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT51), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1038), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT120), .B(new_n957), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1060), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1068), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT62), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n993), .A2(new_n958), .A3(new_n934), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n443), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT123), .B(G1961), .Z(new_n1082));
  AOI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n999), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1073), .A2(new_n1078), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n566), .B2(new_n568), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n530), .A2(new_n565), .A3(G53), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(KEYINPUT114), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(new_n564), .A3(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n1097));
  AND3_X1   g672(.A1(new_n1096), .A2(KEYINPUT115), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT115), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1098), .A2(new_n1099), .B1(new_n1100), .B2(G299), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  INV_X1    g677(.A(G1956), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1079), .A2(new_n1102), .B1(new_n999), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1090), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n999), .A2(new_n741), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n958), .A2(new_n925), .A3(new_n959), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n605), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n604), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT60), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1101), .A2(new_n1090), .A3(new_n1104), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1079), .A2(new_n927), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1005), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n551), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1104), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n1128));
  OAI221_X1 g703(.A(new_n1128), .B1(new_n1100), .B2(G299), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1112), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1106), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1115), .A2(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n993), .A2(new_n934), .A3(new_n1084), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n958), .B(KEYINPUT124), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1083), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1087), .B1(G171), .B2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1136), .B2(G171), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1083), .A2(G301), .A3(new_n1085), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1137), .A2(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1133), .B(new_n1142), .C1(new_n1072), .C2(new_n1071), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1089), .A2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1048), .A2(new_n1057), .B1(new_n1144), .B2(new_n1034), .ZN(new_n1145));
  AND2_X1   g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n942), .B1(new_n935), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT99), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n945), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n955), .B1(new_n1145), .B2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g725(.A1(G229), .A2(new_n464), .A3(G401), .A4(G227), .ZN(new_n1152));
  NAND2_X1  g726(.A1(new_n855), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n923), .A2(new_n1153), .ZN(G308));
  AND2_X1   g728(.A1(new_n922), .A2(new_n920), .ZN(new_n1155));
  NOR3_X1   g729(.A1(new_n907), .A2(new_n910), .A3(new_n920), .ZN(new_n1156));
  OAI211_X1 g730(.A(new_n855), .B(new_n1152), .C1(new_n1155), .C2(new_n1156), .ZN(G225));
endmodule


