//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G134), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n199), .A3(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT67), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n208), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n208), .A2(G143), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G128), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n212), .B(new_n218), .C1(new_n220), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G143), .B(G146), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n219), .A3(G128), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n228), .A2(KEYINPUT68), .A3(new_n212), .A4(new_n218), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n202), .A2(new_n230), .A3(new_n204), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n206), .A2(new_n226), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT66), .B(G116), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G119), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT2), .B(G113), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n242), .A3(G119), .ZN(new_n243));
  INV_X1    g057(.A(new_n234), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n237), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n227), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n250), .B(new_n251), .C1(new_n209), .C2(new_n211), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n200), .A2(KEYINPUT64), .A3(G131), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT64), .A2(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n196), .A2(new_n198), .A3(new_n256), .A4(new_n199), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n232), .A2(new_n248), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n205), .A2(new_n224), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n232), .A2(new_n259), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(KEYINPUT30), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n193), .B(new_n260), .C1(new_n265), .C2(new_n248), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n262), .B1(new_n232), .B2(new_n259), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n247), .B1(new_n268), .B2(new_n263), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n193), .A4(new_n260), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n193), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n260), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n260), .A2(KEYINPUT71), .A3(new_n274), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n261), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n247), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n260), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n277), .B(new_n278), .C1(KEYINPUT70), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n273), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n188), .B1(new_n272), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n232), .A2(new_n248), .A3(new_n259), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n248), .B1(new_n232), .B2(new_n259), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n277), .A3(new_n278), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n273), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n260), .A2(KEYINPUT71), .A3(new_n274), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT71), .B1(new_n260), .B2(new_n274), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n260), .A2(new_n281), .ZN(new_n296));
  INV_X1    g110(.A(new_n279), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n295), .A2(new_n300), .A3(new_n301), .A4(new_n284), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n292), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n269), .A2(new_n260), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(new_n193), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n305), .B2(new_n301), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(KEYINPUT32), .A2(new_n287), .B1(new_n307), .B2(G472), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n287), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT70), .B1(new_n296), .B2(new_n297), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(new_n294), .A3(new_n293), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n193), .B1(new_n313), .B2(new_n284), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n267), .A2(new_n271), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n187), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n310), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT73), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n308), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G217), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(G234), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT75), .B1(new_n324), .B2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(G128), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT75), .B(new_n328), .C1(new_n324), .C2(G128), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G110), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT24), .B(G110), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT74), .B1(new_n324), .B2(G128), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n207), .A3(G119), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n335), .A3(new_n327), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G125), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT76), .ZN(new_n341));
  OR3_X1    g155(.A1(new_n337), .A2(KEYINPUT76), .A3(G125), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n343), .A2(new_n208), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n208), .B1(new_n343), .B2(new_n345), .ZN(new_n347));
  OAI221_X1 g161(.A(new_n331), .B1(new_n332), .B2(new_n336), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  XNOR2_X1  g164(.A(G125), .B(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n208), .ZN(new_n352));
  INV_X1    g166(.A(G110), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n326), .A2(new_n353), .A3(new_n327), .A4(new_n329), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n336), .A2(new_n332), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT77), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT77), .B1(new_n354), .B2(new_n355), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n350), .B(new_n352), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n348), .A2(new_n358), .A3(new_n363), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n321), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n365), .A2(KEYINPUT25), .A3(new_n321), .A4(new_n366), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n323), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n322), .A2(G902), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n210), .B2(G128), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n207), .A2(KEYINPUT90), .A3(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n210), .A2(G128), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n195), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n378), .A2(new_n379), .B1(G128), .B2(new_n210), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G134), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n240), .A2(new_n242), .A3(G122), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n386), .B(new_n387), .C1(new_n233), .C2(G122), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n390));
  OAI21_X1  g204(.A(G107), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n233), .A2(G122), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n235), .B2(G122), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT91), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n386), .B(new_n390), .C1(new_n233), .C2(G122), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n235), .A2(KEYINPUT14), .A3(G122), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(G107), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n393), .A2(new_n387), .B1(new_n384), .B2(G134), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT91), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n383), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n386), .B1(new_n233), .B2(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G107), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n380), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G134), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n404), .A2(new_n388), .B1(new_n407), .B2(new_n384), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n384), .B2(new_n407), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT9), .B(G234), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT78), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n411), .A2(new_n320), .A3(G953), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n402), .B2(new_n409), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n376), .B(new_n321), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n400), .B1(new_n419), .B2(new_n398), .ZN(new_n420));
  INV_X1    g234(.A(new_n401), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n409), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n412), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n417), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n376), .A3(new_n321), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(G234), .A2(G237), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n429), .A2(G952), .A3(new_n361), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n429), .A2(G902), .A3(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n418), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n436));
  XNOR2_X1  g250(.A(G113), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(G104), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G237), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n361), .A3(G214), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n210), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT18), .A2(G131), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n337), .A2(KEYINPUT76), .A3(G125), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n351), .B2(KEYINPUT76), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G146), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n352), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT88), .B1(new_n346), .B2(new_n347), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n343), .A2(new_n208), .A3(new_n345), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n350), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT17), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n444), .B2(G131), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n442), .A2(new_n201), .A3(new_n443), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n441), .A2(new_n210), .ZN(new_n461));
  AOI21_X1  g275(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n442), .A2(new_n464), .A3(new_n201), .A4(new_n443), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n458), .B1(new_n466), .B2(new_n457), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n439), .B(new_n451), .C1(new_n456), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n448), .A2(KEYINPUT19), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n351), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n351), .A2(new_n471), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT87), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n466), .B(new_n350), .C1(new_n475), .C2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n451), .ZN(new_n477));
  INV_X1    g291(.A(new_n439), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(G475), .A2(G902), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n436), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  AOI211_X1 g297(.A(KEYINPUT20), .B(new_n483), .C1(new_n468), .C2(new_n479), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n451), .B1(new_n456), .B2(new_n467), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n486), .B2(new_n468), .ZN(new_n487));
  INV_X1    g301(.A(G475), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n482), .A2(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n435), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G214), .B1(G237), .B2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n243), .A2(KEYINPUT5), .A3(new_n244), .ZN(new_n496));
  INV_X1    g310(.A(G113), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT5), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n234), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n496), .A2(new_n499), .B1(new_n236), .B2(new_n238), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n387), .A2(KEYINPUT81), .A3(G104), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n438), .B2(G107), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n387), .A2(G104), .ZN(new_n504));
  OAI211_X1 g318(.A(G101), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT3), .B1(new_n438), .B2(G107), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT3), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n387), .A3(G104), .ZN(new_n508));
  INV_X1    g322(.A(G101), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n438), .A2(G107), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT82), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n511), .A3(KEYINPUT82), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n500), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n518));
  AND2_X1   g332(.A1(KEYINPUT80), .A2(G101), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT4), .A3(new_n511), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n247), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G110), .B(G122), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT6), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n253), .A2(G125), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n361), .A2(G224), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n228), .A2(new_n339), .A3(new_n212), .A4(new_n218), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n536), .A3(new_n526), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n529), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n505), .A2(new_n511), .A3(KEYINPUT84), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n512), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n500), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n525), .B(KEYINPUT8), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n500), .B2(new_n539), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT85), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n531), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n533), .B2(new_n534), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n496), .A2(new_n499), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n239), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n505), .A2(new_n511), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(KEYINPUT84), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n500), .A2(new_n539), .A3(new_n541), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n543), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n530), .A2(new_n532), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n528), .B1(new_n557), .B2(new_n547), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n321), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n495), .B1(new_n538), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n556), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n529), .A2(new_n535), .A3(new_n537), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n321), .A4(new_n494), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n493), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G221), .B1(new_n411), .B2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n361), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT79), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n228), .A2(new_n212), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n551), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n520), .A2(new_n254), .A3(new_n522), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n226), .A2(new_n229), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n514), .A2(KEYINPUT10), .A3(new_n515), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n570), .B1(new_n579), .B2(new_n258), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n505), .A2(new_n511), .A3(KEYINPUT82), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT82), .B1(new_n505), .B2(new_n511), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n226), .A4(new_n229), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n200), .B(new_n256), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n575), .A4(new_n576), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT83), .A3(new_n570), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n579), .A2(new_n258), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n582), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n570), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n512), .A2(new_n212), .A3(new_n228), .A4(new_n218), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n573), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT12), .B1(new_n594), .B2(new_n258), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n596), .B(new_n587), .C1(new_n573), .C2(new_n593), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n579), .A2(new_n258), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n592), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n591), .A2(G469), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G469), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n580), .A2(new_n598), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n570), .B1(new_n590), .B2(new_n588), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n602), .B(new_n321), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n602), .A2(new_n321), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n566), .B1(new_n601), .B2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n491), .A2(new_n565), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n319), .A2(new_n375), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AOI21_X1  g426(.A(G902), .B1(new_n272), .B2(new_n286), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n591), .A2(G469), .A3(new_n600), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n605), .A3(new_n607), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(new_n375), .A3(new_n566), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n615), .A2(new_n287), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n426), .A2(KEYINPUT33), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n424), .A2(new_n621), .A3(new_n425), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n622), .A3(G478), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n416), .A2(new_n321), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n424), .B2(new_n425), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n416), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n489), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n564), .A2(new_n434), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  INV_X1    g451(.A(new_n468), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n463), .A2(new_n465), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT17), .B1(new_n639), .B2(new_n460), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n452), .B(new_n455), .C1(new_n640), .C2(new_n458), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n439), .B1(new_n641), .B2(new_n451), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n321), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n637), .A2(new_n482), .B1(new_n643), .B2(G475), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n480), .A2(new_n481), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT20), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n480), .A2(new_n436), .A3(new_n481), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(KEYINPUT95), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n418), .A2(new_n428), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n644), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n630), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n619), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n387), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  OAI211_X1 g469(.A(new_n316), .B(new_n490), .C1(new_n613), .C2(new_n614), .ZN(new_n656));
  INV_X1    g470(.A(new_n566), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT10), .B1(new_n551), .B2(new_n572), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n517), .B(new_n521), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(new_n254), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n587), .B1(new_n660), .B2(new_n586), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n592), .B1(new_n599), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n588), .B(new_n570), .C1(new_n597), .C2(new_n595), .ZN(new_n663));
  AOI21_X1  g477(.A(G902), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n606), .B1(new_n664), .B2(new_n602), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n657), .B1(new_n665), .B2(new_n616), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n359), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n373), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n369), .A2(new_n370), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n323), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n666), .A2(new_n564), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n656), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n430), .B1(new_n431), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n649), .A2(new_n644), .A3(new_n648), .A4(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n666), .A3(new_n564), .A4(new_n672), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n319), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XOR2_X1   g498(.A(new_n678), .B(KEYINPUT39), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n609), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT40), .Z(new_n688));
  OAI21_X1  g502(.A(new_n309), .B1(new_n287), .B2(new_n310), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n316), .A2(KEYINPUT73), .A3(new_n317), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n304), .A2(new_n193), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n288), .A2(new_n289), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n693), .B2(new_n273), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n614), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n287), .B2(KEYINPUT32), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n489), .A2(new_n649), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n672), .A2(new_n699), .A3(new_n493), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n560), .A2(new_n563), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n688), .A2(new_n698), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n210), .ZN(G45));
  AND4_X1   g520(.A1(new_n489), .A2(new_n623), .A3(new_n626), .A4(new_n679), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n666), .A3(new_n564), .A4(new_n672), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n319), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT100), .B(G146), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G48));
  OAI21_X1  g526(.A(new_n321), .B1(new_n603), .B2(new_n604), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n714), .A2(new_n566), .A3(new_n605), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n319), .A2(new_n375), .A3(new_n631), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT101), .ZN(new_n717));
  INV_X1    g531(.A(new_n375), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n691), .B2(new_n308), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n631), .A4(new_n715), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT102), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n722), .B(new_n724), .ZN(G15));
  NAND4_X1  g539(.A1(new_n319), .A2(new_n375), .A3(new_n651), .A4(new_n715), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND4_X1  g541(.A1(new_n715), .A2(new_n490), .A3(new_n564), .A4(new_n672), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n691), .B2(new_n308), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n324), .ZN(G21));
  AOI21_X1  g544(.A(new_n193), .B1(new_n295), .B2(new_n290), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n187), .B1(new_n315), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n375), .B(new_n732), .C1(new_n613), .C2(new_n614), .ZN(new_n733));
  INV_X1    g547(.A(new_n699), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n715), .A3(new_n564), .A4(new_n434), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(G122), .Z(G24));
  OAI211_X1 g551(.A(new_n672), .B(new_n732), .C1(new_n613), .C2(new_n614), .ZN(new_n738));
  INV_X1    g552(.A(new_n707), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n715), .A2(new_n564), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n339), .ZN(G27));
  AND3_X1   g556(.A1(new_n560), .A2(new_n563), .A3(new_n492), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n617), .A3(new_n744), .A4(new_n566), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(new_n666), .B2(new_n743), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n319), .A2(new_n748), .A3(new_n375), .A4(new_n707), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(KEYINPUT104), .A3(new_n750), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n718), .B1(new_n308), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n739), .A2(new_n750), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n748), .A3(KEYINPUT105), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n307), .A2(G472), .ZN(new_n760));
  OAI211_X1 g574(.A(KEYINPUT32), .B(new_n187), .C1(new_n314), .C2(new_n315), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n375), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n560), .A2(new_n563), .A3(new_n492), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT103), .B1(new_n609), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n707), .A4(new_n745), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n759), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n753), .A2(new_n754), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND4_X1  g585(.A1(new_n319), .A2(new_n748), .A3(new_n375), .A4(new_n680), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NOR2_X1   g587(.A1(new_n627), .A2(new_n489), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(KEYINPUT43), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n672), .B1(new_n615), .B2(new_n287), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT44), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n780), .B2(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n765), .B1(new_n780), .B2(KEYINPUT44), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n591), .A2(new_n600), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT106), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n602), .B1(new_n789), .B2(new_n790), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n788), .B1(new_n794), .B2(new_n606), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n793), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n607), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n605), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(new_n566), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n782), .A2(KEYINPUT108), .A3(new_n783), .A4(new_n784), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n787), .A2(new_n685), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(new_n319), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n718), .A3(new_n707), .A4(new_n743), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n798), .A2(new_n566), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n804), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n337), .ZN(G42));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n805), .A2(new_n808), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n714), .A2(new_n605), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n657), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n776), .A2(new_n430), .A3(new_n777), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n733), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n743), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT117), .Z(new_n818));
  NOR2_X1   g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n492), .B1(KEYINPUT118), .B2(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n704), .A2(new_n816), .A3(new_n715), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(KEYINPUT118), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n824), .ZN(new_n826));
  INV_X1    g640(.A(new_n813), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n815), .A2(new_n657), .A3(new_n827), .A4(new_n765), .ZN(new_n828));
  INV_X1    g642(.A(new_n738), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n489), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n375), .A2(new_n715), .A3(new_n430), .A4(new_n743), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n698), .A2(new_n831), .A3(new_n627), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n826), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n811), .B1(new_n819), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT51), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n811), .B(new_n837), .C1(new_n819), .C2(new_n834), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n828), .A2(new_n756), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n361), .A2(G952), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n698), .A2(new_n832), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n629), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n815), .A2(new_n740), .A3(new_n733), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n841), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n836), .A2(new_n838), .A3(new_n846), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n733), .A2(new_n735), .B1(new_n656), .B2(new_n673), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n729), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n418), .A2(new_n428), .A3(KEYINPUT110), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT110), .B1(new_n418), .B2(new_n428), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n831), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT111), .B(new_n831), .C1(new_n850), .C2(new_n851), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n629), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n630), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n619), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n849), .A2(new_n611), .A3(new_n726), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n721), .B2(new_n717), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n691), .A2(new_n308), .B1(new_n681), .B2(new_n708), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n741), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n672), .A2(new_n678), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n666), .A3(new_n564), .A4(new_n734), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n697), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n861), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n865), .B1(new_n691), .B2(new_n696), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n862), .A2(new_n869), .A3(KEYINPUT52), .A4(new_n741), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n738), .A2(new_n739), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n748), .A2(new_n872), .A3(KEYINPUT112), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n766), .A2(new_n745), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n321), .B1(new_n314), .B2(new_n315), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G472), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n672), .A3(new_n707), .A4(new_n732), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n609), .A2(new_n765), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n672), .A2(new_n648), .A3(new_n644), .A4(new_n679), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n882), .A2(new_n850), .A3(new_n851), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n319), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n880), .A2(new_n772), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n860), .A2(new_n871), .A3(new_n770), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n886), .A2(KEYINPUT114), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n848), .ZN(new_n889));
  INV_X1    g703(.A(new_n728), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n319), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n611), .A2(new_n889), .A3(new_n891), .A4(new_n858), .ZN(new_n892));
  INV_X1    g706(.A(new_n726), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n885), .A3(new_n722), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n754), .A2(new_n769), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT104), .B1(new_n749), .B2(new_n750), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n319), .B1(new_n682), .B2(new_n709), .ZN(new_n900));
  INV_X1    g714(.A(new_n741), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n867), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT113), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT52), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT114), .B1(new_n886), .B2(new_n887), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n888), .B(KEYINPUT54), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(KEYINPUT52), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n863), .A2(new_n861), .A3(new_n867), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n895), .A2(new_n898), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n908), .B1(new_n912), .B2(KEYINPUT53), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n894), .A2(new_n885), .A3(new_n722), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n904), .A2(new_n914), .A3(KEYINPUT53), .A4(new_n770), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n886), .A2(KEYINPUT115), .A3(new_n887), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n907), .B1(KEYINPUT54), .B2(new_n917), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n847), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n704), .B1(KEYINPUT49), .B2(new_n827), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n718), .A2(new_n657), .A3(new_n493), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n922), .A3(new_n774), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT109), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n924), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n919), .B1(new_n697), .B2(new_n926), .ZN(G75));
  AND2_X1   g741(.A1(new_n917), .A2(G902), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(G210), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n529), .A2(new_n537), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n535), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n361), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n917), .B(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n606), .B(KEYINPUT57), .Z(new_n940));
  OAI22_X1  g754(.A1(new_n939), .A2(new_n940), .B1(new_n604), .B2(new_n603), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n928), .A2(new_n794), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(G54));
  NAND3_X1  g757(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n479), .A3(new_n468), .ZN(new_n945));
  INV_X1    g759(.A(new_n936), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .A4(new_n480), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G60));
  AND2_X1   g762(.A1(new_n620), .A2(new_n622), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n624), .B(KEYINPUT59), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n946), .B1(new_n939), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n950), .B1(new_n918), .B2(new_n951), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G63));
  INV_X1    g769(.A(KEYINPUT120), .ZN(new_n956));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT60), .Z(new_n958));
  AOI21_X1  g772(.A(new_n372), .B1(new_n917), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n956), .B1(new_n959), .B2(new_n936), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n916), .A2(new_n915), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT115), .B1(new_n886), .B2(new_n887), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n372), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(KEYINPUT120), .A3(new_n946), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n917), .A2(new_n669), .A3(new_n958), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n960), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n967), .A4(new_n946), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n936), .B1(new_n963), .B2(new_n964), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n967), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n970), .A2(new_n976), .ZN(G66));
  XOR2_X1   g791(.A(new_n860), .B(KEYINPUT122), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n361), .ZN(new_n979));
  INV_X1    g793(.A(G224), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n432), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n931), .B1(G898), .B2(new_n361), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G69));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n734), .A2(new_n564), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n806), .A2(new_n686), .A3(new_n764), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n863), .A2(new_n772), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n809), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(new_n801), .A3(new_n361), .A4(new_n770), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n265), .B(new_n475), .Z(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(G900), .B2(G953), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n705), .A2(new_n741), .A3(new_n862), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT62), .ZN(new_n995));
  INV_X1    g809(.A(new_n809), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n719), .A2(new_n685), .A3(new_n881), .A4(new_n856), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n995), .A2(new_n801), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n998), .A2(new_n361), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n991), .B(KEYINPUT123), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n985), .B(new_n993), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n990), .A2(new_n992), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n998), .B2(new_n361), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT124), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n361), .B1(G227), .B2(G900), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(G72));
  XNOR2_X1  g823(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n989), .A2(new_n801), .A3(new_n770), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n978), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n305), .ZN(new_n1015));
  INV_X1    g829(.A(new_n692), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1012), .B1(new_n304), .B2(new_n193), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n888), .B(new_n1018), .C1(new_n905), .C2(new_n906), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1015), .A2(new_n946), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1012), .B1(new_n998), .B2(new_n978), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(KEYINPUT126), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1023), .B(new_n1012), .C1(new_n998), .C2(new_n978), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1022), .A2(new_n1016), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1022), .A2(KEYINPUT127), .A3(new_n1016), .A4(new_n1024), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(G57));
endmodule


