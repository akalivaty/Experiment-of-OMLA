//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n211), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G77), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n223), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT68), .Z(new_n233));
  AOI211_X1 g0033(.A(new_n219), .B(new_n233), .C1(KEYINPUT1), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G58), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(G1698), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(new_n228), .B2(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n259), .A3(G274), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n262), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(G226), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n212), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n202), .A2(G20), .ZN(new_n273));
  XOR2_X1   g0073(.A(KEYINPUT8), .B(G58), .Z(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G20), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n274), .A2(new_n276), .B1(G150), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n272), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n271), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n205), .A2(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G50), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G50), .B2(new_n280), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n269), .A2(G169), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n261), .A2(new_n268), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G179), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n279), .A2(new_n285), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT9), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n269), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n291), .A2(KEYINPUT9), .B1(new_n287), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n294), .A2(KEYINPUT10), .A3(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G107), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n256), .A2(new_n226), .B1(new_n302), .B2(new_n252), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n307), .A2(new_n236), .A3(G1698), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n260), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n265), .B1(G244), .B2(new_n267), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G169), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  INV_X1    g0113(.A(new_n276), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT70), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n227), .A2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(new_n274), .ZN(new_n317));
  INV_X1    g0117(.A(new_n277), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT70), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n271), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n283), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n282), .A2(new_n324), .B1(new_n228), .B2(new_n281), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n312), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n311), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n321), .A2(new_n325), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n311), .B2(G190), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n293), .B2(new_n311), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n301), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n252), .A2(G226), .A3(new_n253), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n264), .B1(new_n226), .B2(new_n266), .C1(new_n338), .C2(new_n259), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT13), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n343), .A3(G169), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n344), .C1(new_n327), .C2(new_n340), .ZN(new_n345));
  INV_X1    g0145(.A(new_n282), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n346), .A2(new_n216), .A3(new_n322), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n225), .A2(G20), .ZN(new_n348));
  INV_X1    g0148(.A(G13), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G1), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n348), .A2(KEYINPUT12), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT12), .B1(new_n281), .B2(new_n216), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n347), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT11), .ZN(new_n354));
  INV_X1    g0154(.A(G50), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n314), .A2(new_n323), .B1(new_n355), .B2(new_n318), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n271), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n353), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n357), .A2(new_n354), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n340), .A2(new_n295), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n340), .A2(G200), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n334), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n217), .B1(new_n225), .B2(new_n215), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n277), .A2(G159), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n252), .B2(G20), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n307), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n225), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n367), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n252), .A2(new_n374), .A3(G20), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n307), .B2(new_n206), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n369), .A4(new_n372), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n382), .A3(new_n271), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n274), .A2(new_n283), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n346), .B1(new_n384), .B2(KEYINPUT72), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(KEYINPUT72), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n385), .A2(new_n386), .B1(new_n281), .B2(new_n317), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n304), .A2(new_n306), .A3(G226), .A4(G1698), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n304), .A2(new_n306), .A3(G223), .A4(new_n253), .ZN(new_n390));
  INV_X1    g0190(.A(G87), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n390), .C1(new_n275), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n260), .ZN(new_n393));
  INV_X1    g0193(.A(G274), .ZN(new_n394));
  INV_X1    g0194(.A(new_n212), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n258), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n267), .A2(G232), .B1(new_n396), .B2(new_n263), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n397), .A3(G179), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n264), .B1(new_n236), .B2(new_n266), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n260), .B2(new_n392), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n398), .B(KEYINPUT73), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT73), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n388), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT18), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n383), .A2(new_n387), .B1(new_n403), .B2(new_n404), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n402), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n393), .A2(new_n397), .A3(G190), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n293), .B1(new_n393), .B2(new_n397), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n383), .A3(new_n387), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n413), .A2(new_n383), .A3(KEYINPUT17), .A4(new_n387), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n416), .A2(KEYINPUT74), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT74), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n407), .B(new_n410), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n366), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G283), .ZN(new_n422));
  INV_X1    g0222(.A(G97), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n206), .C1(G33), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT80), .ZN(new_n425));
  AOI21_X1  g0225(.A(G20), .B1(new_n275), .B2(G97), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n422), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G116), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G20), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n271), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT81), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT20), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n205), .A2(G33), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n280), .A2(new_n438), .A3(new_n212), .A4(new_n270), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n439), .A2(KEYINPUT79), .A3(new_n430), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT79), .B1(new_n439), .B2(new_n430), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n281), .A2(new_n430), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n445), .A2(new_n447), .B1(new_n395), .B2(new_n258), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n205), .A2(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n448), .A2(G270), .B1(new_n396), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n305), .A2(G33), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n456));
  OAI21_X1  g0256(.A(G303), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n304), .A2(new_n306), .A3(G264), .A4(G1698), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n304), .A2(new_n306), .A3(G257), .A4(new_n253), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n260), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G200), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n434), .A2(new_n436), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n432), .B1(new_n425), .B2(new_n428), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT20), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(KEYINPUT81), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n462), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G190), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT81), .B1(new_n465), .B2(KEYINPUT20), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n436), .B(new_n432), .C1(new_n428), .C2(new_n425), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT82), .B1(new_n476), .B2(new_n463), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n462), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G179), .B(new_n469), .C1(new_n472), .C2(new_n475), .ZN(new_n482));
  INV_X1    g0282(.A(new_n480), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(KEYINPUT21), .C1(new_n475), .C2(new_n472), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n304), .A3(new_n306), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G294), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n304), .A2(new_n306), .A3(G257), .A4(G1698), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n488), .A2(new_n304), .A3(new_n306), .A4(KEYINPUT85), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n260), .ZN(new_n496));
  INV_X1    g0296(.A(new_n452), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n447), .B1(new_n497), .B2(new_n450), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G264), .A3(new_n259), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(KEYINPUT86), .A3(G264), .A4(new_n259), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n453), .A2(new_n396), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n496), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n496), .A2(new_n503), .A3(KEYINPUT87), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(G169), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n505), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G179), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n304), .A2(new_n306), .A3(new_n206), .A4(G87), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n252), .A2(new_n515), .A3(new_n206), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G20), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n206), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n302), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n518), .B1(new_n517), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n271), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR3_X1    g0330(.A1(new_n280), .A2(KEYINPUT25), .A3(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT25), .B1(new_n280), .B2(G107), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n302), .C2(new_n439), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT84), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(KEYINPUT83), .B(new_n271), .C1(new_n526), .C2(new_n527), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n512), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n527), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n272), .B1(new_n539), .B2(new_n525), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n534), .B1(new_n540), .B2(KEYINPUT83), .ZN(new_n541));
  AOI21_X1  g0341(.A(G190), .B1(new_n507), .B2(new_n508), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n510), .A2(G200), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n530), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n226), .A2(new_n253), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n229), .A2(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n252), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n259), .B1(new_n548), .B2(new_n519), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n259), .A2(G274), .A3(new_n447), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n259), .A2(G250), .A3(new_n449), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT77), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT77), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n519), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n260), .ZN(new_n558));
  INV_X1    g0358(.A(new_n554), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n552), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  OR2_X1    g0361(.A1(KEYINPUT78), .A2(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(KEYINPUT78), .A2(G87), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n423), .A3(new_n302), .A4(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n206), .B1(new_n337), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n314), .B2(new_n423), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n252), .A2(new_n206), .A3(G68), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n271), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n313), .A2(new_n281), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n439), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G87), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n556), .A2(new_n561), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n560), .A2(new_n401), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n572), .C1(new_n313), .C2(new_n439), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(G179), .C2(new_n560), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n304), .A2(new_n306), .A3(G244), .A4(new_n253), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT75), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n304), .A2(new_n306), .A3(G250), .A4(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n422), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n583), .A3(new_n581), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n259), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n448), .A2(G257), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n504), .ZN(new_n591));
  OR3_X1    g0391(.A1(new_n589), .A2(new_n295), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n423), .A3(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(G97), .B(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(new_n206), .B1(new_n323), .B2(new_n318), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n302), .B1(new_n375), .B2(new_n376), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n271), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n281), .A2(new_n423), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n574), .A2(G97), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n590), .A2(KEYINPUT76), .A3(new_n504), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT76), .B1(new_n590), .B2(new_n504), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n589), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n592), .B(new_n603), .C1(new_n606), .C2(new_n293), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n604), .A2(new_n605), .ZN(new_n608));
  INV_X1    g0408(.A(new_n589), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n327), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n401), .B1(new_n589), .B2(new_n591), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n602), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n580), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n421), .A2(new_n486), .A3(new_n545), .A4(new_n613), .ZN(G372));
  AND3_X1   g0414(.A1(new_n610), .A2(new_n611), .A3(new_n602), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n580), .A2(new_n615), .A3(KEYINPUT26), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n576), .A2(new_n579), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n613), .A2(new_n544), .ZN(new_n621));
  INV_X1    g0421(.A(new_n538), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n485), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n579), .B(new_n620), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n421), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(KEYINPUT88), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n388), .A2(new_n403), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(new_n409), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n365), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n362), .B1(new_n630), .B2(new_n329), .ZN(new_n631));
  INV_X1    g0431(.A(new_n419), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n416), .A2(KEYINPUT74), .A3(new_n417), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n629), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n297), .B(new_n298), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n290), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n626), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n476), .A2(new_n463), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT82), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n470), .A3(new_n468), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n484), .A2(new_n482), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n444), .A2(new_n467), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n350), .A2(new_n206), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n644), .A2(new_n645), .A3(new_n481), .A4(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n485), .A2(new_n646), .A3(new_n652), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n537), .A2(new_n652), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n545), .A2(new_n658), .B1(new_n622), .B2(new_n652), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n640), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n654), .B2(new_n655), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n538), .A2(new_n544), .A3(new_n658), .ZN(new_n663));
  INV_X1    g0463(.A(new_n652), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n538), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(KEYINPUT89), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n538), .A2(new_n652), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n485), .A2(new_n664), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n670), .B2(new_n545), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT90), .Z(G399));
  INV_X1    g0473(.A(new_n209), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n564), .A2(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n218), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n624), .B2(new_n664), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n624), .A2(new_n681), .A3(new_n664), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n545), .A2(new_n486), .A3(new_n613), .A4(new_n664), .ZN(new_n686));
  XOR2_X1   g0486(.A(KEYINPUT93), .B(KEYINPUT30), .Z(new_n687));
  NAND3_X1  g0487(.A1(new_n454), .A2(new_n461), .A3(G179), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n589), .A2(new_n688), .A3(new_n591), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n496), .A2(new_n503), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n560), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n555), .A2(KEYINPUT91), .A3(new_n496), .A4(new_n503), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT92), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT92), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n689), .A2(new_n692), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n687), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n505), .A2(new_n327), .A3(new_n462), .A4(new_n560), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n694), .A2(new_n699), .B1(new_n700), .B2(new_n606), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT31), .B(new_n652), .C1(new_n698), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n686), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n652), .B1(new_n698), .B2(new_n701), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT94), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(KEYINPUT94), .A3(new_n705), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n661), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n685), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n680), .B1(new_n710), .B2(G1), .ZN(G364));
  NOR2_X1   g0511(.A1(new_n349), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n205), .B1(new_n712), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n675), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n662), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(G330), .B2(new_n656), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n212), .B1(G20), .B2(new_n401), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n206), .A2(G179), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n562), .B2(new_n563), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n206), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n721), .B1(G97), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n206), .A2(new_n327), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n295), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n719), .A2(new_n295), .A3(G200), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n725), .B1(new_n355), .B2(new_n729), .C1(new_n302), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n719), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G159), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n733), .A2(KEYINPUT32), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT32), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n727), .A2(G190), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n738), .B2(new_n216), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n726), .A2(G190), .A3(new_n293), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n726), .A2(new_n732), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n252), .B1(new_n740), .B2(new_n215), .C1(new_n228), .C2(new_n741), .ZN(new_n742));
  NOR4_X1   g0542(.A1(new_n731), .A2(new_n735), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n728), .B(KEYINPUT97), .ZN(new_n744));
  INV_X1    g0544(.A(G326), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n720), .B(KEYINPUT98), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G303), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n744), .A2(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n740), .ZN(new_n750));
  INV_X1    g0550(.A(new_n733), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(G322), .B1(new_n751), .B2(G329), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n307), .C1(new_n753), .C2(new_n741), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n737), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n758), .B1(new_n759), .B2(new_n730), .C1(new_n760), .C2(new_n723), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n749), .A2(new_n754), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n718), .B1(new_n743), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n715), .B(KEYINPUT95), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n674), .A2(new_n252), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n218), .ZN(new_n767));
  INV_X1    g0567(.A(new_n250), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G45), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n209), .A2(new_n252), .ZN(new_n770));
  INV_X1    g0570(.A(G355), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(G116), .B2(new_n209), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n769), .B1(KEYINPUT96), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(KEYINPUT96), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n718), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n765), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n763), .B(new_n779), .C1(new_n656), .C2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n717), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  INV_X1    g0583(.A(new_n718), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n776), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n764), .B1(G77), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT99), .Z(new_n787));
  AOI22_X1  g0587(.A1(new_n750), .A2(G294), .B1(new_n751), .B2(G311), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(new_n307), .C1(new_n430), .C2(new_n741), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n730), .A2(new_n391), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G283), .B2(new_n737), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n791), .B1(new_n423), .B2(new_n723), .C1(new_n748), .C2(new_n729), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n789), .B(new_n792), .C1(G107), .C2(new_n746), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n252), .B1(new_n733), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n730), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(G68), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n215), .B2(new_n723), .ZN(new_n798));
  INV_X1    g0598(.A(new_n741), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n750), .A2(G143), .B1(new_n799), .B2(G159), .ZN(new_n800));
  INV_X1    g0600(.A(G150), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(new_n738), .B2(new_n801), .C1(new_n802), .C2(new_n729), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT34), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n798), .B(new_n805), .C1(G50), .C2(new_n746), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n793), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n330), .A2(new_n652), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n332), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n329), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n329), .A2(new_n652), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n787), .B1(new_n784), .B2(new_n808), .C1(new_n814), .C2(new_n776), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n624), .A2(new_n664), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(new_n814), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n704), .A2(new_n705), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT94), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n822), .A2(new_n708), .A3(new_n702), .A4(new_n686), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G330), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n715), .B1(new_n819), .B2(new_n824), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n816), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G384));
  NOR2_X1   g0629(.A1(new_n712), .A2(new_n205), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n624), .A2(new_n664), .A3(new_n814), .ZN(new_n831));
  INV_X1    g0631(.A(new_n813), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n361), .A2(new_n652), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n362), .A2(new_n365), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n361), .B(new_n652), .C1(new_n630), .C2(new_n345), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n216), .B1(new_n375), .B2(new_n376), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n367), .B1(new_n373), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n382), .A3(new_n271), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n387), .ZN(new_n842));
  INV_X1    g0642(.A(new_n650), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n403), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(new_n845), .A3(new_n414), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT37), .B1(new_n408), .B2(new_n402), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n413), .A2(new_n383), .A3(new_n387), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n650), .B1(new_n383), .B2(new_n387), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(KEYINPUT37), .A2(new_n846), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n407), .A2(new_n410), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n632), .B2(new_n633), .ZN(new_n854));
  OAI211_X1 g0654(.A(KEYINPUT38), .B(new_n852), .C1(new_n854), .C2(new_n844), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n844), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n628), .A2(new_n843), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n844), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n420), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n863), .B2(new_n852), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n857), .B(new_n851), .C1(new_n420), .C2(new_n862), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT39), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n416), .A2(new_n417), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT100), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n416), .A2(KEYINPUT100), .A3(new_n417), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n628), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n847), .A2(new_n850), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n850), .A2(new_n627), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n872), .A2(new_n849), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n855), .B(new_n867), .C1(new_n876), .C2(KEYINPUT38), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n345), .A2(new_n361), .A3(new_n664), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n876), .A2(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT101), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n867), .A4(new_n855), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n861), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n638), .B1(new_n421), .B2(new_n685), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT102), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n886), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n855), .B1(new_n876), .B2(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n814), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n835), .B2(new_n836), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n686), .A2(new_n702), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n652), .C1(new_n698), .C2(new_n701), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n705), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n893), .A2(new_n897), .A3(KEYINPUT104), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT104), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n890), .B(new_n892), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(new_n897), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n893), .A2(new_n897), .A3(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT40), .B1(new_n858), .B2(new_n855), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n892), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n421), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n904), .B2(new_n905), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n661), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n911), .B2(new_n909), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n830), .B1(new_n889), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n889), .B2(new_n913), .ZN(new_n915));
  INV_X1    g0715(.A(new_n596), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n430), .B(new_n214), .C1(new_n916), .C2(KEYINPUT35), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(KEYINPUT35), .B2(new_n916), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  INV_X1    g0719(.A(new_n218), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n227), .C1(new_n215), .C2(new_n225), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(G50), .B2(new_n216), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n349), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(new_n919), .A3(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n573), .A2(new_n575), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n652), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n580), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n579), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT105), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT106), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n602), .A2(new_n652), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n607), .A2(new_n612), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n615), .A2(new_n652), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT107), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT107), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND4_X1   g0742(.A1(new_n485), .A2(new_n538), .A3(new_n544), .A4(new_n664), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT42), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n938), .B(new_n939), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT42), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(new_n943), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n615), .B1(new_n946), .B2(new_n622), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n945), .B(new_n948), .C1(new_n949), .C2(new_n652), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT108), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n951), .B1(new_n950), .B2(new_n952), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n934), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n667), .A2(new_n942), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n950), .A2(new_n952), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n959));
  INV_X1    g0759(.A(new_n934), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n953), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n956), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n954), .A2(new_n955), .A3(new_n934), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n959), .B2(new_n953), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n963), .A2(new_n964), .B1(new_n667), .B2(new_n942), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n675), .B(KEYINPUT41), .Z(new_n966));
  OAI211_X1 g0766(.A(new_n942), .B(KEYINPUT44), .C1(new_n668), .C2(new_n943), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n946), .B2(new_n671), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n671), .B1(new_n941), .B2(new_n940), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n946), .A2(new_n671), .A3(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n970), .A2(new_n975), .A3(new_n667), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n667), .B1(new_n970), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT109), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n657), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n943), .B1(new_n659), .B2(new_n669), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n662), .A2(KEYINPUT109), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n944), .B1(new_n665), .B2(new_n670), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(KEYINPUT109), .A3(new_n662), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n710), .A2(KEYINPUT110), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n684), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n682), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n986), .A3(new_n824), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT110), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n978), .A2(new_n987), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n966), .B1(new_n993), .B2(new_n710), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n962), .B(new_n965), .C1(new_n994), .C2(new_n714), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n778), .B1(new_n209), .B2(new_n313), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n766), .B2(new_n242), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n765), .A2(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n740), .A2(new_n748), .B1(new_n733), .B2(new_n755), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n252), .B(new_n999), .C1(G283), .C2(new_n799), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n730), .A2(new_n423), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n723), .A2(new_n302), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G294), .C2(new_n737), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n720), .A2(new_n430), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1003), .C1(KEYINPUT46), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n746), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n744), .B2(new_n753), .ZN(new_n1007));
  INV_X1    g0807(.A(G143), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n744), .A2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n724), .A2(G68), .B1(new_n796), .B2(new_n227), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n720), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n737), .A2(G159), .B1(new_n1011), .B2(G58), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n307), .B1(new_n750), .B2(G150), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G50), .A2(new_n799), .B1(new_n751), .B2(G137), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1005), .A2(new_n1007), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT47), .Z(new_n1017));
  OAI221_X1 g0817(.A(new_n998), .B1(new_n784), .B2(new_n1017), .C1(new_n932), .C2(new_n780), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n995), .A2(new_n1018), .ZN(G387));
  NAND2_X1  g0819(.A1(new_n987), .A2(new_n992), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n675), .B(KEYINPUT113), .Z(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n710), .C2(new_n986), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n659), .A2(new_n777), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n770), .A2(new_n677), .B1(G107), .B2(new_n209), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n239), .A2(new_n446), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT111), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n677), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n274), .A2(new_n355), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT50), .Z(new_n1030));
  AOI211_X1 g0830(.A(new_n674), .B(new_n252), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1024), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n778), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n764), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n728), .A2(G159), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT112), .Z(new_n1036));
  OAI22_X1  g0836(.A1(new_n740), .A2(new_n355), .B1(new_n741), .B2(new_n216), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n307), .B(new_n1037), .C1(G150), .C2(new_n751), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n228), .A2(new_n720), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n1001), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n723), .A2(new_n313), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n274), .B2(new_n737), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n750), .A2(G317), .B1(new_n799), .B2(G303), .ZN(new_n1044));
  INV_X1    g0844(.A(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n753), .B2(new_n738), .C1(new_n744), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n724), .A2(G283), .B1(new_n1011), .B2(G294), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n307), .B1(new_n733), .B2(new_n745), .C1(new_n430), .C2(new_n730), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1043), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1034), .B1(new_n1057), .B2(new_n718), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n986), .A2(new_n714), .B1(new_n1023), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1022), .A2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n247), .A2(new_n766), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1033), .B1(G97), .B2(new_n674), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n765), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n729), .A2(new_n755), .B1(new_n753), .B2(new_n740), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n738), .A2(new_n748), .B1(new_n730), .B2(new_n302), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n307), .B1(new_n733), .B2(new_n1045), .C1(new_n760), .C2(new_n741), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n723), .A2(new_n430), .B1(new_n720), .B2(new_n759), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n738), .A2(new_n355), .B1(new_n720), .B2(new_n225), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n252), .B1(new_n733), .B2(new_n1008), .C1(new_n317), .C2(new_n741), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n723), .A2(new_n323), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n790), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G150), .A2(new_n728), .B1(new_n750), .B2(G159), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1065), .A2(new_n1069), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1063), .B1(new_n784), .B2(new_n1077), .C1(new_n946), .C2(new_n780), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n978), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n713), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1020), .A2(new_n1079), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT115), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT115), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1020), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n993), .A2(new_n1021), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1080), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G390));
  NAND2_X1  g0889(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n867), .B1(new_n858), .B2(new_n855), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n883), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n880), .B1(new_n833), .B2(new_n837), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n709), .A2(KEYINPUT116), .A3(new_n814), .A4(new_n837), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n823), .A2(G330), .A3(new_n837), .A4(new_n814), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT116), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1093), .A2(new_n890), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(G330), .B(new_n892), .C1(new_n898), .C2(new_n899), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1093), .B1(new_n878), .B2(new_n883), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1093), .A2(new_n890), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1092), .A2(new_n775), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n764), .B1(new_n274), .B2(new_n785), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n740), .A2(new_n794), .B1(new_n741), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n307), .B(new_n1112), .C1(G125), .C2(new_n751), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n720), .A2(new_n801), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n737), .A2(G137), .B1(new_n796), .B2(G50), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G159), .A2(new_n724), .B1(new_n728), .B2(G128), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n728), .A2(G283), .B1(new_n799), .B2(G97), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n302), .B2(new_n738), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT118), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1072), .B1(G68), .B2(new_n796), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n307), .B1(new_n733), .B2(new_n760), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G116), .B2(new_n750), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(new_n747), .C2(new_n391), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1118), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1110), .B1(new_n1126), .B2(new_n718), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1108), .A2(new_n714), .B1(new_n1109), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n833), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1129));
  OAI211_X1 g0929(.A(G330), .B(new_n814), .C1(new_n898), .C2(new_n899), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n837), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n823), .A2(G330), .A3(new_n814), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1131), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1103), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1134), .B1(new_n1137), .B2(new_n833), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n833), .ZN(new_n1139));
  AOI211_X1 g0939(.A(KEYINPUT117), .B(new_n1139), .C1(new_n1103), .C2(new_n1136), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1133), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n906), .A2(new_n421), .A3(G330), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n887), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1108), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1021), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1108), .B1(new_n1144), .B2(new_n1141), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1128), .B1(new_n1146), .B2(new_n1147), .ZN(G378));
  NOR2_X1   g0948(.A1(new_n291), .A2(new_n650), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n636), .A2(new_n290), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n301), .A2(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n837), .A2(new_n814), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n904), .B2(new_n905), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(KEYINPUT40), .A2(new_n900), .B1(new_n1161), .B2(new_n907), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1159), .B1(new_n1162), .B2(new_n661), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1156), .A2(KEYINPUT120), .A3(new_n1157), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT120), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n909), .A2(G330), .A3(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1163), .A2(new_n885), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n885), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1166), .A2(new_n775), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n715), .B1(G50), .B2(new_n785), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n252), .A2(G41), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G283), .B2(new_n751), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n302), .B2(new_n740), .C1(new_n313), .C2(new_n741), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1039), .B(new_n1176), .C1(G68), .C2(new_n724), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n728), .A2(G116), .B1(new_n796), .B2(G58), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n423), .C2(new_n738), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT119), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1174), .B(new_n355), .C1(G33), .C2(G41), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n728), .A2(G125), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n738), .B2(new_n794), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n750), .A2(G128), .B1(new_n799), .B2(G137), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n720), .B2(new_n1111), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G150), .C2(new_n724), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n796), .A2(G159), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1173), .B1(new_n1195), .B2(new_n718), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1171), .A2(new_n714), .B1(new_n1172), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1141), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1144), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1158), .B1(new_n909), .B2(G330), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n661), .B(new_n1166), .C1(new_n901), .C2(new_n908), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n886), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1163), .A2(new_n1168), .A3(new_n885), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(KEYINPUT57), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1143), .B1(new_n1108), .B2(new_n1141), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1021), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1197), .B1(new_n1201), .B2(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n966), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1143), .B(new_n1133), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1131), .A2(new_n775), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n764), .B1(G68), .B2(new_n785), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n740), .A2(new_n802), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n252), .B1(new_n741), .B2(new_n801), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G128), .C2(new_n751), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n746), .A2(G159), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n724), .A2(G50), .B1(new_n796), .B2(G58), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1111), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G132), .A2(new_n728), .B1(new_n737), .B2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n728), .A2(G294), .B1(new_n799), .B2(G107), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n430), .B2(new_n738), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT121), .Z(new_n1226));
  OAI21_X1  g1026(.A(new_n307), .B1(new_n740), .B2(new_n759), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1041), .B(new_n1227), .C1(G77), .C2(new_n796), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n746), .A2(G97), .B1(G303), .B2(new_n751), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT122), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1223), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1215), .B1(new_n1232), .B2(new_n718), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1141), .A2(new_n714), .B1(new_n1214), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1213), .A2(new_n1234), .ZN(G381));
  INV_X1    g1035(.A(KEYINPUT123), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(G375), .B(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(G378), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1088), .A2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1240), .A2(G387), .A3(G381), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(new_n1238), .A3(new_n1241), .ZN(G407));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(G343), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1237), .A2(new_n1238), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G407), .A2(new_n1245), .A3(G213), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(G407), .A2(new_n1245), .A3(KEYINPUT124), .A4(G213), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(G409));
  OAI211_X1 g1050(.A(G378), .B(new_n1197), .C1(new_n1201), .C2(new_n1208), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1210), .A2(new_n1199), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n1021), .A3(new_n1145), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1254), .A2(new_n1207), .A3(new_n966), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1172), .A2(new_n1196), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1254), .B2(new_n713), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1253), .B(new_n1128), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1244), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1021), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1137), .A2(new_n833), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT117), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1137), .A2(new_n1134), .A3(new_n833), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1265), .A2(KEYINPUT60), .A3(new_n1143), .A4(new_n1133), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1212), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1234), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT125), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1272), .A3(new_n1234), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(G384), .A3(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1269), .A2(new_n1272), .A3(new_n1234), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1272), .B1(new_n1269), .B2(new_n1234), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n828), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1259), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1244), .A2(G2897), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1275), .A2(new_n1276), .A3(new_n828), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1270), .A2(KEYINPUT125), .A3(G384), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1244), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1274), .A2(new_n1277), .A3(G2897), .A4(new_n1244), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1259), .A2(new_n1278), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1280), .A2(new_n1289), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1088), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1086), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n995), .B(new_n1018), .C1(new_n1295), .C2(new_n1080), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(new_n782), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1300), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1297), .A2(new_n1298), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1293), .A2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1259), .A2(new_n1278), .A3(KEYINPUT63), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1279), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1308), .A2(new_n1290), .A3(new_n1289), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1305), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1238), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1251), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1306), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1313), .A2(new_n1317), .A3(new_n1251), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1318), .A2(new_n1278), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1304), .A2(KEYINPUT127), .A3(new_n1314), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1316), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1316), .B2(new_n1320), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


