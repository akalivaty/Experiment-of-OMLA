

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U549 ( .A1(n677), .A2(n764), .ZN(n721) );
  XNOR2_X1 U550 ( .A(n690), .B(n689), .ZN(n734) );
  XNOR2_X1 U551 ( .A(n688), .B(KEYINPUT102), .ZN(n689) );
  INV_X1 U552 ( .A(KEYINPUT31), .ZN(n688) );
  NOR2_X2 U553 ( .A1(n527), .A2(n526), .ZN(G160) );
  NOR2_X1 U554 ( .A1(n737), .A2(n736), .ZN(n513) );
  NOR2_X1 U555 ( .A1(n972), .A2(n695), .ZN(n701) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n712) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n716) );
  XNOR2_X1 U558 ( .A(n717), .B(n716), .ZN(n720) );
  NAND2_X1 U559 ( .A1(n720), .A2(n719), .ZN(n733) );
  NOR2_X1 U560 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U561 ( .A1(G8), .A2(n721), .ZN(n762) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n864) );
  NOR2_X1 U564 ( .A1(G651), .A2(n625), .ZN(n640) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n515) );
  INV_X1 U566 ( .A(G2105), .ZN(n524) );
  AND2_X1 U567 ( .A1(n524), .A2(G2104), .ZN(n869) );
  NAND2_X1 U568 ( .A1(G101), .A2(n869), .ZN(n514) );
  XNOR2_X1 U569 ( .A(n515), .B(n514), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n864), .A2(G113), .ZN(n516) );
  XOR2_X1 U571 ( .A(KEYINPUT67), .B(n516), .Z(n519) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n517), .Z(n868) );
  NAND2_X1 U573 ( .A1(n868), .A2(G137), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n519), .A2(n518), .ZN(n521) );
  INV_X1 U575 ( .A(KEYINPUT68), .ZN(n520) );
  XNOR2_X1 U576 ( .A(n521), .B(n520), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n527) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n524), .ZN(n865) );
  NAND2_X1 U579 ( .A1(G125), .A2(n865), .ZN(n525) );
  XNOR2_X1 U580 ( .A(KEYINPUT65), .B(n525), .ZN(n526) );
  XOR2_X1 U581 ( .A(G651), .B(KEYINPUT70), .Z(n534) );
  NOR2_X1 U582 ( .A1(G543), .A2(n534), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n528), .Z(n639) );
  NAND2_X1 U584 ( .A1(G63), .A2(n639), .ZN(n530) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n625) );
  NAND2_X1 U586 ( .A1(G51), .A2(n640), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n531), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n532), .B(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U591 ( .A1(G89), .A2(n645), .ZN(n533) );
  XNOR2_X1 U592 ( .A(n533), .B(KEYINPUT4), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n625), .A2(n534), .ZN(n636) );
  NAND2_X1 U594 ( .A1(G76), .A2(n636), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U596 ( .A(KEYINPUT76), .B(n537), .Z(n538) );
  XNOR2_X1 U597 ( .A(KEYINPUT5), .B(n538), .ZN(n539) );
  NOR2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(n541), .Z(G168) );
  XNOR2_X1 U600 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U601 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U602 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  NAND2_X1 U604 ( .A1(G108), .A2(G120), .ZN(n542) );
  NOR2_X1 U605 ( .A1(G237), .A2(n542), .ZN(n543) );
  NAND2_X1 U606 ( .A1(G69), .A2(n543), .ZN(n820) );
  NAND2_X1 U607 ( .A1(n820), .A2(G567), .ZN(n549) );
  NOR2_X1 U608 ( .A1(G219), .A2(G220), .ZN(n544) );
  XNOR2_X1 U609 ( .A(KEYINPUT22), .B(n544), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n545), .A2(G96), .ZN(n546) );
  NOR2_X1 U611 ( .A1(G218), .A2(n546), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT90), .B(n547), .Z(n821) );
  NAND2_X1 U613 ( .A1(n821), .A2(G2106), .ZN(n548) );
  AND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(G319) );
  NAND2_X1 U615 ( .A1(G77), .A2(n636), .ZN(n551) );
  NAND2_X1 U616 ( .A1(G90), .A2(n645), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT9), .B(n552), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G64), .A2(n639), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G52), .A2(n640), .ZN(n553) );
  AND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(G301) );
  INV_X1 U623 ( .A(G301), .ZN(G171) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U625 ( .A1(G135), .A2(n868), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n557), .B(KEYINPUT78), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G123), .A2(n865), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n558), .B(KEYINPUT18), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n864), .A2(G111), .ZN(n559) );
  NAND2_X1 U630 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U631 ( .A1(G99), .A2(n869), .ZN(n561) );
  XNOR2_X1 U632 ( .A(KEYINPUT79), .B(n561), .ZN(n562) );
  NOR2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n939) );
  XNOR2_X1 U635 ( .A(G2096), .B(n939), .ZN(n566) );
  OR2_X1 U636 ( .A1(G2100), .A2(n566), .ZN(G156) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n816) );
  NAND2_X1 U641 ( .A1(n816), .A2(G567), .ZN(n568) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U643 ( .A1(G56), .A2(n639), .ZN(n569) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n569), .Z(n575) );
  NAND2_X1 U645 ( .A1(G81), .A2(n645), .ZN(n570) );
  XNOR2_X1 U646 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U647 ( .A1(G68), .A2(n636), .ZN(n571) );
  NAND2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  NOR2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n640), .A2(G43), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n972) );
  INV_X1 U653 ( .A(G860), .ZN(n605) );
  OR2_X1 U654 ( .A1(n972), .A2(n605), .ZN(G153) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G66), .A2(n639), .ZN(n579) );
  NAND2_X1 U657 ( .A1(G92), .A2(n645), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n584) );
  NAND2_X1 U659 ( .A1(G79), .A2(n636), .ZN(n581) );
  NAND2_X1 U660 ( .A1(G54), .A2(n640), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U662 ( .A(KEYINPUT75), .B(n582), .Z(n583) );
  NOR2_X1 U663 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U664 ( .A(KEYINPUT15), .B(n585), .Z(n963) );
  OR2_X1 U665 ( .A1(n963), .A2(G868), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G53), .A2(n640), .ZN(n588) );
  XNOR2_X1 U668 ( .A(n588), .B(KEYINPUT72), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G78), .A2(n636), .ZN(n590) );
  NAND2_X1 U670 ( .A1(G65), .A2(n639), .ZN(n589) );
  NAND2_X1 U671 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U672 ( .A1(G91), .A2(n645), .ZN(n591) );
  XNOR2_X1 U673 ( .A(KEYINPUT71), .B(n591), .ZN(n592) );
  NOR2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n595), .A2(n594), .ZN(G299) );
  XNOR2_X1 U676 ( .A(KEYINPUT77), .B(G868), .ZN(n596) );
  NOR2_X1 U677 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U679 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n605), .A2(G559), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n599), .A2(n963), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n972), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n963), .A2(G868), .ZN(n601) );
  NOR2_X1 U685 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G559), .A2(n963), .ZN(n604) );
  XOR2_X1 U688 ( .A(n972), .B(n604), .Z(n658) );
  NAND2_X1 U689 ( .A1(n605), .A2(n658), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G80), .A2(n636), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n606), .B(KEYINPUT80), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n640), .A2(G55), .ZN(n608) );
  NAND2_X1 U693 ( .A1(G93), .A2(n645), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U695 ( .A1(G67), .A2(n639), .ZN(n609) );
  XNOR2_X1 U696 ( .A(KEYINPUT81), .B(n609), .ZN(n610) );
  NOR2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n656) );
  XNOR2_X1 U699 ( .A(n614), .B(n656), .ZN(G145) );
  NAND2_X1 U700 ( .A1(G72), .A2(n636), .ZN(n616) );
  NAND2_X1 U701 ( .A1(G60), .A2(n639), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U703 ( .A1(G85), .A2(n645), .ZN(n617) );
  XNOR2_X1 U704 ( .A(KEYINPUT69), .B(n617), .ZN(n618) );
  NOR2_X1 U705 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n640), .A2(G47), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n621), .A2(n620), .ZN(G290) );
  NAND2_X1 U708 ( .A1(G49), .A2(n640), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U711 ( .A1(n639), .A2(n624), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n625), .A2(G87), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G50), .A2(n640), .ZN(n628) );
  XNOR2_X1 U715 ( .A(n628), .B(KEYINPUT84), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G75), .A2(n636), .ZN(n630) );
  NAND2_X1 U717 ( .A1(G62), .A2(n639), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U719 ( .A1(G88), .A2(n645), .ZN(n631) );
  XNOR2_X1 U720 ( .A(KEYINPUT85), .B(n631), .ZN(n632) );
  NOR2_X1 U721 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  XOR2_X1 U724 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n638) );
  NAND2_X1 U725 ( .A1(G73), .A2(n636), .ZN(n637) );
  XNOR2_X1 U726 ( .A(n638), .B(n637), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G61), .A2(n639), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G48), .A2(n640), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G86), .A2(n645), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U733 ( .A(KEYINPUT83), .B(n648), .Z(G305) );
  INV_X1 U734 ( .A(G868), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n649), .A2(n656), .ZN(n650) );
  XNOR2_X1 U736 ( .A(n650), .B(KEYINPUT88), .ZN(n662) );
  XOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n651) );
  XNOR2_X1 U738 ( .A(G288), .B(n651), .ZN(n652) );
  XNOR2_X1 U739 ( .A(G290), .B(n652), .ZN(n654) );
  INV_X1 U740 ( .A(G299), .ZN(n965) );
  XNOR2_X1 U741 ( .A(n965), .B(G166), .ZN(n653) );
  XNOR2_X1 U742 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U743 ( .A(n655), .B(G305), .ZN(n657) );
  XNOR2_X1 U744 ( .A(n657), .B(n656), .ZN(n881) );
  XNOR2_X1 U745 ( .A(n881), .B(n658), .ZN(n659) );
  XNOR2_X1 U746 ( .A(n659), .B(KEYINPUT87), .ZN(n660) );
  NAND2_X1 U747 ( .A1(G868), .A2(n660), .ZN(n661) );
  NAND2_X1 U748 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XNOR2_X1 U750 ( .A(n663), .B(KEYINPUT89), .ZN(n664) );
  XNOR2_X1 U751 ( .A(n664), .B(KEYINPUT20), .ZN(n665) );
  NAND2_X1 U752 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n667), .A2(G2072), .ZN(G158) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n668) );
  XNOR2_X1 U756 ( .A(KEYINPUT91), .B(n668), .ZN(n669) );
  NAND2_X1 U757 ( .A1(n669), .A2(G319), .ZN(n670) );
  XOR2_X1 U758 ( .A(KEYINPUT92), .B(n670), .Z(n819) );
  NAND2_X1 U759 ( .A1(G36), .A2(n819), .ZN(G176) );
  NAND2_X1 U760 ( .A1(G138), .A2(n868), .ZN(n672) );
  NAND2_X1 U761 ( .A1(G102), .A2(n869), .ZN(n671) );
  NAND2_X1 U762 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U763 ( .A1(G114), .A2(n864), .ZN(n674) );
  NAND2_X1 U764 ( .A1(G126), .A2(n865), .ZN(n673) );
  NAND2_X1 U765 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U766 ( .A1(n676), .A2(n675), .ZN(G164) );
  XOR2_X1 U767 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n763) );
  INV_X1 U769 ( .A(n763), .ZN(n677) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n764) );
  NOR2_X1 U771 ( .A1(G1966), .A2(n762), .ZN(n736) );
  NOR2_X1 U772 ( .A1(G2084), .A2(n721), .ZN(n735) );
  NOR2_X1 U773 ( .A1(n736), .A2(n735), .ZN(n678) );
  NAND2_X1 U774 ( .A1(G8), .A2(n678), .ZN(n679) );
  XNOR2_X1 U775 ( .A(KEYINPUT30), .B(n679), .ZN(n681) );
  INV_X1 U776 ( .A(KEYINPUT101), .ZN(n680) );
  XNOR2_X1 U777 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U778 ( .A1(n682), .A2(G168), .ZN(n687) );
  INV_X1 U779 ( .A(n721), .ZN(n705) );
  NOR2_X1 U780 ( .A1(n705), .A2(G1961), .ZN(n683) );
  XOR2_X1 U781 ( .A(KEYINPUT96), .B(n683), .Z(n685) );
  XNOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .ZN(n914) );
  NAND2_X1 U783 ( .A1(n705), .A2(n914), .ZN(n684) );
  NAND2_X1 U784 ( .A1(n685), .A2(n684), .ZN(n718) );
  NOR2_X1 U785 ( .A1(G171), .A2(n718), .ZN(n686) );
  NOR2_X1 U786 ( .A1(n687), .A2(n686), .ZN(n690) );
  XOR2_X1 U787 ( .A(G1996), .B(KEYINPUT98), .Z(n905) );
  NOR2_X1 U788 ( .A1(n721), .A2(n905), .ZN(n692) );
  XNOR2_X1 U789 ( .A(KEYINPUT26), .B(KEYINPUT99), .ZN(n691) );
  XNOR2_X1 U790 ( .A(n692), .B(n691), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n721), .A2(G1341), .ZN(n693) );
  NAND2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n963), .A2(n701), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n721), .A2(G1348), .ZN(n696) );
  XNOR2_X1 U795 ( .A(n696), .B(KEYINPUT100), .ZN(n698) );
  NAND2_X1 U796 ( .A1(n705), .A2(G2067), .ZN(n697) );
  NAND2_X1 U797 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U798 ( .A1(n700), .A2(n699), .ZN(n703) );
  OR2_X1 U799 ( .A1(n963), .A2(n701), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n710) );
  NAND2_X1 U801 ( .A1(G1956), .A2(n721), .ZN(n704) );
  XNOR2_X1 U802 ( .A(KEYINPUT97), .B(n704), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n705), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U804 ( .A(n706), .B(KEYINPUT27), .ZN(n707) );
  NOR2_X1 U805 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n965), .A2(n711), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n965), .A2(n711), .ZN(n713) );
  XNOR2_X1 U809 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n718), .A2(G171), .ZN(n719) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n762), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n721), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n724), .A2(G303), .ZN(n726) );
  AND2_X1 U816 ( .A1(n733), .A2(n726), .ZN(n725) );
  NAND2_X1 U817 ( .A1(n734), .A2(n725), .ZN(n730) );
  INV_X1 U818 ( .A(n726), .ZN(n727) );
  OR2_X1 U819 ( .A1(n727), .A2(G286), .ZN(n728) );
  AND2_X1 U820 ( .A1(n728), .A2(G8), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n732) );
  XOR2_X1 U822 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n731) );
  XNOR2_X1 U823 ( .A(n732), .B(n731), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n738) );
  AND2_X1 U825 ( .A1(G8), .A2(n735), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n513), .ZN(n753) );
  NAND2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n961) );
  AND2_X1 U828 ( .A1(n753), .A2(n961), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n752), .A2(n739), .ZN(n743) );
  INV_X1 U830 ( .A(n961), .ZN(n741) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n964) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NOR2_X1 U833 ( .A1(n964), .A2(n960), .ZN(n740) );
  OR2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  AND2_X1 U835 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n762), .A2(n744), .ZN(n745) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n745), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n964), .A2(KEYINPUT33), .ZN(n746) );
  NOR2_X1 U839 ( .A1(n746), .A2(n762), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n982), .A2(n749), .ZN(n758) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n750) );
  NAND2_X1 U842 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT104), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n756), .A2(n762), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U848 ( .A(KEYINPUT105), .B(n759), .ZN(n804) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XOR2_X1 U850 ( .A(n760), .B(KEYINPUT24), .Z(n761) );
  NOR2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n802) );
  NOR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n807) );
  NAND2_X1 U853 ( .A1(G105), .A2(n869), .ZN(n765) );
  XNOR2_X1 U854 ( .A(n765), .B(KEYINPUT38), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G141), .A2(n868), .ZN(n767) );
  NAND2_X1 U856 ( .A1(G129), .A2(n865), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U858 ( .A1(G117), .A2(n864), .ZN(n768) );
  XNOR2_X1 U859 ( .A(KEYINPUT95), .B(n768), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n875) );
  NOR2_X1 U862 ( .A1(G1996), .A2(n875), .ZN(n933) );
  NAND2_X1 U863 ( .A1(n875), .A2(G1996), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G131), .A2(n868), .ZN(n774) );
  NAND2_X1 U865 ( .A1(G119), .A2(n865), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G107), .A2(n864), .ZN(n776) );
  NAND2_X1 U868 ( .A1(G95), .A2(n869), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U871 ( .A(KEYINPUT94), .B(n779), .Z(n859) );
  NAND2_X1 U872 ( .A1(n859), .A2(G1991), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n937) );
  NAND2_X1 U874 ( .A1(n937), .A2(n807), .ZN(n806) );
  INV_X1 U875 ( .A(n806), .ZN(n784) );
  NOR2_X1 U876 ( .A1(G1986), .A2(G290), .ZN(n782) );
  NOR2_X1 U877 ( .A1(G1991), .A2(n859), .ZN(n942) );
  NOR2_X1 U878 ( .A1(n782), .A2(n942), .ZN(n783) );
  NOR2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U880 ( .A1(n933), .A2(n785), .ZN(n786) );
  XNOR2_X1 U881 ( .A(KEYINPUT39), .B(n786), .ZN(n797) );
  NAND2_X1 U882 ( .A1(n868), .A2(G140), .ZN(n787) );
  XOR2_X1 U883 ( .A(KEYINPUT93), .B(n787), .Z(n789) );
  NAND2_X1 U884 ( .A1(n869), .A2(G104), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G116), .A2(n864), .ZN(n792) );
  NAND2_X1 U888 ( .A1(G128), .A2(n865), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U892 ( .A(KEYINPUT36), .B(n796), .ZN(n858) );
  XNOR2_X1 U893 ( .A(G2067), .B(KEYINPUT37), .ZN(n798) );
  NOR2_X1 U894 ( .A1(n858), .A2(n798), .ZN(n950) );
  NAND2_X1 U895 ( .A1(n807), .A2(n950), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n797), .A2(n805), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n858), .A2(n798), .ZN(n947) );
  NAND2_X1 U898 ( .A1(n799), .A2(n947), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n807), .A2(n800), .ZN(n801) );
  XOR2_X1 U900 ( .A(KEYINPUT106), .B(n801), .Z(n811) );
  NOR2_X1 U901 ( .A1(n802), .A2(n811), .ZN(n803) );
  AND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n809) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n969) );
  AND2_X1 U905 ( .A1(n969), .A2(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n815) );
  XOR2_X1 U909 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U913 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(G188) );
  XNOR2_X1 U916 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G108), .ZN(G238) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  XOR2_X1 U923 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n823) );
  XNOR2_X1 U924 ( .A(G2678), .B(KEYINPUT43), .ZN(n822) );
  XNOR2_X1 U925 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U926 ( .A(KEYINPUT42), .B(G2090), .Z(n825) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2072), .ZN(n824) );
  XNOR2_X1 U928 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U929 ( .A(n827), .B(n826), .Z(n829) );
  XNOR2_X1 U930 ( .A(G2096), .B(G2100), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n831) );
  XOR2_X1 U932 ( .A(G2084), .B(G2078), .Z(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1976), .B(G1971), .Z(n833) );
  XNOR2_X1 U935 ( .A(G1966), .B(G1961), .ZN(n832) );
  XNOR2_X1 U936 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U937 ( .A(n834), .B(G2474), .Z(n836) );
  XNOR2_X1 U938 ( .A(G1981), .B(G1956), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1986), .Z(n838) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(G229) );
  NAND2_X1 U944 ( .A1(G124), .A2(n865), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U946 ( .A1(n864), .A2(G112), .ZN(n842) );
  NAND2_X1 U947 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G136), .A2(n868), .ZN(n845) );
  NAND2_X1 U949 ( .A1(G100), .A2(n869), .ZN(n844) );
  NAND2_X1 U950 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U951 ( .A1(n847), .A2(n846), .ZN(G162) );
  XNOR2_X1 U952 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n849) );
  XNOR2_X1 U953 ( .A(n939), .B(KEYINPUT112), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U955 ( .A(G164), .B(n850), .ZN(n863) );
  NAND2_X1 U956 ( .A1(G139), .A2(n868), .ZN(n852) );
  NAND2_X1 U957 ( .A1(G103), .A2(n869), .ZN(n851) );
  NAND2_X1 U958 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G115), .A2(n864), .ZN(n854) );
  NAND2_X1 U960 ( .A1(G127), .A2(n865), .ZN(n853) );
  NAND2_X1 U961 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U962 ( .A(KEYINPUT47), .B(n855), .Z(n856) );
  NOR2_X1 U963 ( .A1(n857), .A2(n856), .ZN(n925) );
  XNOR2_X1 U964 ( .A(n858), .B(n925), .ZN(n861) );
  XNOR2_X1 U965 ( .A(G160), .B(n859), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n879) );
  NAND2_X1 U968 ( .A1(G118), .A2(n864), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G130), .A2(n865), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G142), .A2(n868), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G106), .A2(n869), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(G162), .B(n877), .Z(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U979 ( .A1(G37), .A2(n880), .ZN(G395) );
  XOR2_X1 U980 ( .A(n881), .B(G286), .Z(n883) );
  XNOR2_X1 U981 ( .A(G171), .B(n963), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n884), .B(n972), .ZN(n885) );
  NOR2_X1 U984 ( .A1(G37), .A2(n885), .ZN(G397) );
  XOR2_X1 U985 ( .A(G2451), .B(G2443), .Z(n887) );
  XNOR2_X1 U986 ( .A(G2427), .B(G2454), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(n888), .B(G2446), .Z(n890) );
  XNOR2_X1 U989 ( .A(G1341), .B(G1348), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U991 ( .A(G2435), .B(KEYINPUT108), .Z(n892) );
  XNOR2_X1 U992 ( .A(G2430), .B(G2438), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(n894), .B(n893), .Z(n895) );
  NAND2_X1 U995 ( .A1(G14), .A2(n895), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G319), .A2(n902), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n896) );
  XOR2_X1 U998 ( .A(KEYINPUT49), .B(n896), .Z(n897) );
  XNOR2_X1 U999 ( .A(n897), .B(KEYINPUT113), .ZN(n898) );
  NOR2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n901) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(n902), .ZN(G401) );
  XNOR2_X1 U1005 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n903) );
  XNOR2_X1 U1006 ( .A(n903), .B(G34), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(G2084), .B(n904), .ZN(n921) );
  XNOR2_X1 U1008 ( .A(G2090), .B(G35), .ZN(n919) );
  XNOR2_X1 U1009 ( .A(n905), .B(G32), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(G2072), .B(G33), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(G25), .B(G1991), .ZN(n906) );
  NOR2_X1 U1012 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1013 ( .A1(G28), .A2(n908), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(KEYINPUT118), .B(G2067), .ZN(n909) );
  XNOR2_X1 U1015 ( .A(G26), .B(n909), .ZN(n910) );
  NOR2_X1 U1016 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n916) );
  XOR2_X1 U1018 ( .A(G27), .B(n914), .Z(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1020 ( .A(KEYINPUT53), .B(n917), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(G29), .A2(KEYINPUT55), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n922), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(G11), .A2(n923), .ZN(n958) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n952) );
  OR2_X1 U1027 ( .A1(n952), .A2(n924), .ZN(n956) );
  XNOR2_X1 U1028 ( .A(G164), .B(G2078), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n925), .ZN(n926) );
  XNOR2_X1 U1030 ( .A(n926), .B(KEYINPUT116), .ZN(n927) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(n929), .B(KEYINPUT50), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(KEYINPUT117), .B(n930), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G162), .ZN(n931) );
  XNOR2_X1 U1035 ( .A(n931), .B(KEYINPUT115), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n934), .Z(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n946) );
  INV_X1 U1039 ( .A(n937), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(G160), .B(G2084), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n938), .B(KEYINPUT114), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(n951), .B(KEYINPUT52), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(G29), .A2(n954), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n1017) );
  XOR2_X1 U1053 ( .A(G1961), .B(G171), .Z(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n978) );
  XNOR2_X1 U1056 ( .A(n963), .B(G1348), .ZN(n976) );
  XOR2_X1 U1057 ( .A(n964), .B(KEYINPUT122), .Z(n967) );
  XNOR2_X1 U1058 ( .A(n965), .B(G1956), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G1341), .B(n972), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(KEYINPUT123), .B(n979), .ZN(n986) );
  XOR2_X1 U1068 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n984) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n980), .B(KEYINPUT120), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1072 ( .A(n984), .B(n983), .Z(n985) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .Z(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(n989), .ZN(n1014) );
  XNOR2_X1 U1077 ( .A(G1348), .B(KEYINPUT59), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n990), .B(G4), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(G1981), .B(G6), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G19), .B(G1341), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G20), .B(G1956), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1085 ( .A(KEYINPUT60), .B(n997), .Z(n999) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G21), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT126), .B(n1000), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G5), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1001), .B(KEYINPUT125), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G24), .B(G1986), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(G1976), .B(G23), .Z(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1011), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(G16), .A2(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1015), .Z(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

