

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n655), .A2(n654), .ZN(n671) );
  NOR2_X1 U550 ( .A1(G651), .A2(n568), .ZN(n799) );
  BUF_X1 U551 ( .A(n688), .Z(n689) );
  NOR2_X2 U552 ( .A1(G164), .A2(G1384), .ZN(n684) );
  AND2_X1 U553 ( .A1(n725), .A2(n514), .ZN(n675) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(n674), .ZN(n514) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n637) );
  INV_X1 U556 ( .A(n998), .ZN(n718) );
  AND2_X1 U557 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U558 ( .A(n591), .B(KEYINPUT73), .ZN(n595) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  XOR2_X1 U560 ( .A(G543), .B(KEYINPUT0), .Z(n536) );
  OR2_X1 U561 ( .A1(n539), .A2(n568), .ZN(n540) );
  INV_X1 U562 ( .A(KEYINPUT15), .ZN(n610) );
  NAND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XNOR2_X1 U564 ( .A(n515), .B(KEYINPUT67), .ZN(n890) );
  NAND2_X1 U565 ( .A1(n890), .A2(G114), .ZN(n519) );
  XOR2_X1 U566 ( .A(KEYINPUT68), .B(n516), .Z(n517) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(n517), .ZN(n688) );
  NAND2_X1 U568 ( .A1(G138), .A2(n688), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n519), .A2(n518), .ZN(n525) );
  XNOR2_X1 U570 ( .A(KEYINPUT65), .B(G2104), .ZN(n521) );
  AND2_X1 U571 ( .A1(n521), .A2(G2105), .ZN(n520) );
  XNOR2_X1 U572 ( .A(KEYINPUT66), .B(n520), .ZN(n530) );
  BUF_X1 U573 ( .A(n530), .Z(n891) );
  NAND2_X1 U574 ( .A1(G126), .A2(n891), .ZN(n523) );
  NOR2_X1 U575 ( .A1(G2105), .A2(n521), .ZN(n526) );
  BUF_X1 U576 ( .A(n526), .Z(n894) );
  NAND2_X1 U577 ( .A1(n894), .A2(G102), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U579 ( .A1(n525), .A2(n524), .ZN(G164) );
  NAND2_X1 U580 ( .A1(G137), .A2(n688), .ZN(n529) );
  NAND2_X1 U581 ( .A1(G101), .A2(n526), .ZN(n527) );
  XOR2_X1 U582 ( .A(KEYINPUT23), .B(n527), .Z(n528) );
  NAND2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G113), .A2(n890), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G125), .A2(n530), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U587 ( .A1(n534), .A2(n533), .ZN(G160) );
  INV_X1 U588 ( .A(G651), .ZN(n539) );
  NOR2_X1 U589 ( .A1(G543), .A2(n539), .ZN(n535) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n535), .Z(n794) );
  NAND2_X1 U591 ( .A1(G64), .A2(n794), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT69), .B(n536), .Z(n568) );
  NAND2_X1 U593 ( .A1(G52), .A2(n799), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n796) );
  NAND2_X1 U596 ( .A1(G90), .A2(n796), .ZN(n542) );
  XOR2_X2 U597 ( .A(KEYINPUT70), .B(n540), .Z(n800) );
  NAND2_X1 U598 ( .A1(G77), .A2(n800), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U601 ( .A1(n545), .A2(n544), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G63), .A2(n794), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G51), .A2(n799), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT6), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n549), .B(KEYINPUT79), .ZN(n556) );
  XNOR2_X1 U607 ( .A(KEYINPUT5), .B(KEYINPUT78), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n796), .A2(G89), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G76), .A2(n800), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n554), .B(n553), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  NAND2_X1 U615 ( .A1(G88), .A2(n796), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G75), .A2(n800), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G62), .A2(n794), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G50), .A2(n799), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G166) );
  INV_X1 U622 ( .A(G166), .ZN(G303) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT80), .B(n564), .ZN(G286) );
  NAND2_X1 U625 ( .A1(G49), .A2(n799), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U628 ( .A1(n794), .A2(n567), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G87), .A2(n568), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT87), .B(n569), .Z(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(G288) );
  AND2_X1 U632 ( .A1(G72), .A2(n800), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G85), .A2(n796), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G47), .A2(n799), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n794), .A2(G60), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(G290) );
  NAND2_X1 U639 ( .A1(n800), .A2(G73), .ZN(n578) );
  XNOR2_X1 U640 ( .A(n578), .B(KEYINPUT2), .ZN(n585) );
  NAND2_X1 U641 ( .A1(G86), .A2(n796), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G61), .A2(n794), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n799), .A2(G48), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT88), .B(n581), .Z(n582) );
  NOR2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(G305) );
  NAND2_X1 U648 ( .A1(G40), .A2(G160), .ZN(n586) );
  XNOR2_X1 U649 ( .A(n586), .B(KEYINPUT93), .ZN(n682) );
  NAND2_X2 U650 ( .A1(n684), .A2(n682), .ZN(n656) );
  NAND2_X1 U651 ( .A1(G8), .A2(n656), .ZN(n729) );
  INV_X1 U652 ( .A(G1996), .ZN(n945) );
  NOR2_X1 U653 ( .A1(n656), .A2(n945), .ZN(n588) );
  XOR2_X1 U654 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n587) );
  XNOR2_X1 U655 ( .A(n588), .B(n587), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n656), .A2(G1341), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n616) );
  NAND2_X1 U658 ( .A1(G68), .A2(n800), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT72), .B(KEYINPUT12), .Z(n593) );
  NAND2_X1 U660 ( .A1(G81), .A2(n796), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n593), .B(n592), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U663 ( .A(KEYINPUT13), .B(KEYINPUT74), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n597), .B(n596), .ZN(n602) );
  NAND2_X1 U665 ( .A1(n794), .A2(G56), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT14), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G43), .A2(n799), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n995) );
  NAND2_X1 U670 ( .A1(n799), .A2(G54), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G79), .A2(n800), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U673 ( .A(KEYINPUT77), .B(n605), .Z(n609) );
  NAND2_X1 U674 ( .A1(G92), .A2(n796), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G66), .A2(n794), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  OR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  XNOR2_X2 U678 ( .A(n611), .B(n610), .ZN(n996) );
  NAND2_X1 U679 ( .A1(G1348), .A2(n656), .ZN(n613) );
  INV_X1 U680 ( .A(n656), .ZN(n639) );
  NAND2_X1 U681 ( .A1(G2067), .A2(n639), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n996), .A2(n617), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n995), .A2(n614), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n619) );
  NOR2_X1 U686 ( .A1(n617), .A2(n996), .ZN(n618) );
  NOR2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n632) );
  XNOR2_X1 U688 ( .A(KEYINPUT98), .B(G1956), .ZN(n929) );
  NAND2_X1 U689 ( .A1(n656), .A2(n929), .ZN(n623) );
  INV_X1 U690 ( .A(n656), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n620), .A2(G2072), .ZN(n621) );
  XOR2_X1 U692 ( .A(KEYINPUT27), .B(n621), .Z(n622) );
  NAND2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n624), .B(KEYINPUT99), .ZN(n633) );
  NAND2_X1 U695 ( .A1(G65), .A2(n794), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G53), .A2(n799), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G91), .A2(n796), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G78), .A2(n800), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n1012) );
  NAND2_X1 U702 ( .A1(n633), .A2(n1012), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n633), .A2(n1012), .ZN(n634) );
  XOR2_X1 U705 ( .A(n634), .B(KEYINPUT28), .Z(n635) );
  NAND2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n638), .B(n637), .ZN(n643) );
  INV_X1 U708 ( .A(G1961), .ZN(n918) );
  NAND2_X1 U709 ( .A1(n656), .A2(n918), .ZN(n641) );
  XNOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U711 ( .A1(n639), .A2(n944), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n647) );
  NAND2_X1 U713 ( .A1(n647), .A2(G171), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n664) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n729), .ZN(n652) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n656), .ZN(n651) );
  NOR2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G8), .A2(n644), .ZN(n645) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n645), .ZN(n646) );
  NOR2_X1 U720 ( .A1(G168), .A2(n646), .ZN(n649) );
  NOR2_X1 U721 ( .A1(G171), .A2(n647), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U723 ( .A(KEYINPUT31), .B(n650), .Z(n662) );
  AND2_X1 U724 ( .A1(n664), .A2(n662), .ZN(n655) );
  AND2_X1 U725 ( .A1(G8), .A2(n651), .ZN(n653) );
  OR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n654) );
  INV_X1 U727 ( .A(G8), .ZN(n661) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n729), .ZN(n658) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n656), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n659), .A2(G303), .ZN(n660) );
  OR2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n665) );
  AND2_X1 U733 ( .A1(n662), .A2(n665), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n668) );
  INV_X1 U735 ( .A(n665), .ZN(n666) );
  OR2_X1 U736 ( .A1(n666), .A2(G286), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT32), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n725) );
  NOR2_X1 U740 ( .A1(G288), .A2(G1976), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT100), .ZN(n1007) );
  NOR2_X1 U742 ( .A1(G1971), .A2(G303), .ZN(n1014) );
  XOR2_X1 U743 ( .A(n1014), .B(KEYINPUT101), .Z(n673) );
  NOR2_X1 U744 ( .A1(n1007), .A2(n673), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(KEYINPUT103), .ZN(n676) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  NAND2_X1 U747 ( .A1(n676), .A2(n1005), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT104), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n729), .A2(n678), .ZN(n679) );
  OR2_X2 U750 ( .A1(n679), .A2(KEYINPUT33), .ZN(n721) );
  INV_X1 U751 ( .A(n1007), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n729), .A2(n680), .ZN(n681) );
  NAND2_X1 U753 ( .A1(KEYINPUT33), .A2(n681), .ZN(n707) );
  XNOR2_X1 U754 ( .A(G1986), .B(G290), .ZN(n1006) );
  INV_X1 U755 ( .A(n682), .ZN(n683) );
  NOR2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n751) );
  NAND2_X1 U757 ( .A1(n1006), .A2(n751), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n685), .B(KEYINPUT94), .ZN(n706) );
  XOR2_X1 U759 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n687) );
  NAND2_X1 U760 ( .A1(G105), .A2(n894), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n687), .B(n686), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n890), .A2(G117), .ZN(n691) );
  NAND2_X1 U763 ( .A1(G141), .A2(n689), .ZN(n690) );
  NAND2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U766 ( .A1(G129), .A2(n891), .ZN(n694) );
  NAND2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n883) );
  NAND2_X1 U768 ( .A1(G1996), .A2(n883), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n894), .A2(G95), .ZN(n697) );
  NAND2_X1 U770 ( .A1(G131), .A2(n689), .ZN(n696) );
  NAND2_X1 U771 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U772 ( .A(KEYINPUT95), .B(n698), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n891), .A2(G119), .ZN(n700) );
  NAND2_X1 U774 ( .A1(G107), .A2(n890), .ZN(n699) );
  AND2_X1 U775 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U776 ( .A1(n702), .A2(n701), .ZN(n885) );
  NAND2_X1 U777 ( .A1(G1991), .A2(n885), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n974) );
  NAND2_X1 U779 ( .A1(n974), .A2(n751), .ZN(n705) );
  XOR2_X1 U780 ( .A(KEYINPUT97), .B(n705), .Z(n739) );
  AND2_X1 U781 ( .A1(n706), .A2(n739), .ZN(n733) );
  AND2_X1 U782 ( .A1(n707), .A2(n733), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n894), .A2(G104), .ZN(n709) );
  NAND2_X1 U784 ( .A1(G140), .A2(n689), .ZN(n708) );
  NAND2_X1 U785 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U786 ( .A(KEYINPUT34), .B(n710), .ZN(n715) );
  NAND2_X1 U787 ( .A1(G116), .A2(n890), .ZN(n712) );
  NAND2_X1 U788 ( .A1(G128), .A2(n891), .ZN(n711) );
  NAND2_X1 U789 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U790 ( .A(KEYINPUT35), .B(n713), .Z(n714) );
  NOR2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U792 ( .A(KEYINPUT36), .B(n716), .ZN(n903) );
  XNOR2_X1 U793 ( .A(KEYINPUT37), .B(G2067), .ZN(n748) );
  NOR2_X1 U794 ( .A1(n903), .A2(n748), .ZN(n965) );
  NAND2_X1 U795 ( .A1(n751), .A2(n965), .ZN(n746) );
  AND2_X1 U796 ( .A1(n717), .A2(n746), .ZN(n719) );
  XNOR2_X1 U797 ( .A(G1981), .B(G305), .ZN(n998) );
  NAND2_X1 U798 ( .A1(n721), .A2(n720), .ZN(n737) );
  INV_X1 U799 ( .A(n746), .ZN(n735) );
  NAND2_X1 U800 ( .A1(G8), .A2(G166), .ZN(n722) );
  NOR2_X1 U801 ( .A1(G2090), .A2(n722), .ZN(n723) );
  XNOR2_X1 U802 ( .A(KEYINPUT105), .B(n723), .ZN(n724) );
  NAND2_X1 U803 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U804 ( .A1(n726), .A2(n729), .ZN(n731) );
  NOR2_X1 U805 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U806 ( .A(n727), .B(KEYINPUT24), .Z(n728) );
  OR2_X1 U807 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U808 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U812 ( .A(n738), .B(KEYINPUT106), .ZN(n753) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n883), .ZN(n983) );
  INV_X1 U814 ( .A(n739), .ZN(n742) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n885), .ZN(n975) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U817 ( .A1(n975), .A2(n740), .ZN(n741) );
  NOR2_X1 U818 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U819 ( .A(KEYINPUT107), .B(n743), .Z(n744) );
  NOR2_X1 U820 ( .A1(n983), .A2(n744), .ZN(n745) );
  XNOR2_X1 U821 ( .A(n745), .B(KEYINPUT39), .ZN(n747) );
  NAND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U823 ( .A1(n903), .A2(n748), .ZN(n964) );
  NAND2_X1 U824 ( .A1(n749), .A2(n964), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U827 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n754) );
  XNOR2_X1 U828 ( .A(n755), .B(n754), .ZN(G329) );
  XOR2_X1 U829 ( .A(G2430), .B(G2443), .Z(n757) );
  XNOR2_X1 U830 ( .A(KEYINPUT109), .B(G2451), .ZN(n756) );
  XNOR2_X1 U831 ( .A(n757), .B(n756), .ZN(n764) );
  XOR2_X1 U832 ( .A(G2435), .B(G2427), .Z(n759) );
  XNOR2_X1 U833 ( .A(G2446), .B(G2454), .ZN(n758) );
  XNOR2_X1 U834 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U835 ( .A(n760), .B(G2438), .Z(n762) );
  XNOR2_X1 U836 ( .A(G1348), .B(G1341), .ZN(n761) );
  XNOR2_X1 U837 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n764), .B(n763), .ZN(n765) );
  AND2_X1 U839 ( .A1(n765), .A2(G14), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U841 ( .A(n995), .ZN(n792) );
  XNOR2_X1 U842 ( .A(G860), .B(KEYINPUT75), .ZN(n772) );
  OR2_X1 U843 ( .A1(n792), .A2(n772), .ZN(G153) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  INV_X1 U846 ( .A(G108), .ZN(G238) );
  INV_X1 U847 ( .A(G120), .ZN(G236) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U850 ( .A(n766), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U851 ( .A(G567), .ZN(n825) );
  NOR2_X1 U852 ( .A1(n825), .A2(G223), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U854 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n769) );
  INV_X1 U856 ( .A(G868), .ZN(n815) );
  NAND2_X1 U857 ( .A1(n996), .A2(n815), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(G284) );
  XNOR2_X1 U859 ( .A(n1012), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U860 ( .A1(G868), .A2(G286), .ZN(n771) );
  NAND2_X1 U861 ( .A1(G299), .A2(n815), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n772), .A2(G559), .ZN(n773) );
  INV_X1 U864 ( .A(n996), .ZN(n791) );
  NAND2_X1 U865 ( .A1(n773), .A2(n791), .ZN(n774) );
  XNOR2_X1 U866 ( .A(n774), .B(KEYINPUT81), .ZN(n775) );
  XOR2_X1 U867 ( .A(KEYINPUT16), .B(n775), .Z(G148) );
  NAND2_X1 U868 ( .A1(n791), .A2(G868), .ZN(n776) );
  NOR2_X1 U869 ( .A1(G559), .A2(n776), .ZN(n777) );
  XNOR2_X1 U870 ( .A(n777), .B(KEYINPUT82), .ZN(n779) );
  NOR2_X1 U871 ( .A1(n792), .A2(G868), .ZN(n778) );
  NOR2_X1 U872 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U873 ( .A1(G99), .A2(n894), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n890), .A2(G111), .ZN(n781) );
  NAND2_X1 U875 ( .A1(G135), .A2(n689), .ZN(n780) );
  NAND2_X1 U876 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n891), .A2(G123), .ZN(n782) );
  XOR2_X1 U878 ( .A(KEYINPUT18), .B(n782), .Z(n783) );
  NOR2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U881 ( .A(n787), .B(KEYINPUT83), .ZN(n973) );
  XOR2_X1 U882 ( .A(n973), .B(G2096), .Z(n789) );
  XNOR2_X1 U883 ( .A(G2100), .B(KEYINPUT84), .ZN(n788) );
  NOR2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U885 ( .A(KEYINPUT85), .B(n790), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G559), .A2(n791), .ZN(n793) );
  XNOR2_X1 U887 ( .A(n793), .B(n792), .ZN(n812) );
  NOR2_X1 U888 ( .A1(n812), .A2(G860), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G67), .A2(n794), .ZN(n795) );
  XNOR2_X1 U890 ( .A(n795), .B(KEYINPUT86), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n796), .A2(G93), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n799), .A2(G55), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G80), .A2(n800), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n814) );
  XOR2_X1 U897 ( .A(n805), .B(n814), .Z(G145) );
  XOR2_X1 U898 ( .A(KEYINPUT19), .B(KEYINPUT89), .Z(n806) );
  XNOR2_X1 U899 ( .A(G288), .B(n806), .ZN(n809) );
  XNOR2_X1 U900 ( .A(G166), .B(G290), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(G299), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n809), .B(n808), .ZN(n811) );
  XOR2_X1 U903 ( .A(G305), .B(n814), .Z(n810) );
  XNOR2_X1 U904 ( .A(n811), .B(n810), .ZN(n909) );
  XOR2_X1 U905 ( .A(n812), .B(n909), .Z(n813) );
  NAND2_X1 U906 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(G295) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(KEYINPUT90), .Z(n819) );
  NAND2_X1 U910 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n820), .ZN(n821) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G236), .A2(G238), .ZN(n823) );
  NAND2_X1 U917 ( .A1(G69), .A2(n823), .ZN(n824) );
  NOR2_X1 U918 ( .A1(G237), .A2(n824), .ZN(n841) );
  NOR2_X1 U919 ( .A1(n841), .A2(n825), .ZN(n832) );
  NOR2_X1 U920 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U922 ( .A1(G218), .A2(n827), .ZN(n828) );
  XOR2_X1 U923 ( .A(KEYINPUT91), .B(n828), .Z(n829) );
  NAND2_X1 U924 ( .A1(G96), .A2(n829), .ZN(n842) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n842), .ZN(n830) );
  XOR2_X1 U926 ( .A(KEYINPUT92), .B(n830), .Z(n831) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(G319) );
  INV_X1 U928 ( .A(G319), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U932 ( .A(G223), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n835), .A2(G2106), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U936 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U938 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(KEYINPUT111), .B(n840), .Z(G188) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(n841), .ZN(n843) );
  NOR2_X1 U943 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT112), .B(n844), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2084), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n847), .B(G2100), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U953 ( .A(KEYINPUT113), .B(G2678), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U956 ( .A(G1971), .B(G1986), .Z(n855) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n865) );
  XOR2_X1 U959 ( .A(G2474), .B(KEYINPUT41), .Z(n857) );
  XNOR2_X1 U960 ( .A(G1956), .B(KEYINPUT116), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U962 ( .A(G1976), .B(G1981), .Z(n859) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1961), .ZN(n858) );
  XNOR2_X1 U964 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U965 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U966 ( .A(KEYINPUT115), .B(KEYINPUT114), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U969 ( .A1(G112), .A2(n890), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G100), .A2(n894), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n891), .A2(G124), .ZN(n868) );
  XOR2_X1 U973 ( .A(KEYINPUT117), .B(n868), .Z(n869) );
  XNOR2_X1 U974 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G136), .A2(n689), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G115), .A2(n890), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G127), .A2(n891), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n876), .B(KEYINPUT47), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G103), .A2(n894), .ZN(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G139), .A2(n689), .ZN(n879) );
  XNOR2_X1 U985 ( .A(KEYINPUT119), .B(n879), .ZN(n880) );
  NOR2_X1 U986 ( .A1(n881), .A2(n880), .ZN(n967) );
  XOR2_X1 U987 ( .A(G160), .B(n967), .Z(n882) );
  XNOR2_X1 U988 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U989 ( .A(n973), .B(n884), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n885), .B(G162), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n887), .B(n886), .ZN(n905) );
  XOR2_X1 U992 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n889) );
  XNOR2_X1 U993 ( .A(G164), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U994 ( .A(n889), .B(n888), .ZN(n901) );
  NAND2_X1 U995 ( .A1(G118), .A2(n890), .ZN(n893) );
  NAND2_X1 U996 ( .A1(G130), .A2(n891), .ZN(n892) );
  NAND2_X1 U997 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n894), .A2(G106), .ZN(n896) );
  NAND2_X1 U999 ( .A1(G142), .A2(n689), .ZN(n895) );
  NAND2_X1 U1000 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U1001 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U1002 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1003 ( .A(n901), .B(n900), .Z(n902) );
  XOR2_X1 U1004 ( .A(n903), .B(n902), .Z(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(n996), .B(KEYINPUT120), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n995), .B(G171), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n908), .B(n907), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(G286), .B(n909), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n914), .ZN(n915) );
  AND2_X1 U1016 ( .A1(G319), .A2(n915), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1021 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n940) );
  XOR2_X1 U1022 ( .A(G1966), .B(G21), .Z(n920) );
  XNOR2_X1 U1023 ( .A(n918), .B(G5), .ZN(n919) );
  NAND2_X1 U1024 ( .A1(n920), .A2(n919), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(G1971), .B(G22), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(G23), .B(G1976), .ZN(n921) );
  NOR2_X1 U1027 ( .A1(n922), .A2(n921), .ZN(n924) );
  XOR2_X1 U1028 ( .A(G1986), .B(G24), .Z(n923) );
  NAND2_X1 U1029 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1030 ( .A(KEYINPUT58), .B(n925), .ZN(n926) );
  NOR2_X1 U1031 ( .A1(n927), .A2(n926), .ZN(n938) );
  XOR2_X1 U1032 ( .A(G1348), .B(KEYINPUT59), .Z(n928) );
  XNOR2_X1 U1033 ( .A(G4), .B(n928), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(G20), .B(n929), .ZN(n930) );
  NOR2_X1 U1035 ( .A1(n931), .A2(n930), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(G1981), .B(G6), .ZN(n932) );
  NOR2_X1 U1038 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1039 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1040 ( .A(KEYINPUT60), .B(n936), .Z(n937) );
  NAND2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1042 ( .A(n940), .B(n939), .ZN(n941) );
  OR2_X1 U1043 ( .A1(G16), .A2(n941), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(G11), .A2(n942), .ZN(n993) );
  XOR2_X1 U1045 ( .A(G1991), .B(G25), .Z(n943) );
  NAND2_X1 U1046 ( .A1(n943), .A2(G28), .ZN(n950) );
  XOR2_X1 U1047 ( .A(n944), .B(G27), .Z(n947) );
  XOR2_X1 U1048 ( .A(n945), .B(G32), .Z(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1050 ( .A(KEYINPUT124), .B(n948), .Z(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(n955), .B(KEYINPUT53), .ZN(n958) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1060 ( .A(KEYINPUT123), .B(G2090), .Z(n959) );
  XNOR2_X1 U1061 ( .A(G35), .B(n959), .ZN(n960) );
  NOR2_X1 U1062 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1063 ( .A1(G29), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1064 ( .A(n963), .B(KEYINPUT55), .ZN(n991) );
  INV_X1 U1065 ( .A(n964), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(G2072), .B(n967), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(G164), .B(G2078), .ZN(n968) );
  XNOR2_X1 U1069 ( .A(n968), .B(KEYINPUT122), .ZN(n969) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1071 ( .A(n971), .B(KEYINPUT50), .ZN(n979) );
  XOR2_X1 U1072 ( .A(G2084), .B(G160), .Z(n972) );
  NOR2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1080 ( .A(KEYINPUT51), .B(n984), .Z(n985) );
  XNOR2_X1 U1081 ( .A(n985), .B(KEYINPUT121), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1083 ( .A(KEYINPUT52), .B(n988), .Z(n989) );
  NAND2_X1 U1084 ( .A1(G29), .A2(n989), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1023) );
  XNOR2_X1 U1087 ( .A(G16), .B(KEYINPUT125), .ZN(n994) );
  XNOR2_X1 U1088 ( .A(n994), .B(KEYINPUT56), .ZN(n1020) );
  XNOR2_X1 U1089 ( .A(n995), .B(G1341), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n996), .B(G1348), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(G1966), .B(G168), .Z(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(KEYINPUT57), .B(n999), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1018) );
  NAND2_X1 U1096 ( .A1(G1971), .A2(G303), .ZN(n1004) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(G1956), .B(n1012), .Z(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(KEYINPUT126), .B(n1021), .Z(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

