

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801;

  AND2_X1 U372 ( .A1(n465), .A2(n470), .ZN(n728) );
  AND2_X1 U373 ( .A1(n417), .A2(n466), .ZN(n729) );
  BUF_X1 U374 ( .A(n788), .Z(n792) );
  AND2_X1 U375 ( .A1(n649), .A2(n428), .ZN(n427) );
  AND2_X1 U376 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U377 ( .A(n577), .B(KEYINPUT42), .ZN(n680) );
  BUF_X1 U378 ( .A(n615), .Z(n351) );
  XNOR2_X1 U379 ( .A(n350), .B(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U380 ( .A1(n371), .A2(n448), .ZN(n350) );
  XNOR2_X1 U381 ( .A(n356), .B(n583), .ZN(n615) );
  OR2_X1 U382 ( .A1(n645), .A2(n572), .ZN(n579) );
  XNOR2_X1 U383 ( .A(n357), .B(G469), .ZN(n356) );
  NOR2_X1 U384 ( .A1(n667), .A2(G902), .ZN(n421) );
  XNOR2_X1 U385 ( .A(n403), .B(G119), .ZN(n513) );
  XNOR2_X1 U386 ( .A(n512), .B(G104), .ZN(n542) );
  XNOR2_X1 U387 ( .A(G146), .B(G125), .ZN(n521) );
  XNOR2_X1 U388 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n390) );
  XNOR2_X1 U389 ( .A(G119), .B(G128), .ZN(n391) );
  XNOR2_X2 U390 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X2 U391 ( .A1(n382), .A2(n379), .ZN(n623) );
  OR2_X2 U392 ( .A1(n722), .A2(n525), .ZN(n530) );
  NOR2_X2 U393 ( .A1(n767), .A2(n766), .ZN(n769) );
  XNOR2_X1 U394 ( .A(G137), .B(G113), .ZN(n442) );
  NOR2_X2 U395 ( .A1(G953), .A2(G237), .ZN(n541) );
  AND2_X2 U396 ( .A1(n378), .A2(n525), .ZN(n449) );
  AND2_X2 U397 ( .A1(n398), .A2(n358), .ZN(n396) );
  AND2_X2 U398 ( .A1(n438), .A2(n434), .ZN(n433) );
  XNOR2_X2 U399 ( .A(n368), .B(n662), .ZN(n685) );
  NAND2_X2 U400 ( .A1(n433), .A2(n431), .ZN(n664) );
  NAND2_X1 U401 ( .A1(n774), .A2(n782), .ZN(n639) );
  INV_X1 U402 ( .A(n734), .ZN(n732) );
  NOR2_X1 U403 ( .A1(G902), .A2(n707), .ZN(n548) );
  INV_X2 U404 ( .A(G953), .ZN(n793) );
  NAND2_X1 U405 ( .A1(n593), .A2(n598), .ZN(n566) );
  XNOR2_X1 U406 ( .A(n542), .B(n513), .ZN(n410) );
  NAND2_X1 U407 ( .A1(n432), .A2(n436), .ZN(n431) );
  NAND2_X1 U408 ( .A1(n627), .A2(n626), .ZN(n628) );
  AND2_X1 U409 ( .A1(n384), .A2(n364), .ZN(n382) );
  XNOR2_X1 U410 ( .A(n387), .B(n386), .ZN(n550) );
  XNOR2_X1 U411 ( .A(G110), .B(KEYINPUT92), .ZN(n473) );
  XNOR2_X1 U412 ( .A(n416), .B(n469), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n416), .B(n469), .ZN(n666) );
  XNOR2_X1 U414 ( .A(n419), .B(KEYINPUT94), .ZN(n629) );
  NOR2_X2 U415 ( .A1(n666), .A2(n729), .ZN(n353) );
  NOR2_X1 U416 ( .A1(n352), .A2(n729), .ZN(n354) );
  BUF_X1 U417 ( .A(n763), .Z(n355) );
  NOR2_X1 U418 ( .A1(n352), .A2(n729), .ZN(n719) );
  XNOR2_X1 U419 ( .A(n357), .B(G469), .ZN(n584) );
  NOR2_X2 U420 ( .A1(n712), .A2(G902), .ZN(n357) );
  XNOR2_X2 U421 ( .A(n399), .B(KEYINPUT40), .ZN(n683) );
  NAND2_X2 U422 ( .A1(n396), .A2(n394), .ZN(n399) );
  XNOR2_X2 U423 ( .A(n628), .B(KEYINPUT35), .ZN(n682) );
  INV_X1 U424 ( .A(G902), .ZN(n508) );
  INV_X1 U425 ( .A(KEYINPUT95), .ZN(n445) );
  XNOR2_X1 U426 ( .A(n446), .B(n442), .ZN(n441) );
  XNOR2_X1 U427 ( .A(G116), .B(KEYINPUT5), .ZN(n446) );
  AND2_X1 U428 ( .A1(n435), .A2(n681), .ZN(n434) );
  NAND2_X1 U429 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X1 U430 ( .A(KEYINPUT4), .B(G131), .ZN(n489) );
  AND2_X1 U431 ( .A1(n503), .A2(n455), .ZN(n454) );
  NAND2_X1 U432 ( .A1(n731), .A2(KEYINPUT30), .ZN(n455) );
  INV_X1 U433 ( .A(n579), .ZN(n407) );
  XNOR2_X1 U434 ( .A(G116), .B(G107), .ZN(n557) );
  INV_X1 U435 ( .A(KEYINPUT65), .ZN(n469) );
  OR2_X1 U436 ( .A1(n642), .A2(n641), .ZN(n644) );
  XNOR2_X1 U437 ( .A(n630), .B(KEYINPUT6), .ZN(n651) );
  NAND2_X1 U438 ( .A1(n550), .A2(G221), .ZN(n385) );
  NOR2_X1 U439 ( .A1(n793), .A2(G952), .ZN(n725) );
  INV_X1 U440 ( .A(n786), .ZN(n437) );
  AND2_X1 U441 ( .A1(n786), .A2(KEYINPUT81), .ZN(n439) );
  INV_X1 U442 ( .A(KEYINPUT81), .ZN(n436) );
  NAND2_X1 U443 ( .A1(n430), .A2(n658), .ZN(n428) );
  INV_X1 U444 ( .A(G237), .ZN(n507) );
  XOR2_X1 U445 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n483) );
  XOR2_X1 U446 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n534) );
  XNOR2_X1 U447 ( .A(G131), .B(KEYINPUT97), .ZN(n533) );
  XNOR2_X1 U448 ( .A(G143), .B(G140), .ZN(n536) );
  XNOR2_X1 U449 ( .A(G104), .B(G101), .ZN(n495) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n499) );
  NAND2_X1 U451 ( .A1(n377), .A2(KEYINPUT109), .ZN(n376) );
  NAND2_X1 U452 ( .A1(n745), .A2(n616), .ZN(n373) );
  XNOR2_X1 U453 ( .A(n548), .B(n547), .ZN(n597) );
  XNOR2_X1 U454 ( .A(n546), .B(G475), .ZN(n547) );
  XNOR2_X1 U455 ( .A(n443), .B(n441), .ZN(n504) );
  XNOR2_X1 U456 ( .A(n444), .B(n445), .ZN(n443) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n393), .B(n473), .ZN(n392) );
  NAND2_X1 U459 ( .A1(n477), .A2(n476), .ZN(n393) );
  INV_X1 U460 ( .A(KEYINPUT8), .ZN(n386) );
  NAND2_X1 U461 ( .A1(n793), .A2(G234), .ZN(n387) );
  XNOR2_X1 U462 ( .A(G122), .B(KEYINPUT7), .ZN(n556) );
  XOR2_X1 U463 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n555) );
  XNOR2_X1 U464 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n518) );
  XNOR2_X1 U465 ( .A(KEYINPUT86), .B(KEYINPUT4), .ZN(n520) );
  INV_X1 U466 ( .A(KEYINPUT80), .ZN(n418) );
  INV_X1 U467 ( .A(n625), .ZN(n626) );
  NAND2_X1 U468 ( .A1(n381), .A2(n380), .ZN(n379) );
  INV_X1 U469 ( .A(KEYINPUT108), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n353), .A2(G472), .ZN(n668) );
  XNOR2_X1 U471 ( .A(n410), .B(n515), .ZN(n693) );
  NAND2_X1 U472 ( .A1(n395), .A2(n532), .ZN(n394) );
  AND2_X1 U473 ( .A1(n653), .A2(n413), .ZN(n654) );
  AND2_X1 U474 ( .A1(n652), .A2(n414), .ZN(n413) );
  INV_X1 U475 ( .A(n779), .ZN(n567) );
  NAND2_X1 U476 ( .A1(n354), .A2(G217), .ZN(n699) );
  INV_X1 U477 ( .A(n651), .ZN(n448) );
  INV_X1 U478 ( .A(n731), .ZN(n402) );
  AND2_X1 U479 ( .A1(n567), .A2(n397), .ZN(n358) );
  NOR2_X1 U480 ( .A1(n800), .A2(n778), .ZN(n359) );
  AND2_X1 U481 ( .A1(n402), .A2(n458), .ZN(n360) );
  XNOR2_X1 U482 ( .A(n415), .B(n447), .ZN(n361) );
  OR2_X1 U483 ( .A1(n595), .A2(KEYINPUT47), .ZN(n362) );
  INV_X1 U484 ( .A(KEYINPUT30), .ZN(n458) );
  INV_X1 U485 ( .A(n655), .ZN(n414) );
  AND2_X1 U486 ( .A1(n734), .A2(n447), .ZN(n363) );
  OR2_X1 U487 ( .A1(n402), .A2(n383), .ZN(n364) );
  XOR2_X1 U488 ( .A(n667), .B(KEYINPUT62), .Z(n365) );
  XNOR2_X1 U489 ( .A(KEYINPUT15), .B(G902), .ZN(n663) );
  INV_X1 U490 ( .A(KEYINPUT84), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n606), .B(KEYINPUT48), .ZN(n366) );
  NAND2_X1 U492 ( .A1(KEYINPUT84), .A2(KEYINPUT44), .ZN(n367) );
  NAND2_X1 U493 ( .A1(n685), .A2(n470), .ZN(n378) );
  NAND2_X1 U494 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U495 ( .A1(n660), .A2(n659), .ZN(n369) );
  XNOR2_X1 U496 ( .A(n650), .B(KEYINPUT83), .ZN(n370) );
  NAND2_X1 U497 ( .A1(n615), .A2(n616), .ZN(n374) );
  OR2_X1 U498 ( .A1(n615), .A2(n745), .ZN(n635) );
  NOR2_X1 U499 ( .A1(n375), .A2(n372), .ZN(n371) );
  NAND2_X1 U500 ( .A1(n374), .A2(n373), .ZN(n372) );
  NOR2_X1 U501 ( .A1(n376), .A2(n615), .ZN(n375) );
  INV_X1 U502 ( .A(n745), .ZN(n377) );
  NOR2_X1 U503 ( .A1(n731), .A2(n589), .ZN(n380) );
  INV_X1 U504 ( .A(n610), .ZN(n381) );
  INV_X1 U505 ( .A(n589), .ZN(n383) );
  NAND2_X1 U506 ( .A1(n610), .A2(n589), .ZN(n384) );
  NAND2_X1 U507 ( .A1(n623), .A2(n622), .ZN(n401) );
  XNOR2_X1 U508 ( .A(n388), .B(n385), .ZN(n480) );
  XNOR2_X1 U509 ( .A(n392), .B(n389), .ZN(n388) );
  NAND2_X1 U510 ( .A1(n602), .A2(n734), .ZN(n415) );
  INV_X1 U511 ( .A(n596), .ZN(n395) );
  OR2_X1 U512 ( .A1(n734), .A2(n447), .ZN(n397) );
  NAND2_X1 U513 ( .A1(n596), .A2(n363), .ZN(n398) );
  XNOR2_X1 U514 ( .A(n665), .B(n418), .ZN(n417) );
  BUF_X1 U515 ( .A(n682), .Z(n420) );
  AND2_X1 U516 ( .A1(n433), .A2(n431), .ZN(n400) );
  BUF_X1 U517 ( .A(n645), .Z(n655) );
  NOR2_X1 U518 ( .A1(n605), .A2(n461), .ZN(n460) );
  XNOR2_X2 U519 ( .A(n401), .B(KEYINPUT0), .ZN(n642) );
  XNOR2_X2 U520 ( .A(G101), .B(KEYINPUT3), .ZN(n403) );
  NAND2_X1 U521 ( .A1(n404), .A2(n426), .ZN(n429) );
  NAND2_X1 U522 ( .A1(n405), .A2(KEYINPUT84), .ZN(n404) );
  INV_X1 U523 ( .A(n682), .ZN(n405) );
  INV_X1 U524 ( .A(n408), .ZN(n409) );
  NAND2_X1 U525 ( .A1(n408), .A2(n360), .ZN(n452) );
  XNOR2_X2 U526 ( .A(n578), .B(n406), .ZN(n408) );
  AND2_X1 U527 ( .A1(n414), .A2(n409), .ZN(n656) );
  NAND2_X1 U528 ( .A1(n408), .A2(n407), .ZN(n574) );
  NOR2_X1 U529 ( .A1(n408), .A2(n458), .ZN(n450) );
  NAND2_X1 U530 ( .A1(n411), .A2(n658), .ZN(n660) );
  NAND2_X1 U531 ( .A1(n412), .A2(n359), .ZN(n411) );
  INV_X1 U532 ( .A(n420), .ZN(n412) );
  XNOR2_X2 U533 ( .A(n457), .B(n511), .ZN(n596) );
  XNOR2_X2 U534 ( .A(n664), .B(KEYINPUT78), .ZN(n788) );
  NAND2_X1 U535 ( .A1(n468), .A2(n449), .ZN(n416) );
  NOR2_X2 U536 ( .A1(n584), .A2(n614), .ZN(n419) );
  XNOR2_X2 U537 ( .A(n634), .B(KEYINPUT96), .ZN(n774) );
  NAND2_X1 U538 ( .A1(n683), .A2(n680), .ZN(n464) );
  XNOR2_X2 U539 ( .A(n421), .B(G472), .ZN(n578) );
  NOR2_X1 U540 ( .A1(n451), .A2(n450), .ZN(n453) );
  NAND2_X1 U541 ( .A1(n422), .A2(n763), .ZN(n424) );
  INV_X1 U542 ( .A(n633), .ZN(n422) );
  XNOR2_X1 U543 ( .A(n642), .B(KEYINPUT90), .ZN(n633) );
  BUF_X2 U544 ( .A(n610), .Z(n423) );
  XNOR2_X1 U545 ( .A(n424), .B(n472), .ZN(n627) );
  NAND2_X1 U546 ( .A1(n682), .A2(n367), .ZN(n426) );
  NAND2_X1 U547 ( .A1(n429), .A2(n427), .ZN(n650) );
  INV_X1 U548 ( .A(n440), .ZN(n432) );
  NAND2_X1 U549 ( .A1(n440), .A2(n439), .ZN(n438) );
  XNOR2_X1 U550 ( .A(n459), .B(n366), .ZN(n440) );
  NAND2_X1 U551 ( .A1(n541), .A2(G210), .ZN(n444) );
  INV_X1 U552 ( .A(n532), .ZN(n447) );
  NAND2_X1 U553 ( .A1(n362), .A2(n784), .ZN(n461) );
  NAND2_X1 U554 ( .A1(n467), .A2(n466), .ZN(n465) );
  NAND2_X1 U555 ( .A1(n452), .A2(n454), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n456), .A2(n453), .ZN(n457) );
  XNOR2_X1 U557 ( .A(n629), .B(KEYINPUT112), .ZN(n456) );
  NAND2_X1 U558 ( .A1(n462), .A2(n460), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n464), .B(n463), .ZN(n462) );
  INV_X1 U560 ( .A(KEYINPUT46), .ZN(n463) );
  INV_X1 U561 ( .A(n685), .ZN(n466) );
  INV_X1 U562 ( .A(n792), .ZN(n467) );
  NAND2_X1 U563 ( .A1(n788), .A2(n470), .ZN(n468) );
  INV_X1 U564 ( .A(KEYINPUT2), .ZN(n470) );
  XNOR2_X2 U565 ( .A(n485), .B(n484), .ZN(n570) );
  AND2_X1 U566 ( .A1(n581), .A2(n567), .ZN(n471) );
  XOR2_X1 U567 ( .A(n624), .B(KEYINPUT69), .Z(n472) );
  XNOR2_X1 U568 ( .A(n536), .B(n535), .ZN(n537) );
  BUF_X1 U569 ( .A(n712), .Z(n715) );
  INV_X1 U570 ( .A(n725), .ZN(n669) );
  BUF_X1 U571 ( .A(n698), .Z(n700) );
  BUF_X1 U572 ( .A(n683), .Z(n684) );
  INV_X1 U573 ( .A(KEYINPUT91), .ZN(n474) );
  NAND2_X1 U574 ( .A1(KEYINPUT77), .A2(n474), .ZN(n477) );
  INV_X1 U575 ( .A(KEYINPUT77), .ZN(n475) );
  NAND2_X1 U576 ( .A1(n475), .A2(KEYINPUT91), .ZN(n476) );
  XNOR2_X1 U577 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n521), .B(n478), .ZN(n539) );
  INV_X1 U579 ( .A(G137), .ZN(n479) );
  XNOR2_X1 U580 ( .A(n479), .B(G140), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n539), .B(n491), .ZN(n791) );
  XNOR2_X1 U582 ( .A(n480), .B(n791), .ZN(n698) );
  NAND2_X1 U583 ( .A1(n698), .A2(n508), .ZN(n485) );
  NAND2_X1 U584 ( .A1(G234), .A2(n663), .ZN(n481) );
  XNOR2_X1 U585 ( .A(KEYINPUT20), .B(n481), .ZN(n486) );
  NAND2_X1 U586 ( .A1(n486), .A2(G217), .ZN(n482) );
  XOR2_X1 U587 ( .A(n483), .B(n482), .Z(n484) );
  NAND2_X1 U588 ( .A1(n486), .A2(G221), .ZN(n487) );
  XNOR2_X1 U589 ( .A(n487), .B(KEYINPUT21), .ZN(n741) );
  INV_X1 U590 ( .A(n741), .ZN(n640) );
  NAND2_X1 U591 ( .A1(n570), .A2(n640), .ZN(n614) );
  XNOR2_X2 U592 ( .A(G143), .B(G128), .ZN(n516) );
  INV_X1 U593 ( .A(G134), .ZN(n488) );
  XNOR2_X2 U594 ( .A(n516), .B(n488), .ZN(n551) );
  XNOR2_X2 U595 ( .A(n551), .B(n489), .ZN(n789) );
  XNOR2_X2 U596 ( .A(n789), .B(G146), .ZN(n505) );
  NAND2_X1 U597 ( .A1(n793), .A2(G227), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n490), .B(KEYINPUT72), .ZN(n493) );
  INV_X1 U599 ( .A(n491), .ZN(n492) );
  XNOR2_X1 U600 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U601 ( .A(G107), .B(G110), .ZN(n494) );
  XNOR2_X1 U602 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U603 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U604 ( .A(n505), .B(n498), .ZN(n712) );
  XNOR2_X1 U605 ( .A(n499), .B(KEYINPUT14), .ZN(n500) );
  NAND2_X1 U606 ( .A1(G952), .A2(n500), .ZN(n759) );
  NOR2_X1 U607 ( .A1(n759), .A2(G953), .ZN(n619) );
  NAND2_X1 U608 ( .A1(G902), .A2(n500), .ZN(n617) );
  OR2_X1 U609 ( .A1(n793), .A2(n617), .ZN(n501) );
  NOR2_X1 U610 ( .A1(n501), .A2(G900), .ZN(n502) );
  NOR2_X1 U611 ( .A1(n619), .A2(n502), .ZN(n571) );
  INV_X1 U612 ( .A(n571), .ZN(n503) );
  XOR2_X1 U613 ( .A(n504), .B(n513), .Z(n506) );
  XNOR2_X1 U614 ( .A(n505), .B(n506), .ZN(n667) );
  NAND2_X1 U615 ( .A1(n508), .A2(n507), .ZN(n526) );
  NAND2_X1 U616 ( .A1(n526), .A2(G214), .ZN(n510) );
  INV_X1 U617 ( .A(KEYINPUT88), .ZN(n509) );
  XNOR2_X1 U618 ( .A(n510), .B(n509), .ZN(n731) );
  INV_X1 U619 ( .A(KEYINPUT70), .ZN(n511) );
  XNOR2_X2 U620 ( .A(G122), .B(G113), .ZN(n512) );
  XNOR2_X1 U621 ( .A(KEYINPUT16), .B(G110), .ZN(n514) );
  XNOR2_X1 U622 ( .A(n557), .B(n514), .ZN(n515) );
  NAND2_X1 U623 ( .A1(n793), .A2(G224), .ZN(n517) );
  XNOR2_X1 U624 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U625 ( .A(n516), .B(n519), .ZN(n523) );
  XNOR2_X1 U626 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U627 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U628 ( .A(n693), .B(n524), .ZN(n722) );
  INV_X1 U629 ( .A(n663), .ZN(n525) );
  NAND2_X1 U630 ( .A1(n526), .A2(G210), .ZN(n528) );
  INV_X1 U631 ( .A(KEYINPUT87), .ZN(n527) );
  XNOR2_X1 U632 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X2 U633 ( .A(n530), .B(n529), .ZN(n610) );
  XNOR2_X2 U634 ( .A(n423), .B(KEYINPUT38), .ZN(n734) );
  INV_X1 U635 ( .A(KEYINPUT68), .ZN(n531) );
  XNOR2_X1 U636 ( .A(n531), .B(KEYINPUT39), .ZN(n532) );
  XNOR2_X1 U637 ( .A(n534), .B(n533), .ZN(n538) );
  INV_X1 U638 ( .A(KEYINPUT98), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n538), .B(n537), .ZN(n540) );
  XNOR2_X1 U640 ( .A(n540), .B(n539), .ZN(n545) );
  NAND2_X1 U641 ( .A1(G214), .A2(n541), .ZN(n543) );
  XOR2_X1 U642 ( .A(n543), .B(n542), .Z(n544) );
  XNOR2_X1 U643 ( .A(n545), .B(n544), .ZN(n707) );
  XNOR2_X1 U644 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n546) );
  INV_X1 U645 ( .A(KEYINPUT100), .ZN(n549) );
  XNOR2_X1 U646 ( .A(n597), .B(n549), .ZN(n593) );
  XNOR2_X1 U647 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n563) );
  NAND2_X1 U648 ( .A1(n550), .A2(G217), .ZN(n553) );
  BUF_X1 U649 ( .A(n551), .Z(n552) );
  XNOR2_X1 U650 ( .A(n553), .B(n552), .ZN(n561) );
  XNOR2_X1 U651 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n554) );
  XNOR2_X1 U652 ( .A(n555), .B(n554), .ZN(n559) );
  XNOR2_X1 U653 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U654 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U655 ( .A(n561), .B(n560), .ZN(n702) );
  NOR2_X1 U656 ( .A1(G902), .A2(n702), .ZN(n562) );
  XNOR2_X1 U657 ( .A(n563), .B(n562), .ZN(n565) );
  INV_X1 U658 ( .A(G478), .ZN(n564) );
  XNOR2_X1 U659 ( .A(n565), .B(n564), .ZN(n598) );
  XNOR2_X2 U660 ( .A(n566), .B(KEYINPUT106), .ZN(n779) );
  AND2_X1 U661 ( .A1(n597), .A2(n598), .ZN(n736) );
  NAND2_X1 U662 ( .A1(n736), .A2(n402), .ZN(n568) );
  NOR2_X1 U663 ( .A1(n568), .A2(n732), .ZN(n569) );
  XNOR2_X1 U664 ( .A(n569), .B(KEYINPUT41), .ZN(n753) );
  BUF_X1 U665 ( .A(n570), .Z(n645) );
  OR2_X1 U666 ( .A1(n741), .A2(n571), .ZN(n572) );
  INV_X1 U667 ( .A(KEYINPUT28), .ZN(n573) );
  XNOR2_X1 U668 ( .A(n574), .B(n573), .ZN(n576) );
  INV_X1 U669 ( .A(n356), .ZN(n575) );
  NAND2_X1 U670 ( .A1(n576), .A2(n575), .ZN(n587) );
  OR2_X1 U671 ( .A1(n753), .A2(n587), .ZN(n577) );
  INV_X1 U672 ( .A(n578), .ZN(n630) );
  NOR2_X1 U673 ( .A1(n651), .A2(n579), .ZN(n580) );
  XNOR2_X1 U674 ( .A(n580), .B(KEYINPUT110), .ZN(n581) );
  NAND2_X1 U675 ( .A1(n471), .A2(n402), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n607), .A2(n423), .ZN(n582) );
  XNOR2_X1 U677 ( .A(n582), .B(KEYINPUT36), .ZN(n586) );
  XNOR2_X1 U678 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n583) );
  INV_X1 U679 ( .A(n351), .ZN(n585) );
  NAND2_X1 U680 ( .A1(n586), .A2(n585), .ZN(n784) );
  INV_X1 U681 ( .A(n587), .ZN(n590) );
  INV_X1 U682 ( .A(KEYINPUT71), .ZN(n588) );
  XNOR2_X1 U683 ( .A(n588), .B(KEYINPUT19), .ZN(n589) );
  NAND2_X1 U684 ( .A1(n590), .A2(n623), .ZN(n592) );
  INV_X1 U685 ( .A(KEYINPUT74), .ZN(n591) );
  XNOR2_X2 U686 ( .A(n592), .B(n591), .ZN(n675) );
  OR2_X1 U687 ( .A1(n593), .A2(n598), .ZN(n674) );
  INV_X1 U688 ( .A(KEYINPUT107), .ZN(n594) );
  XNOR2_X1 U689 ( .A(n674), .B(n594), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n779), .A2(n612), .ZN(n638) );
  NAND2_X1 U691 ( .A1(n675), .A2(n638), .ZN(n595) );
  NAND2_X1 U692 ( .A1(n595), .A2(KEYINPUT47), .ZN(n603) );
  BUF_X1 U693 ( .A(n596), .Z(n602) );
  INV_X1 U694 ( .A(n597), .ZN(n600) );
  INV_X1 U695 ( .A(n598), .ZN(n599) );
  NAND2_X1 U696 ( .A1(n600), .A2(n599), .ZN(n625) );
  NOR2_X1 U697 ( .A1(n625), .A2(n423), .ZN(n601) );
  NAND2_X1 U698 ( .A1(n602), .A2(n601), .ZN(n679) );
  NAND2_X1 U699 ( .A1(n603), .A2(n679), .ZN(n604) );
  XNOR2_X1 U700 ( .A(n604), .B(KEYINPUT76), .ZN(n605) );
  INV_X1 U701 ( .A(KEYINPUT82), .ZN(n606) );
  XNOR2_X1 U702 ( .A(n607), .B(KEYINPUT111), .ZN(n608) );
  NAND2_X1 U703 ( .A1(n608), .A2(n351), .ZN(n609) );
  XNOR2_X1 U704 ( .A(n609), .B(KEYINPUT43), .ZN(n611) );
  NAND2_X1 U705 ( .A1(n611), .A2(n423), .ZN(n786) );
  INV_X1 U706 ( .A(n612), .ZN(n613) );
  NAND2_X1 U707 ( .A1(n361), .A2(n613), .ZN(n681) );
  BUF_X1 U708 ( .A(n614), .Z(n745) );
  INV_X1 U709 ( .A(KEYINPUT109), .ZN(n616) );
  INV_X1 U710 ( .A(G898), .ZN(n689) );
  NAND2_X1 U711 ( .A1(G953), .A2(n689), .ZN(n694) );
  NOR2_X1 U712 ( .A1(n694), .A2(n617), .ZN(n618) );
  OR2_X1 U713 ( .A1(n619), .A2(n618), .ZN(n621) );
  INV_X1 U714 ( .A(KEYINPUT89), .ZN(n620) );
  XNOR2_X1 U715 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U716 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n624) );
  BUF_X1 U717 ( .A(n629), .Z(n631) );
  INV_X1 U718 ( .A(n630), .ZN(n743) );
  NAND2_X1 U719 ( .A1(n631), .A2(n743), .ZN(n632) );
  OR2_X1 U720 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U721 ( .A1(n635), .A2(n743), .ZN(n750) );
  OR2_X1 U722 ( .A1(n750), .A2(n642), .ZN(n637) );
  INV_X1 U723 ( .A(KEYINPUT31), .ZN(n636) );
  XNOR2_X1 U724 ( .A(n637), .B(n636), .ZN(n782) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n736), .A2(n640), .ZN(n641) );
  INV_X1 U727 ( .A(KEYINPUT22), .ZN(n643) );
  XNOR2_X1 U728 ( .A(n644), .B(n643), .ZN(n653) );
  AND2_X1 U729 ( .A1(n653), .A2(n351), .ZN(n657) );
  AND2_X1 U730 ( .A1(n651), .A2(n655), .ZN(n646) );
  AND2_X1 U731 ( .A1(n657), .A2(n646), .ZN(n770) );
  INV_X1 U732 ( .A(n770), .ZN(n647) );
  NOR2_X1 U733 ( .A1(n448), .A2(n351), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n654), .B(KEYINPUT32), .ZN(n800) );
  AND2_X1 U735 ( .A1(n657), .A2(n656), .ZN(n778) );
  INV_X1 U736 ( .A(KEYINPUT44), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n359), .A2(KEYINPUT44), .ZN(n659) );
  XNOR2_X1 U738 ( .A(KEYINPUT79), .B(KEYINPUT45), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT64), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n400), .A2(KEYINPUT2), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n668), .B(n365), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n671), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U744 ( .A1(n675), .A2(n567), .ZN(n673) );
  XOR2_X1 U745 ( .A(G146), .B(KEYINPUT115), .Z(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G48) );
  INV_X1 U747 ( .A(n674), .ZN(n773) );
  NAND2_X1 U748 ( .A1(n675), .A2(n773), .ZN(n677) );
  XOR2_X1 U749 ( .A(G128), .B(KEYINPUT29), .Z(n676) );
  XNOR2_X1 U750 ( .A(n677), .B(n676), .ZN(G30) );
  XNOR2_X1 U751 ( .A(G143), .B(KEYINPUT114), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n679), .B(n678), .ZN(G45) );
  XNOR2_X1 U753 ( .A(n680), .B(G137), .ZN(G39) );
  XNOR2_X1 U754 ( .A(n681), .B(G134), .ZN(G36) );
  XOR2_X1 U755 ( .A(G122), .B(n420), .Z(G24) );
  XNOR2_X1 U756 ( .A(n684), .B(G131), .ZN(G33) );
  NOR2_X1 U757 ( .A1(n685), .A2(G953), .ZN(n692) );
  NAND2_X1 U758 ( .A1(G224), .A2(G953), .ZN(n686) );
  XNOR2_X1 U759 ( .A(n686), .B(KEYINPUT61), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(KEYINPUT125), .ZN(n688) );
  NOR2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U762 ( .A(n690), .B(KEYINPUT126), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U764 ( .A(n693), .ZN(n695) );
  NAND2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n697), .B(n696), .ZN(G69) );
  XOR2_X1 U767 ( .A(n700), .B(n699), .Z(n701) );
  NOR2_X1 U768 ( .A1(n701), .A2(n725), .ZN(G66) );
  NAND2_X1 U769 ( .A1(n354), .A2(G478), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT124), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n705), .A2(n725), .ZN(G63) );
  NAND2_X1 U773 ( .A1(n353), .A2(G475), .ZN(n709) );
  XNOR2_X1 U774 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U776 ( .A1(n710), .A2(n725), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U778 ( .A1(n354), .A2(G469), .ZN(n717) );
  XOR2_X1 U779 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n713) );
  XNOR2_X1 U780 ( .A(n713), .B(KEYINPUT58), .ZN(n714) );
  XNOR2_X1 U781 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n718), .A2(n725), .ZN(G54) );
  NAND2_X1 U784 ( .A1(n719), .A2(G210), .ZN(n724) );
  XNOR2_X1 U785 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n720) );
  XNOR2_X1 U786 ( .A(n720), .B(KEYINPUT55), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U788 ( .A(n724), .B(n723), .ZN(n726) );
  NOR2_X1 U789 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U790 ( .A(n727), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U791 ( .A(KEYINPUT75), .B(n728), .Z(n730) );
  NOR2_X1 U792 ( .A1(n730), .A2(n729), .ZN(n767) );
  NOR2_X1 U793 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U794 ( .A1(n638), .A2(n733), .ZN(n739) );
  NOR2_X1 U795 ( .A1(n734), .A2(n402), .ZN(n735) );
  XNOR2_X1 U796 ( .A(n735), .B(KEYINPUT119), .ZN(n737) );
  NAND2_X1 U797 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U798 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U799 ( .A1(n740), .A2(n355), .ZN(n756) );
  NAND2_X1 U800 ( .A1(n414), .A2(n741), .ZN(n742) );
  XOR2_X1 U801 ( .A(KEYINPUT49), .B(n742), .Z(n744) );
  NAND2_X1 U802 ( .A1(n744), .A2(n743), .ZN(n749) );
  NAND2_X1 U803 ( .A1(n351), .A2(n745), .ZN(n747) );
  XOR2_X1 U804 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n746) );
  XNOR2_X1 U805 ( .A(n747), .B(n746), .ZN(n748) );
  OR2_X1 U806 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U808 ( .A(KEYINPUT51), .B(n752), .Z(n754) );
  INV_X1 U809 ( .A(n753), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n754), .A2(n762), .ZN(n755) );
  AND2_X1 U811 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U812 ( .A(n757), .B(KEYINPUT52), .ZN(n758) );
  XNOR2_X1 U813 ( .A(KEYINPUT120), .B(n758), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U815 ( .A1(n761), .A2(G953), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n355), .A2(n762), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U818 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n768) );
  XNOR2_X1 U819 ( .A(n769), .B(n768), .ZN(G75) );
  XNOR2_X1 U820 ( .A(G101), .B(n770), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n771), .B(KEYINPUT113), .ZN(G3) );
  NOR2_X1 U822 ( .A1(n779), .A2(n774), .ZN(n772) );
  XOR2_X1 U823 ( .A(G104), .B(n772), .Z(G6) );
  NOR2_X1 U824 ( .A1(n774), .A2(n674), .ZN(n776) );
  XNOR2_X1 U825 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n775) );
  XNOR2_X1 U826 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U827 ( .A(G107), .B(n777), .ZN(G9) );
  XOR2_X1 U828 ( .A(G110), .B(n778), .Z(G12) );
  NOR2_X1 U829 ( .A1(n779), .A2(n782), .ZN(n780) );
  XOR2_X1 U830 ( .A(KEYINPUT116), .B(n780), .Z(n781) );
  XNOR2_X1 U831 ( .A(G113), .B(n781), .ZN(G15) );
  NOR2_X1 U832 ( .A1(n674), .A2(n782), .ZN(n783) );
  XOR2_X1 U833 ( .A(G116), .B(n783), .Z(G18) );
  XOR2_X1 U834 ( .A(n784), .B(G125), .Z(n785) );
  XNOR2_X1 U835 ( .A(n785), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U836 ( .A(G140), .B(n786), .Z(n787) );
  XNOR2_X1 U837 ( .A(n787), .B(KEYINPUT117), .ZN(G42) );
  BUF_X1 U838 ( .A(n789), .Z(n790) );
  XNOR2_X1 U839 ( .A(n790), .B(n791), .ZN(n795) );
  XNOR2_X1 U840 ( .A(n792), .B(n795), .ZN(n794) );
  NAND2_X1 U841 ( .A1(n794), .A2(n793), .ZN(n799) );
  XNOR2_X1 U842 ( .A(n795), .B(G227), .ZN(n796) );
  NAND2_X1 U843 ( .A1(n796), .A2(G900), .ZN(n797) );
  NAND2_X1 U844 ( .A1(n797), .A2(G953), .ZN(n798) );
  NAND2_X1 U845 ( .A1(n799), .A2(n798), .ZN(G72) );
  XNOR2_X1 U846 ( .A(G119), .B(KEYINPUT127), .ZN(n801) );
  XNOR2_X1 U847 ( .A(n801), .B(n800), .ZN(G21) );
endmodule

