//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XNOR2_X1  g0004(.A(KEYINPUT65), .B(G20), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n202), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT66), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n210), .B(new_n215), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  OAI211_X1 g0048(.A(G1), .B(G13), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G274), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n206), .B1(G33), .B2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(new_n252), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(G226), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n258), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(G1698), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT69), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(G223), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n249), .B(KEYINPUT70), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n257), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G200), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n206), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  INV_X1    g0072(.A(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n247), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n205), .A2(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n280), .A2(new_n273), .A3(G1), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n270), .ZN(new_n282));
  INV_X1    g0082(.A(G50), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n251), .B2(G20), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n282), .A2(new_n284), .B1(new_n283), .B2(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT9), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n268), .B(new_n287), .C1(new_n288), .C2(new_n267), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT10), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT71), .B(G179), .Z(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n267), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n267), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n286), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n276), .A2(new_n261), .B1(new_n273), .B2(G68), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT74), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n283), .B2(new_n274), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  OAI211_X1 g0101(.A(KEYINPUT11), .B(new_n270), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n280), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G20), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n306));
  INV_X1    g0106(.A(G68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n251), .B2(G20), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n305), .A2(new_n306), .B1(new_n282), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n270), .B1(new_n300), .B2(new_n301), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT11), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n253), .B1(G238), .B2(new_n256), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n249), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  INV_X1    g0118(.A(G232), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G226), .B2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n318), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n315), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(G169), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(G179), .A3(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n332), .B2(G169), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n314), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(G200), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n329), .A2(G190), .A3(new_n331), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n339), .A2(new_n310), .A3(new_n313), .A4(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n282), .B(G77), .C1(G1), .C2(new_n273), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n304), .A2(KEYINPUT73), .A3(G77), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT73), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n281), .B2(new_n261), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n277), .ZN(new_n347));
  NOR2_X1   g0147(.A1(G20), .A2(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n273), .A2(KEYINPUT65), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT65), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n347), .A2(new_n348), .B1(new_n352), .B2(G77), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n276), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n346), .B1(new_n270), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n264), .A2(G238), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n259), .A2(G232), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT72), .B1(new_n325), .B2(new_n358), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n325), .A2(KEYINPUT72), .A3(new_n358), .ZN(new_n360));
  INV_X1    g0160(.A(G107), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n258), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n317), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n253), .B1(G244), .B2(new_n256), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n356), .B1(new_n365), .B2(new_n294), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n291), .A3(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n356), .B1(new_n365), .B2(new_n288), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n363), .B2(new_n364), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n297), .A2(new_n338), .A3(new_n341), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT77), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n323), .A2(new_n324), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n322), .A2(KEYINPUT75), .A3(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(G223), .A2(G1698), .ZN(new_n381));
  INV_X1    g0181(.A(G226), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n376), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n378), .B2(new_n379), .ZN(new_n389));
  INV_X1    g0189(.A(new_n387), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n389), .A2(KEYINPUT77), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n317), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n256), .A2(KEYINPUT78), .A3(G232), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n249), .A2(new_n252), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n319), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n253), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n292), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT77), .B1(new_n389), .B2(new_n390), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n322), .A2(KEYINPUT75), .A3(G33), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n258), .B2(new_n377), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n376), .B(new_n387), .C1(new_n401), .C2(new_n384), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n266), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n393), .A2(new_n396), .ZN(new_n404));
  INV_X1    g0204(.A(new_n253), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G159), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT76), .B1(new_n274), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT76), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n348), .A2(new_n411), .A3(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G58), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n307), .ZN(new_n415));
  OAI21_X1  g0215(.A(G20), .B1(new_n415), .B2(new_n201), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n401), .B2(new_n273), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n205), .A2(new_n419), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n380), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n418), .B(KEYINPUT16), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n325), .B2(new_n205), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n273), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n323), .B2(new_n324), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n425), .A2(new_n307), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n424), .B1(new_n428), .B2(new_n417), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n423), .A2(new_n429), .A3(new_n270), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n277), .B1(new_n251), .B2(G20), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n282), .B1(new_n281), .B2(new_n277), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n408), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n408), .A2(new_n436), .A3(new_n433), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n430), .A2(new_n432), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n392), .A2(G190), .A3(new_n397), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n403), .B2(new_n406), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n438), .A2(KEYINPUT17), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n430), .A4(new_n432), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n435), .A2(new_n437), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n375), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n249), .A2(new_n450), .A3(G250), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n249), .A2(G274), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT79), .B1(new_n452), .B2(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n250), .A2(new_n454), .A3(new_n450), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G244), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n457), .B(new_n259), .C1(new_n378), .C2(new_n379), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n380), .A2(G244), .A3(G1698), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT80), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n247), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n259), .A2(G238), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n380), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n447), .B(new_n456), .C1(new_n468), .C2(new_n317), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n458), .B2(KEYINPUT80), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n460), .A2(new_n461), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n317), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n456), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT81), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(G200), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n457), .B1(new_n378), .B2(new_n379), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT80), .B1(new_n476), .B2(G1698), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n401), .A2(new_n465), .B1(new_n247), .B2(new_n463), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n266), .B1(new_n479), .B2(new_n459), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n447), .B1(new_n480), .B2(new_n456), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n472), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(G190), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n354), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n304), .ZN(new_n485));
  INV_X1    g0285(.A(new_n270), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT19), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n205), .B1(new_n487), .B2(new_n318), .ZN(new_n488));
  NOR2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  INV_X1    g0289(.A(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n205), .A2(G33), .A3(G97), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n488), .A2(new_n491), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n380), .A2(G68), .A3(new_n205), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n486), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n251), .A2(G33), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n486), .A2(new_n304), .A3(new_n496), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n485), .B(new_n495), .C1(G87), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n475), .A2(new_n483), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n294), .B1(new_n469), .B2(new_n474), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n481), .A2(new_n291), .A3(new_n482), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n495), .A2(new_n485), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n282), .A2(new_n496), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n354), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT82), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT82), .ZN(new_n507));
  NOR4_X1   g0307(.A1(new_n495), .A2(new_n507), .A3(new_n485), .A4(new_n504), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n501), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n499), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n499), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT83), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n361), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  AND2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n489), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n352), .B1(G77), .B2(new_n348), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT7), .B1(new_n352), .B2(new_n258), .ZN(new_n520));
  INV_X1    g0320(.A(new_n427), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n270), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n304), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G97), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n503), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  NOR2_X1   g0331(.A1(KEYINPUT5), .A2(G41), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(new_n249), .A3(G274), .A4(new_n449), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n254), .B1(new_n533), .B2(new_n449), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G257), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G250), .A2(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(KEYINPUT4), .A2(G244), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(G1698), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n541), .B2(new_n325), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n380), .A2(G244), .A3(new_n259), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n534), .B(new_n536), .C1(new_n545), .C2(new_n266), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n530), .B1(G200), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n546), .A2(new_n288), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n528), .B1(new_n523), .B2(new_n270), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n546), .B2(new_n294), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n545), .A2(new_n266), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(new_n291), .A3(new_n534), .A4(new_n536), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n547), .A2(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT22), .A2(G87), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n401), .A2(new_n352), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n325), .B2(new_n490), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(G20), .B2(new_n361), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n560), .B1(new_n464), .B2(new_n273), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n352), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT23), .B1(new_n273), .B2(G107), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT86), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n557), .A2(new_n561), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT85), .B1(new_n555), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n380), .A2(KEYINPUT22), .A3(G87), .A4(new_n205), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n557), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n567), .B2(new_n571), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n270), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n281), .A2(KEYINPUT25), .A3(new_n361), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT87), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT25), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n304), .B2(G107), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n579), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(G107), .B2(new_n497), .ZN(new_n582));
  INV_X1    g0382(.A(G294), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n247), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G257), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G1698), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G250), .B2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n379), .B2(new_n378), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n317), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n535), .A2(G264), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n534), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n371), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G190), .B2(new_n591), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n575), .A2(new_n582), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n553), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n585), .A2(new_n259), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G264), .B2(new_n259), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n379), .B2(new_n378), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n325), .A2(G303), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT84), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n599), .C1(new_n401), .C2(new_n597), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n317), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n269), .A2(new_n206), .B1(G20), .B2(new_n463), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n537), .B1(new_n527), .B2(G33), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n352), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n304), .A2(G116), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n497), .B2(G116), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n449), .B1(new_n531), .B2(new_n532), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(G270), .A3(new_n249), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n534), .A2(G179), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n605), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n534), .A2(new_n615), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n605), .A2(G190), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n266), .B1(new_n601), .B2(new_n603), .ZN(new_n621));
  OAI21_X1  g0421(.A(G200), .B1(new_n621), .B2(new_n618), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(new_n622), .A3(new_n610), .A4(new_n612), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n605), .A2(new_n619), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n294), .B1(new_n610), .B2(new_n612), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n624), .C1(new_n618), .C2(new_n621), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n617), .B(new_n623), .C1(new_n627), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n591), .A2(new_n294), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(G179), .B2(new_n591), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n575), .B2(new_n582), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n595), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n446), .A2(new_n512), .A3(new_n514), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n296), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n435), .A2(new_n437), .ZN(new_n637));
  INV_X1    g0437(.A(new_n338), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n341), .B2(new_n369), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n441), .A2(new_n444), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(new_n642), .B2(new_n290), .ZN(new_n643));
  INV_X1    g0443(.A(new_n446), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n502), .A2(new_n505), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n472), .A2(new_n473), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n294), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n501), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT88), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT88), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n617), .B1(new_n627), .B2(new_n629), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n594), .B(new_n553), .C1(new_n651), .C2(new_n633), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(G200), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n483), .A2(new_n498), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n649), .B(new_n650), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n550), .A2(new_n552), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n514), .A2(KEYINPUT26), .A3(new_n512), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n655), .B2(new_n657), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n656), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n643), .B1(new_n644), .B2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(new_n633), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n594), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n575), .A2(new_n582), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n205), .A2(new_n303), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n633), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n651), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n613), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n623), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(G330), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n681), .A2(KEYINPUT89), .ZN(new_n682));
  INV_X1    g0482(.A(new_n676), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(G330), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT89), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n677), .A2(new_n672), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n665), .A2(new_n687), .A3(new_n673), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n633), .A2(new_n671), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n213), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n491), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n208), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n514), .A2(new_n634), .A3(new_n512), .A4(new_n671), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT91), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n536), .B1(new_n545), .B2(new_n266), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n616), .A2(new_n589), .A3(new_n590), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n702), .A3(new_n621), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n481), .A2(new_n482), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n481), .A2(new_n703), .A3(KEYINPUT30), .A4(new_n482), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n591), .A2(new_n291), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n619), .B2(new_n605), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT90), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n646), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n472), .A2(KEYINPUT90), .A3(new_n473), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n709), .A2(new_n711), .A3(new_n546), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(new_n707), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(new_n672), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n700), .B1(new_n715), .B2(KEYINPUT31), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n714), .B2(new_n672), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n699), .B(new_n716), .C1(new_n719), .C2(new_n700), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n662), .B2(new_n672), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n655), .A2(new_n660), .A3(new_n657), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n514), .A2(new_n512), .A3(new_n658), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n660), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT29), .B(new_n671), .C1(new_n727), .C2(new_n656), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n722), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n698), .B1(new_n729), .B2(G1), .ZN(G364));
  NOR2_X1   g0530(.A1(new_n352), .A2(new_n280), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n251), .B1(new_n731), .B2(G45), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n694), .A2(KEYINPUT92), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  INV_X1    g0534(.A(new_n732), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n693), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n692), .A2(new_n325), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G355), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G116), .B2(new_n213), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n692), .A2(new_n380), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n448), .B2(new_n209), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n242), .A2(new_n448), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n273), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT93), .Z(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(G20), .B2(new_n294), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n738), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n352), .A2(KEYINPUT96), .A3(new_n288), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT96), .B1(new_n352), .B2(new_n288), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n371), .A2(G179), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT99), .Z(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n273), .A2(new_n288), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n325), .B1(new_n765), .B2(G87), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n352), .B1(new_n288), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n291), .A2(new_n205), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n766), .B1(new_n527), .B2(new_n770), .C1(new_n774), .C2(new_n307), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n771), .A2(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n771), .A2(KEYINPUT94), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(new_n371), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n775), .B1(G77), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n756), .A2(new_n768), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n409), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n785));
  NOR2_X1   g0585(.A1(new_n778), .A2(new_n288), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n784), .A2(new_n785), .B1(new_n786), .B2(G58), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT95), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n772), .B2(new_n288), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n771), .A2(KEYINPUT95), .A3(G190), .A4(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n783), .A2(new_n788), .B1(G50), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n762), .A2(new_n780), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n761), .A2(G283), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n258), .B1(new_n765), .B2(G303), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT33), .B(G317), .Z(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n583), .B2(new_n770), .C1(new_n774), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G329), .B2(new_n781), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n792), .A2(G326), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G311), .A2(new_n779), .B1(new_n786), .B2(G322), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n795), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n753), .B1(new_n803), .B2(new_n750), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n749), .B(KEYINPUT100), .Z(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n680), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n684), .A2(new_n737), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n680), .A2(G330), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G396));
  AND3_X1   g0609(.A1(new_n366), .A2(new_n367), .A3(new_n671), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n370), .A2(new_n372), .B1(new_n356), .B2(new_n671), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n368), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n659), .A2(new_n661), .ZN(new_n813));
  INV_X1    g0613(.A(new_n656), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n812), .B1(new_n815), .B2(new_n671), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT103), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n374), .A2(new_n671), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n662), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n818), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n815), .A2(KEYINPUT103), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n816), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n722), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n737), .B1(new_n822), .B2(new_n722), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n786), .A2(G143), .B1(G150), .B2(new_n773), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  INV_X1    g0627(.A(new_n792), .ZN(new_n828));
  INV_X1    g0628(.A(new_n779), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n826), .B1(new_n827), .B2(new_n828), .C1(new_n409), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT102), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n761), .A2(G68), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n380), .B1(new_n770), .B2(new_n414), .C1(new_n764), .C2(new_n283), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G132), .B2(new_n781), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n786), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n463), .A2(new_n829), .B1(new_n839), .B2(new_n583), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G303), .B2(new_n792), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n761), .A2(G87), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n258), .B1(new_n769), .B2(G97), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n361), .B2(new_n764), .C1(new_n774), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G311), .B2(new_n781), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  AOI21_X1  g0648(.A(new_n751), .B1(new_n838), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n747), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n751), .A2(new_n850), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n738), .B1(G77), .B2(new_n851), .C1(new_n812), .C2(new_n850), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n824), .A2(new_n825), .B1(new_n849), .B2(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n207), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OR3_X1    g0657(.A1(new_n208), .A2(new_n261), .A3(new_n415), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n283), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n251), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n423), .A2(new_n270), .ZN(new_n863));
  INV_X1    g0663(.A(new_n421), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n307), .B1(new_n864), .B2(new_n401), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT7), .B1(new_n380), .B2(G20), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n867), .B2(new_n418), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n432), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n445), .A2(new_n670), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n670), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n442), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n408), .A2(new_n869), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n433), .A2(new_n670), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n434), .A2(new_n876), .A3(new_n877), .A4(new_n442), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n862), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n870), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n877), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n445), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n878), .A2(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n434), .A2(new_n442), .A3(new_n877), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n878), .A2(KEYINPUT104), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n862), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n882), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n883), .B1(new_n893), .B2(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n638), .A2(new_n671), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n894), .A2(new_n895), .B1(new_n637), .B2(new_n670), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n314), .A2(new_n672), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n338), .A2(new_n341), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n314), .B(new_n672), .C1(new_n336), .C2(new_n337), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n821), .A2(new_n819), .ZN(new_n902));
  INV_X1    g0702(.A(new_n810), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n881), .A2(new_n882), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n896), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n728), .A2(new_n724), .A3(new_n446), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n907), .A2(new_n643), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(G330), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n900), .A2(new_n812), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n719), .B2(new_n699), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n892), .A2(new_n882), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n881), .B2(new_n882), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(KEYINPUT40), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n719), .A2(new_n699), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n446), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n910), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n251), .B2(new_n731), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n909), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n861), .B1(new_n923), .B2(new_n924), .ZN(G367));
  INV_X1    g0725(.A(new_n686), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n553), .B1(new_n549), .B2(new_n671), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n658), .A2(new_n672), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n688), .A2(new_n930), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  OAI21_X1  g0735(.A(new_n657), .B1(new_n927), .B2(new_n664), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n671), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n498), .A2(new_n671), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n655), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n649), .A2(new_n650), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n938), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT105), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(KEYINPUT105), .A3(new_n943), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n941), .A2(new_n942), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n937), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n933), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n946), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n949), .B(new_n933), .C1(new_n951), .C2(new_n944), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n932), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n949), .B1(new_n951), .B2(new_n944), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT106), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n931), .A3(new_n952), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n690), .A2(new_n930), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n688), .A2(new_n689), .A3(new_n929), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n926), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n688), .B1(new_n676), .B2(new_n687), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(new_n684), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n729), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n729), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n693), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n735), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n805), .B(new_n939), .C1(new_n940), .C2(new_n938), .ZN(new_n977));
  INV_X1    g0777(.A(new_n752), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n213), .B2(new_n354), .C1(new_n743), .C2(new_n238), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n401), .B1(new_n770), .B2(new_n361), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n764), .A2(new_n463), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(G294), .C2(new_n773), .ZN(new_n983));
  INV_X1    g0783(.A(new_n760), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n984), .A2(G97), .B1(G317), .B2(new_n781), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n792), .A2(G311), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G283), .A2(new_n779), .B1(new_n786), .B2(G303), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n985), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n782), .A2(new_n827), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n760), .A2(new_n261), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n774), .A2(new_n409), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n258), .B1(new_n770), .B2(new_n307), .C1(new_n764), .C2(new_n414), .ZN(new_n992));
  NOR4_X1   g0792(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n779), .A2(G50), .B1(G143), .B2(new_n792), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n272), .C2(new_n839), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI211_X1 g0797(.A(new_n738), .B(new_n979), .C1(new_n997), .C2(new_n751), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n958), .A2(new_n976), .B1(new_n977), .B2(new_n998), .ZN(G387));
  OR2_X1    g0799(.A1(new_n235), .A2(new_n448), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n695), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n1000), .A2(new_n742), .B1(new_n1001), .B2(new_n739), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n695), .B(new_n448), .C1(new_n307), .C2(new_n261), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n347), .B2(new_n283), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n277), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1002), .A2(new_n1007), .B1(G107), .B2(new_n213), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n737), .B1(new_n1008), .B2(new_n978), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n676), .B2(new_n805), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n764), .A2(new_n261), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n401), .B(new_n1011), .C1(new_n484), .C2(new_n769), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n277), .B2(new_n774), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G150), .B2(new_n781), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n792), .A2(G159), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n786), .B1(new_n779), .B2(G68), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n761), .A2(G97), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n779), .A2(G303), .B1(G311), .B2(new_n773), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n786), .A2(G317), .B1(G322), .B2(new_n792), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT48), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(KEYINPUT48), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n765), .A2(G294), .B1(G283), .B2(new_n769), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT107), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n380), .B1(new_n781), .B2(G326), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n463), .C2(new_n760), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1018), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1010), .B1(new_n1031), .B2(new_n750), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n969), .B2(new_n735), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n970), .A2(new_n693), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n729), .A2(new_n969), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(G393));
  NOR2_X1   g0836(.A1(new_n929), .A2(new_n749), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n743), .A2(new_n245), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n978), .B1(new_n213), .B2(new_n527), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n738), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n786), .A2(G311), .B1(G317), .B2(new_n792), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n325), .B1(new_n764), .B2(new_n844), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n781), .B2(G322), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n762), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n773), .A2(G303), .B1(G116), .B2(new_n769), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n829), .B2(new_n583), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT108), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n401), .B1(new_n765), .B2(G68), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n261), .B2(new_n770), .C1(new_n774), .C2(new_n283), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G143), .B2(new_n781), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n842), .B(new_n1052), .C1(new_n277), .C2(new_n829), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n786), .A2(G159), .B1(G150), .B2(new_n792), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1046), .A2(new_n1049), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT109), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1037), .B(new_n1040), .C1(new_n1057), .C2(new_n750), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n966), .B2(new_n735), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n972), .A2(new_n693), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n966), .A2(new_n971), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT110), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  INV_X1    g0869(.A(new_n895), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n893), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n811), .A2(new_n368), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n671), .B(new_n1072), .C1(new_n727), .C2(new_n656), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n903), .ZN(new_n1074));
  OAI211_X1 g0874(.A(KEYINPUT111), .B(new_n1071), .C1(new_n1074), .C2(new_n901), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT111), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n901), .B1(new_n1073), .B2(new_n903), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1071), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n894), .B1(new_n904), .B2(new_n1070), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n910), .B(new_n911), .C1(new_n699), .C2(new_n719), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n720), .A2(G330), .A3(new_n812), .A4(new_n900), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1080), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n918), .A2(G330), .A3(new_n812), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n901), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1089), .A2(new_n1085), .A3(new_n903), .A4(new_n1073), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n720), .A2(G330), .A3(new_n812), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1083), .B1(new_n1091), .B2(new_n901), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n810), .B1(new_n821), .B2(new_n819), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n446), .A2(new_n918), .A3(G330), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n907), .A2(new_n643), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT112), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1094), .A2(KEYINPUT112), .A3(new_n1096), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1087), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n693), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1080), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1083), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n735), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n894), .A2(new_n747), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n738), .B1(new_n347), .B2(new_n851), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n325), .B1(new_n769), .B2(G159), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n765), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT53), .B1(new_n765), .B2(G150), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1113), .B1(new_n774), .B2(new_n827), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n829), .A2(new_n1117), .B1(new_n1118), .B2(new_n828), .ZN(new_n1119));
  INV_X1    g0919(.A(G132), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n839), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n782), .A2(new_n1122), .B1(new_n760), .B2(new_n283), .ZN(new_n1123));
  OR4_X1    g0923(.A1(new_n1116), .A2(new_n1119), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n779), .A2(G97), .B1(G107), .B2(new_n773), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n844), .B2(new_n828), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT113), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n325), .B1(new_n770), .B2(new_n261), .C1(new_n764), .C2(new_n490), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n782), .A2(new_n583), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(G116), .C2(new_n786), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n835), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1124), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT114), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n751), .B1(new_n1134), .B2(KEYINPUT114), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1112), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT115), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1111), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1105), .A2(new_n1110), .A3(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT122), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n916), .B2(new_n910), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n915), .A2(new_n912), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT40), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n912), .B2(new_n913), .ZN(new_n1147));
  OAI211_X1 g0947(.A(KEYINPUT120), .B(G330), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n286), .A2(new_n670), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n297), .B(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1143), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n917), .A2(new_n1152), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n906), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n906), .A3(new_n1155), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1104), .B2(new_n1096), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1141), .B1(new_n1161), .B2(new_n694), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1096), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1109), .B2(new_n1101), .ZN(new_n1164));
  OAI211_X1 g0964(.A(KEYINPUT122), .B(new_n693), .C1(new_n1164), .C2(new_n1160), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1154), .A2(new_n1167), .A3(new_n1155), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(new_n1157), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1162), .A2(new_n1165), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n732), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1152), .A2(new_n747), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n738), .B1(G50), .B2(new_n851), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT119), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n984), .A2(G58), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT116), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n380), .A2(G41), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1179), .B(new_n1011), .C1(new_n781), .C2(G283), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT117), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n792), .A2(G116), .B1(G68), .B2(new_n769), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT118), .Z(new_n1184));
  OAI22_X1  g0984(.A1(new_n839), .A2(new_n361), .B1(new_n527), .B2(new_n774), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n484), .B2(new_n779), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT58), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G33), .A2(G41), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1178), .A2(G50), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n769), .A2(G150), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n764), .B2(new_n1117), .C1(new_n774), .C2(new_n1120), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G137), .B2(new_n779), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n1122), .B2(new_n828), .C1(new_n1118), .C2(new_n839), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n781), .A2(G124), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n1191), .C1(new_n409), .C2(new_n760), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1196), .B2(KEYINPUT59), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1192), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1189), .A2(new_n1190), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1175), .B1(new_n1202), .B2(new_n750), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1172), .B1(new_n1173), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1171), .A2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n901), .A2(new_n747), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n738), .B1(G68), .B2(new_n851), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n761), .A2(G77), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n258), .B1(new_n769), .B2(new_n484), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n527), .B2(new_n764), .C1(new_n774), .C2(new_n463), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G303), .B2(new_n781), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n792), .A2(G294), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G107), .A2(new_n779), .B1(new_n786), .B2(G283), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1208), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1177), .A2(new_n380), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT123), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n765), .A2(G159), .B1(G50), .B2(new_n769), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n774), .B2(new_n1117), .C1(new_n782), .C2(new_n1118), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G137), .B2(new_n786), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n779), .A2(G150), .B1(G132), .B2(new_n792), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1214), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1207), .B1(new_n1222), .B2(new_n750), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1094), .A2(new_n735), .B1(new_n1206), .B2(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1102), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1226), .B2(new_n974), .ZN(G381));
  INV_X1    g1027(.A(G375), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT124), .ZN(new_n1229));
  INV_X1    g1029(.A(G378), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(KEYINPUT124), .ZN(new_n1231));
  OR3_X1    g1031(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1233), .ZN(G407));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G407), .A2(new_n1237), .A3(G213), .ZN(G409));
  XOR2_X1   g1038(.A(G393), .B(G396), .Z(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(G387), .A2(new_n1066), .A3(new_n1064), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1068), .A2(G387), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G387), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1067), .B2(new_n1065), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1068), .A2(G387), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1239), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1243), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1171), .A2(G378), .A3(new_n1204), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1164), .A2(new_n974), .A3(new_n1169), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1158), .A2(new_n735), .A3(new_n1159), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1173), .A2(new_n1203), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1230), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1236), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1224), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1226), .A2(KEYINPUT60), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n694), .B1(new_n1225), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1257), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(G384), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(G384), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1264), .A2(KEYINPUT63), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1249), .B1(new_n1256), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT125), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1236), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1250), .A2(KEYINPUT125), .A3(new_n1255), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1236), .A2(G2897), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1262), .A2(new_n1263), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1272), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1269), .A2(new_n1270), .A3(new_n1264), .A4(new_n1271), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1266), .A2(new_n1276), .A3(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1248), .B1(new_n1281), .B2(new_n1256), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1277), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1256), .A2(KEYINPUT62), .A3(new_n1264), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1287), .B(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1280), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1280), .B(KEYINPUT127), .C1(new_n1286), .C2(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(G405));
  NOR2_X1   g1094(.A1(new_n1228), .A2(G378), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1250), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1297), .B(new_n1264), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(new_n1289), .ZN(G402));
endmodule


