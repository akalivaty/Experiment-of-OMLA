//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n207), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n219), .B1(new_n201), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n217), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(new_n207), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n211), .A2(G13), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT0), .Z(new_n237));
  NOR4_X1   g0037(.A1(new_n228), .A2(new_n229), .A3(new_n234), .A4(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n243));
  XNOR2_X1  g0043(.A(G226), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G238), .B(G244), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G77), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n256), .A2(KEYINPUT69), .A3(G222), .A4(new_n257), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n260), .A2(new_n266), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n270), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n271), .A2(G190), .A3(new_n278), .A4(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n280), .B1(new_n269), .B2(new_n270), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(KEYINPUT73), .A3(G190), .A4(new_n278), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G1), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n207), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n292), .A2(KEYINPUT70), .A3(new_n233), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT70), .B1(new_n292), .B2(new_n233), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n290), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n232), .A2(G1), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(G50), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n261), .B2(G20), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n232), .A2(KEYINPUT72), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(KEYINPUT8), .A2(G58), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT8), .A2(G58), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT71), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n308), .A3(new_n305), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n303), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G20), .A2(G33), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G150), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n232), .B1(new_n206), .B2(new_n207), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n310), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n295), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n291), .B(new_n299), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT9), .ZN(new_n319));
  INV_X1    g0119(.A(new_n314), .ZN(new_n320));
  INV_X1    g0120(.A(new_n315), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n307), .A2(new_n309), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n320), .B(new_n321), .C1(new_n322), .C2(new_n303), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n295), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT9), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n291), .A4(new_n299), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n284), .A2(new_n286), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n285), .A2(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT10), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n284), .A2(new_n286), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n319), .A2(new_n326), .ZN(new_n332));
  AND4_X1   g0132(.A1(KEYINPUT10), .A2(new_n331), .A3(new_n329), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n335));
  INV_X1    g0135(.A(G107), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n256), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n270), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n275), .A2(G244), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n281), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n289), .A2(G77), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G20), .A2(G77), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n344), .B1(new_n306), .B2(new_n312), .C1(new_n303), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n292), .A2(new_n233), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n347), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n298), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n214), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n341), .A2(new_n342), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n340), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n330), .A2(new_n333), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G20), .B1(G159), .B2(new_n311), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n256), .B2(G20), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT76), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n263), .A2(G33), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT7), .B(new_n232), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n366), .B2(new_n363), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT16), .B(new_n360), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n202), .B1(new_n362), .B2(new_n366), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n201), .A2(new_n202), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n206), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n311), .A2(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n347), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n213), .A2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n256), .B(new_n378), .C1(G223), .C2(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n272), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n272), .A2(G232), .A3(new_n274), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(new_n280), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G190), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n322), .A2(new_n297), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n296), .B1(new_n290), .B2(new_n322), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n379), .A2(new_n380), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n270), .ZN(new_n388));
  INV_X1    g0188(.A(new_n382), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n281), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n377), .A2(new_n384), .A3(new_n386), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n377), .A2(new_n386), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n383), .A2(G179), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n383), .B2(new_n354), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n272), .A2(G238), .A3(new_n274), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G226), .A2(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n220), .B2(G1698), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n256), .B1(G33), .B2(G97), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n404), .B(new_n281), .C1(new_n407), .C2(new_n272), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT13), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G200), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n220), .A2(G1698), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(G226), .B2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n413), .B2(new_n265), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n280), .B1(new_n414), .B2(new_n270), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT13), .A4(new_n404), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n202), .A2(G20), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n423), .B1(new_n207), .B2(new_n312), .C1(new_n303), .C2(new_n214), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n202), .B2(new_n350), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT11), .B1(new_n424), .B2(new_n295), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n423), .A2(G1), .A3(new_n287), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT12), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n410), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n421), .A2(G179), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT75), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n409), .A2(new_n435), .A3(G169), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT75), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n421), .A2(new_n437), .A3(G179), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n408), .B(new_n418), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT14), .B1(new_n439), .B2(new_n354), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n434), .A2(new_n436), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n430), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n318), .B1(new_n328), .B2(G179), .ZN(new_n444));
  AOI21_X1  g0244(.A(G169), .B1(new_n285), .B2(new_n278), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n348), .B1(new_n214), .B2(new_n350), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n341), .B2(G190), .ZN(new_n449));
  INV_X1    g0249(.A(G200), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(new_n341), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  AND4_X1   g0252(.A1(new_n358), .A2(new_n403), .A3(new_n443), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT78), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT78), .A2(G116), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(G33), .A3(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(G238), .A2(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n215), .A2(G1698), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n262), .A2(new_n459), .A3(new_n264), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n272), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n273), .A2(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n279), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n261), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(G250), .B(new_n463), .C1(new_n466), .C2(new_n233), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n462), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G190), .ZN(new_n470));
  INV_X1    g0270(.A(new_n464), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n461), .A2(new_n458), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n467), .C1(new_n472), .C2(new_n272), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G200), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n303), .B2(new_n224), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n256), .A2(new_n232), .A3(G68), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n232), .B1(new_n411), .B2(new_n475), .ZN(new_n478));
  INV_X1    g0278(.A(G87), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(new_n224), .A3(new_n336), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n347), .B1(new_n290), .B2(new_n345), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n273), .A2(G33), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n289), .B(new_n484), .C1(new_n293), .C2(new_n294), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G87), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n470), .A2(new_n474), .A3(new_n483), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n347), .ZN(new_n489));
  INV_X1    g0289(.A(new_n345), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n290), .A2(new_n345), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n469), .A2(new_n342), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n473), .A2(new_n354), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n262), .A2(new_n264), .A3(new_n232), .A4(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT22), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT22), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n256), .A2(new_n500), .A3(new_n232), .A4(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n456), .A2(new_n457), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n232), .A3(G33), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n336), .A2(G20), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT23), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT24), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n499), .B2(new_n501), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(new_n505), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n349), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n225), .A2(G1698), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n256), .B(new_n515), .C1(G250), .C2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n463), .ZN(new_n519));
  OR2_X1    g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  NAND2_X1  g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n270), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n518), .A2(new_n270), .B1(G264), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n463), .B1(new_n520), .B2(new_n521), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G274), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n450), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n506), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n288), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT25), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n486), .A2(G107), .B1(new_n531), .B2(new_n530), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NOR4_X1   g0334(.A1(new_n514), .A2(new_n527), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n524), .A2(new_n526), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G190), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n497), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT79), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n503), .A2(G20), .B1(new_n233), .B2(new_n292), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n542), .B(new_n232), .C1(G33), .C2(new_n224), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(KEYINPUT20), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n457), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT78), .A2(G116), .ZN(new_n546));
  OAI21_X1  g0346(.A(G20), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n347), .A3(new_n543), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT20), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n503), .A2(G20), .A3(new_n288), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n349), .A2(new_n289), .A3(G116), .A4(new_n484), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n523), .A2(G270), .B1(G274), .B2(new_n525), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n257), .A2(G257), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G264), .A2(G1698), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n256), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G303), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n265), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n560), .A3(new_n270), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n450), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n540), .B1(new_n554), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n522), .A2(new_n519), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n272), .A3(G270), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n561), .A2(new_n565), .A3(new_n526), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n565), .A3(new_n526), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  INV_X1    g0369(.A(new_n553), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n544), .B2(new_n550), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT79), .A4(new_n552), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n563), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n554), .A2(G179), .A3(new_n566), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n554), .A2(G169), .A3(new_n568), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n554), .A2(KEYINPUT21), .A3(G169), .A4(new_n568), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n573), .A2(new_n574), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n265), .B2(new_n215), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n542), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n256), .A2(G250), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n257), .B1(new_n584), .B2(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n270), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n523), .A2(G257), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n526), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT7), .B1(new_n265), .B2(new_n232), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n361), .B(G20), .C1(new_n262), .C2(new_n264), .ZN(new_n591));
  OAI21_X1  g0391(.A(G107), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n312), .A2(new_n214), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n224), .A2(new_n336), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G97), .A2(G107), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n336), .A2(KEYINPUT6), .A3(G97), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n592), .B(new_n594), .C1(new_n232), .C2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n347), .B1(G97), .B2(new_n486), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n290), .A2(new_n224), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT77), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n586), .A2(G190), .A3(new_n526), .A4(new_n587), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n589), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n588), .A2(new_n354), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n586), .A2(new_n342), .A3(new_n526), .A4(new_n587), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n486), .A2(G97), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n336), .B1(new_n362), .B2(new_n366), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n232), .B1(new_n598), .B2(new_n599), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n610), .A2(new_n593), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n604), .B(new_n609), .C1(new_n612), .C2(new_n349), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n579), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n509), .A2(KEYINPUT24), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n512), .B1(new_n511), .B2(new_n505), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n347), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n532), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n533), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n536), .A2(new_n354), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n537), .A2(new_n342), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n453), .A2(new_n539), .A3(new_n616), .A4(new_n624), .ZN(G372));
  AND3_X1   g0425(.A1(new_n577), .A2(new_n574), .A3(new_n578), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n624), .ZN(new_n627));
  INV_X1    g0427(.A(new_n615), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n539), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n496), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n488), .A2(new_n496), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n613), .A2(new_n608), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n631), .A2(KEYINPUT26), .A3(new_n607), .A4(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n614), .B2(new_n497), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n630), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n453), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g0438(.A(new_n638), .B(KEYINPUT80), .Z(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT82), .B1(new_n330), .B2(new_n333), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n331), .A2(new_n332), .A3(new_n329), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT10), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n327), .A2(KEYINPUT10), .A3(new_n329), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT82), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT81), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT18), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT18), .B1(new_n394), .B2(new_n396), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT81), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n441), .A2(new_n442), .B1(new_n357), .B2(new_n431), .ZN(new_n653));
  INV_X1    g0453(.A(new_n393), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n651), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n446), .B1(new_n647), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n639), .A2(new_n656), .ZN(G369));
  NOR2_X1   g0457(.A1(new_n287), .A2(G20), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n273), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n626), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT84), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT83), .B1(new_n624), .B2(new_n664), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n514), .A2(new_n532), .A3(new_n534), .ZN(new_n669));
  INV_X1    g0469(.A(new_n527), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n538), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n621), .A2(new_n664), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n668), .B1(new_n673), .B2(new_n624), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n624), .A3(new_n672), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT83), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n667), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n673), .A2(new_n624), .ZN(new_n680));
  OAI211_X1 g0480(.A(KEYINPUT84), .B(new_n679), .C1(new_n680), .C2(new_n668), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n666), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n624), .A2(new_n664), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n681), .ZN(new_n685));
  INV_X1    g0485(.A(new_n626), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n554), .A2(new_n664), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n579), .B2(new_n687), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n684), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n235), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n480), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n231), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI211_X1 g0501(.A(KEYINPUT29), .B(new_n664), .C1(new_n629), .C2(new_n636), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n606), .A2(KEYINPUT86), .A3(new_n614), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT86), .B1(new_n606), .B2(new_n614), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n627), .B(new_n539), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n636), .ZN(new_n707));
  INV_X1    g0507(.A(new_n664), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n586), .A2(new_n526), .A3(new_n587), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n473), .A2(new_n568), .A3(new_n342), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n524), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n566), .A2(G179), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n588), .A2(new_n713), .A3(new_n536), .A4(new_n473), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n586), .A2(new_n524), .A3(new_n526), .A4(new_n587), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n566), .A2(new_n469), .A3(G179), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT31), .B1(new_n719), .B2(new_n664), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT85), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n616), .A2(new_n539), .A3(new_n624), .A4(new_n708), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n720), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n722), .B(new_n723), .C1(new_n725), .C2(KEYINPUT85), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n702), .B(new_n709), .C1(G330), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n701), .B1(new_n727), .B2(G1), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT87), .Z(G364));
  INV_X1    g0529(.A(new_n692), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n658), .A2(G45), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n697), .A2(G1), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n690), .A2(new_n691), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n233), .B1(G20), .B2(new_n354), .ZN(new_n735));
  INV_X1    g0535(.A(G190), .ZN(new_n736));
  NOR4_X1   g0536(.A1(new_n232), .A2(new_n736), .A3(new_n450), .A4(G179), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT91), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n256), .B1(new_n739), .B2(G303), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G179), .A2(G200), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n232), .B1(new_n741), .B2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G294), .ZN(new_n744));
  NAND2_X1  g0544(.A1(G20), .A2(G179), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT89), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G322), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n736), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n450), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G311), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n740), .A2(new_n744), .A3(new_n749), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n736), .A2(G20), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT90), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(G179), .A3(new_n450), .ZN(new_n759));
  INV_X1    g0559(.A(new_n741), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G283), .B1(new_n761), .B2(G329), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  NOR2_X1   g0563(.A1(new_n747), .A2(new_n450), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n755), .B(new_n763), .C1(G326), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n737), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n256), .B1(new_n742), .B2(new_n224), .C1(new_n766), .C2(new_n479), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT32), .ZN(new_n768));
  INV_X1    g0568(.A(new_n761), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n761), .A2(KEYINPUT32), .A3(G159), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G68), .A2(new_n752), .B1(new_n751), .B2(G77), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G107), .A2(new_n759), .B1(new_n764), .B2(G50), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G58), .B2(new_n748), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n735), .B1(new_n765), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n778), .B1(new_n689), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n695), .A2(new_n256), .ZN(new_n784));
  INV_X1    g0584(.A(G45), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n230), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n784), .B(new_n786), .C1(new_n251), .C2(new_n785), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n256), .A2(G355), .A3(new_n235), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(G116), .C2(new_n235), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n781), .A2(new_n735), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n732), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT88), .Z(new_n792));
  OAI21_X1  g0592(.A(new_n734), .B1(new_n783), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  NAND2_X1  g0596(.A1(new_n637), .A2(new_n708), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n356), .A2(new_n664), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n448), .A2(new_n664), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n451), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n801), .B2(new_n357), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n357), .B1(new_n451), .B2(new_n800), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n798), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n637), .A2(new_n805), .A3(new_n708), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n726), .A2(G330), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n807), .B(new_n808), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n732), .ZN(new_n810));
  INV_X1    g0610(.A(new_n759), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n202), .B1(new_n769), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n256), .B1(new_n738), .B2(new_n207), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G143), .A2(new_n748), .B1(new_n752), .B2(G150), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  INV_X1    g0616(.A(new_n764), .ZN(new_n817));
  INV_X1    g0617(.A(new_n751), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n770), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n813), .B(new_n814), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n201), .B2(new_n742), .C1(new_n820), .C2(new_n819), .ZN(new_n822));
  INV_X1    g0622(.A(new_n748), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n752), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT95), .B(G283), .Z(new_n827));
  OAI22_X1  g0627(.A1(new_n559), .A2(new_n817), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n504), .B2(new_n751), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n759), .A2(G87), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n769), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G107), .B2(new_n739), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n256), .B1(new_n743), .B2(G97), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n822), .B1(new_n825), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n735), .A2(new_n779), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(new_n735), .B1(new_n214), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n732), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n838), .B(new_n839), .C1(new_n780), .C2(new_n805), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n810), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT35), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n232), .B(new_n233), .C1(new_n600), .C2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(G116), .C1(new_n842), .C2(new_n600), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n231), .A2(new_n214), .A3(new_n372), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT97), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT97), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT98), .B1(new_n202), .B2(G50), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n202), .A2(KEYINPUT98), .A3(G50), .ZN(new_n851));
  OAI211_X1 g0651(.A(G1), .B(new_n287), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n723), .A2(new_n725), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n441), .A2(new_n442), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n442), .A2(new_n664), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n431), .A3(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n442), .B(new_n664), .C1(new_n441), .C2(new_n432), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n855), .A2(new_n805), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n280), .B1(new_n387), .B2(new_n270), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n354), .B1(new_n863), .B2(new_n389), .ZN(new_n864));
  NOR4_X1   g0664(.A1(new_n381), .A2(new_n382), .A3(new_n342), .A4(new_n280), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n360), .B1(new_n367), .B2(new_n368), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n370), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n295), .A3(new_n369), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n869), .B2(new_n386), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n384), .A2(new_n377), .A3(new_n386), .A4(new_n391), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n202), .B1(new_n591), .B2(KEYINPUT76), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n375), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n295), .B1(new_n875), .B2(KEYINPUT16), .ZN(new_n876));
  INV_X1    g0676(.A(new_n369), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n386), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT100), .ZN(new_n879));
  INV_X1    g0679(.A(new_n662), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n385), .A2(new_n296), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n322), .A2(new_n290), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n317), .B1(new_n867), .B2(new_n370), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(new_n369), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT100), .B1(new_n886), .B2(new_n662), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT101), .B(new_n392), .C1(new_n886), .C2(new_n866), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n872), .A2(new_n881), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n394), .A2(new_n880), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n397), .A2(new_n891), .A3(new_n392), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n393), .A2(new_n401), .B1(new_n881), .B2(new_n887), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n893), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n899), .A2(new_n900), .A3(new_n896), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n861), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n651), .A2(new_n652), .A3(new_n393), .ZN(new_n905));
  INV_X1    g0705(.A(new_n891), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n892), .B(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n861), .B(KEYINPUT40), .C1(new_n901), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n453), .A2(new_n855), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n911), .B(new_n912), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(G330), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n901), .B2(new_n909), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n856), .A2(new_n664), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  INV_X1    g0718(.A(new_n888), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n878), .A2(new_n396), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT101), .B1(new_n920), .B2(new_n392), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n887), .A2(new_n881), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n918), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(KEYINPUT38), .B(new_n897), .C1(new_n925), .C2(new_n893), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n900), .B1(new_n899), .B2(new_n896), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT39), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n916), .A2(new_n917), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n651), .A2(new_n652), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n662), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n806), .A2(new_n799), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n860), .B(new_n932), .C1(new_n898), .C2(new_n901), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n453), .B1(new_n709), .B2(new_n702), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n656), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n914), .B(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n658), .A2(new_n273), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n854), .B1(new_n938), .B2(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n613), .A2(new_n664), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n704), .B2(new_n705), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(new_n624), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n664), .B1(new_n943), .B2(new_n614), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n632), .A2(new_n607), .A3(new_n664), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n682), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT42), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n946), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n483), .A2(new_n487), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n664), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n631), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n496), .B2(new_n953), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(KEYINPUT102), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n951), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n946), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n693), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n951), .A2(new_n959), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n960), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n696), .B(KEYINPUT41), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n685), .A2(new_n665), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n969), .A2(new_n730), .A3(new_n682), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n730), .B1(new_n969), .B2(new_n682), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n727), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT103), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n693), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT44), .B1(new_n684), .B2(new_n946), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(new_n961), .C1(new_n682), .C2(new_n683), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT45), .B1(new_n684), .B2(new_n946), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n682), .A2(new_n979), .A3(new_n683), .A4(new_n961), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n975), .B(new_n977), .C1(new_n978), .C2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n693), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(KEYINPUT103), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n975), .A2(new_n977), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n684), .A2(new_n946), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n979), .ZN(new_n986));
  INV_X1    g0786(.A(new_n980), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n988), .A3(new_n693), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n974), .A2(new_n983), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n968), .B1(new_n990), .B2(new_n727), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n731), .A2(G1), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n966), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n256), .B1(new_n766), .B2(new_n201), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n811), .A2(new_n214), .B1(new_n769), .B2(new_n816), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G68), .C2(new_n743), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n207), .A2(new_n818), .B1(new_n823), .B2(new_n313), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G143), .B2(new_n764), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(new_n770), .C2(new_n826), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n742), .A2(new_n336), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n831), .A2(new_n817), .B1(new_n818), .B2(new_n827), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G303), .B2(new_n748), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n759), .A2(G97), .B1(new_n761), .B2(G317), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n738), .A2(new_n455), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT46), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT46), .B1(new_n737), .B2(new_n504), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n256), .B(new_n1006), .C1(new_n752), .C2(G294), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n999), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n732), .B1(new_n1010), .B2(new_n735), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n784), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n790), .B1(new_n235), .B2(new_n345), .C1(new_n241), .C2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(new_n782), .C2(new_n955), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n993), .A2(new_n1014), .ZN(G387));
  AND2_X1   g0815(.A1(new_n761), .A2(G326), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G311), .A2(new_n752), .B1(new_n748), .B2(G317), .ZN(new_n1017));
  INV_X1    g0817(.A(G322), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n559), .B2(new_n818), .C1(new_n1018), .C2(new_n817), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n824), .B2(new_n766), .C1(new_n742), .C2(new_n827), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n256), .B(new_n1016), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n1022), .B2(new_n1021), .C1(new_n503), .C2(new_n811), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n322), .A2(new_n826), .B1(new_n818), .B2(new_n202), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT106), .Z(new_n1026));
  NAND2_X1  g0826(.A1(new_n743), .A2(new_n490), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n256), .C1(new_n766), .C2(new_n214), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n811), .A2(new_n224), .B1(new_n769), .B2(new_n313), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G159), .C2(new_n764), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1026), .B(new_n1030), .C1(new_n207), .C2(new_n823), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n698), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n304), .A2(new_n207), .A3(new_n305), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(KEYINPUT50), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n785), .C1(KEYINPUT50), .C2(new_n1034), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n202), .A2(new_n214), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n784), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT104), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n785), .B2(new_n247), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1033), .A2(new_n235), .A3(new_n256), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G107), .C2(new_n235), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT105), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n781), .B(new_n735), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1032), .A2(new_n735), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n685), .B2(new_n782), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n732), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n970), .A2(new_n971), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1048), .B1(new_n992), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n727), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(new_n696), .A3(new_n972), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(G393));
  AOI21_X1  g0853(.A(new_n693), .B1(new_n984), .B2(new_n988), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n981), .A2(new_n982), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n972), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n696), .A3(new_n990), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G311), .A2(new_n748), .B1(new_n764), .B2(G317), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n265), .B1(new_n766), .B2(new_n827), .C1(new_n818), .C2(new_n824), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n752), .A2(G303), .B1(new_n504), .B2(new_n743), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT109), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n811), .A2(new_n336), .B1(new_n769), .B2(new_n1018), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1061), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(KEYINPUT109), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1059), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n761), .A2(G143), .B1(G68), .B2(new_n737), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT108), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n830), .B1(new_n826), .B2(new_n207), .C1(new_n306), .C2(new_n818), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n764), .B1(new_n748), .B2(G159), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT107), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1069), .B(new_n1070), .C1(new_n1072), .C2(KEYINPUT51), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(KEYINPUT51), .B2(new_n1072), .C1(new_n214), .C2(new_n742), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1074), .B2(new_n265), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n732), .B1(new_n1075), .B2(new_n735), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n790), .B1(new_n224), .B2(new_n235), .C1(new_n254), .C2(new_n1012), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n961), .A2(new_n781), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n992), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1057), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT110), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1057), .A2(new_n1081), .A3(KEYINPUT110), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(G390));
  NAND3_X1  g0886(.A1(new_n453), .A2(G330), .A3(new_n855), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n935), .A2(new_n1087), .A3(new_n656), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT111), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n802), .A2(new_n691), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n860), .B1(new_n726), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1091), .A2(new_n855), .A3(new_n860), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n932), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n664), .B(new_n804), .C1(new_n706), .C2(new_n636), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n798), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n726), .A2(new_n860), .A3(new_n1091), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1091), .A2(new_n855), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n860), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n935), .A2(new_n1087), .A3(KEYINPUT111), .A4(new_n656), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1090), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n917), .B1(new_n932), .B2(new_n860), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n916), .B2(new_n928), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n907), .A2(new_n908), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n900), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n926), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n860), .B1(new_n1095), .B2(new_n798), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n917), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1106), .A2(new_n1112), .A3(new_n1097), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n806), .A2(new_n799), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1114), .B2(new_n1099), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT39), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT39), .B1(new_n1108), .B2(new_n926), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1093), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1104), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1106), .A2(new_n1112), .B1(new_n1099), .B2(new_n1098), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1097), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1090), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(new_n696), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n780), .B1(new_n916), .B2(new_n928), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n761), .A2(G125), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n256), .B(new_n1129), .C1(new_n811), .C2(new_n207), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT112), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n737), .A2(G150), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1132), .A2(KEYINPUT53), .B1(G159), .B2(new_n743), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(KEYINPUT53), .B2(new_n1132), .C1(new_n817), .C2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n812), .A2(new_n823), .B1(new_n818), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1131), .B(new_n1138), .C1(new_n816), .C2(new_n826), .ZN(new_n1139));
  INV_X1    g0939(.A(G283), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n817), .A2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n336), .A2(new_n826), .B1(new_n823), .B2(new_n455), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G97), .B2(new_n751), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n256), .B1(new_n759), .B2(G68), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n824), .A2(new_n769), .B1(new_n738), .B2(new_n479), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G77), .B2(new_n743), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1139), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(new_n735), .B1(new_n322), .B2(new_n837), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1128), .A2(new_n732), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n992), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1127), .A2(KEYINPUT113), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT113), .B1(new_n1127), .B2(new_n1153), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1154), .A2(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n855), .A2(new_n860), .A3(new_n805), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n926), .B2(new_n927), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n910), .B(G330), .C1(new_n1159), .C2(KEYINPUT40), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n318), .A2(new_n880), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT56), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT55), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n647), .B2(new_n447), .ZN(new_n1165));
  AOI211_X1 g0965(.A(KEYINPUT55), .B(new_n446), .C1(new_n640), .C2(new_n646), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT82), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n645), .B1(new_n643), .B2(new_n644), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n447), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT55), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n647), .A2(new_n1164), .A3(new_n447), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n1162), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1160), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n904), .A2(G330), .A3(new_n910), .A4(new_n1174), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n934), .A2(KEYINPUT118), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1176), .A2(new_n1177), .A3(new_n934), .A4(KEYINPUT118), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1090), .A2(new_n1103), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1152), .B2(new_n1102), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1157), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1183), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1121), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1178), .A2(new_n934), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n934), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n1191), .A3(KEYINPUT57), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1185), .A2(new_n1192), .A3(new_n696), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1180), .A2(new_n992), .A3(new_n1181), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n261), .A2(new_n465), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT114), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n207), .C1(G41), .C2(new_n256), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT115), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G116), .A2(new_n764), .B1(new_n751), .B2(new_n490), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n224), .B2(new_n826), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n811), .A2(new_n201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1202), .A2(G41), .A3(new_n256), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n737), .A2(G77), .B1(new_n743), .B2(G68), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n1140), .C2(new_n769), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1201), .B(new_n1205), .C1(G107), .C2(new_n748), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1199), .B1(new_n1206), .B2(KEYINPUT58), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(KEYINPUT58), .B2(new_n1206), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n811), .A2(new_n770), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G132), .A2(new_n752), .B1(new_n751), .B2(G137), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT116), .Z(new_n1211));
  OAI22_X1  g1011(.A1(new_n823), .A2(new_n1134), .B1(new_n313), .B2(new_n742), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G125), .B2(new_n764), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n766), .C2(new_n1136), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1196), .B(new_n1209), .C1(new_n1214), .C2(KEYINPUT59), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT117), .B(G124), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1215), .B1(KEYINPUT59), .B2(new_n1214), .C1(new_n769), .C2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1208), .B(new_n1217), .C1(new_n1198), .C2(new_n1197), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1218), .A2(new_n735), .B1(new_n207), .B2(new_n837), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n839), .C1(new_n780), .C2(new_n1174), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1194), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1193), .A2(new_n1221), .ZN(G375));
  AOI21_X1  g1022(.A(new_n732), .B1(new_n202), .B2(new_n837), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n860), .A2(new_n780), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n812), .A2(new_n817), .B1(new_n826), .B2(new_n1136), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G137), .B2(new_n748), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1134), .A2(new_n769), .B1(new_n738), .B2(new_n770), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(new_n1202), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n751), .A2(G150), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n265), .B1(new_n743), .B2(G50), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G294), .A2(new_n764), .B1(new_n752), .B2(new_n504), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n336), .B2(new_n818), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT122), .Z(new_n1235));
  OAI221_X1 g1035(.A(new_n265), .B1(new_n769), .B2(new_n559), .C1(new_n811), .C2(new_n214), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1027), .B1(new_n823), .B2(new_n1140), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(KEYINPUT123), .B2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1235), .B(new_n1238), .C1(KEYINPUT123), .C2(new_n1237), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n738), .A2(new_n224), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1232), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1224), .B(new_n1225), .C1(new_n735), .C2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n992), .ZN(new_n1244));
  OR3_X1    g1044(.A1(new_n1243), .A2(KEYINPUT120), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT120), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1183), .A2(new_n1243), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n967), .B(KEYINPUT119), .Z(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1125), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(G381));
  INV_X1    g1052(.A(G375), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1127), .A2(new_n1153), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(G384), .A3(G381), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1084), .A2(new_n1014), .A3(new_n993), .A4(new_n1085), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1050), .A2(new_n795), .A3(new_n1052), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(G407));
  NAND2_X1  g1060(.A1(new_n663), .A2(G213), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT124), .Z(new_n1262));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(new_n1255), .C2(new_n1262), .ZN(G409));
  AOI21_X1  g1063(.A(KEYINPUT110), .B1(new_n1057), .B2(new_n1081), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1085), .ZN(new_n1265));
  OAI21_X1  g1065(.A(G387), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1257), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G393), .A2(G396), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1258), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1266), .A2(new_n1257), .A3(new_n1267), .A4(new_n1270), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1193), .B(new_n1221), .C1(new_n1155), .C2(new_n1154), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1191), .A2(new_n992), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1187), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1220), .B(new_n1276), .C1(new_n1277), .C2(new_n1249), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1254), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n696), .B(new_n1125), .C1(new_n1248), .C2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT60), .B1(new_n1183), .B2(new_n1243), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1247), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n810), .A3(new_n840), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1247), .B(G384), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1280), .A2(new_n1261), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1262), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(G2897), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1261), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1292), .A2(G2897), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1287), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1261), .B2(new_n1280), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1289), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1290), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1288), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1274), .A2(new_n1297), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  XOR2_X1   g1101(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1292), .B(new_n1287), .C1(new_n1275), .C2(new_n1279), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT127), .B1(new_n1304), .B2(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1289), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1299), .A2(KEYINPUT62), .A3(new_n1288), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1303), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1301), .B1(new_n1311), .B2(new_n1274), .ZN(G405));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1254), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1275), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1272), .A2(new_n1273), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1287), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1314), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1272), .A2(new_n1273), .A3(new_n1314), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1288), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1322), .ZN(G402));
endmodule


