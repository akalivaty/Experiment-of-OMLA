//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(G50), .ZN(new_n226));
  AND2_X1   g0026(.A1(KEYINPUT64), .A2(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(KEYINPUT64), .A2(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n208), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT0), .Z(new_n234));
  NOR4_X1   g0034(.A1(new_n224), .A2(new_n225), .A3(new_n231), .A4(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  OAI21_X1  g0052(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n206), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n229), .A2(G33), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n230), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(new_n205), .B2(G20), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n265), .A2(new_n267), .B1(new_n266), .B2(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G222), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n272), .B1(new_n216), .B2(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G274), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n282), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(G226), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G200), .ZN(new_n288));
  INV_X1    g0088(.A(new_n287), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G190), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n270), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT70), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n269), .B1(new_n289), .B2(G169), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n293), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n291), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n294), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n274), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n277), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n283), .B1(G238), .B2(new_n285), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT14), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n314), .B2(G179), .ZN(new_n320));
  NOR4_X1   g0120(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT71), .A4(new_n297), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n316), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n261), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n229), .A2(G33), .A3(G77), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G20), .A2(G33), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n264), .B2(new_n261), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n205), .A2(G20), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n263), .A2(KEYINPUT69), .A3(new_n230), .A4(new_n260), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n330), .A2(G68), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n264), .A2(new_n210), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT12), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n328), .A2(new_n333), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n322), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n314), .A2(G190), .ZN(new_n339));
  INV_X1    g0139(.A(new_n337), .ZN(new_n340));
  OAI21_X1  g0140(.A(G200), .B1(new_n312), .B2(new_n313), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT7), .B1(new_n271), .B2(G20), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT7), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n229), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n344), .A2(new_n349), .A3(G68), .ZN(new_n350));
  INV_X1    g0150(.A(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n210), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n201), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n325), .A2(G159), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n353), .A2(KEYINPUT16), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n261), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT64), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n206), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT64), .A2(G20), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT7), .B1(new_n361), .B2(new_n271), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n347), .A2(new_n348), .A3(new_n206), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G68), .A3(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n353), .A2(new_n354), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT16), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT72), .B1(new_n357), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n323), .B1(new_n350), .B2(new_n355), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n364), .A2(new_n365), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(KEYINPUT16), .ZN(new_n371));
  INV_X1    g0171(.A(new_n258), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n265), .A2(new_n331), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n258), .A2(new_n264), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT73), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n367), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n307), .A2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n271), .B(new_n378), .C1(G223), .C2(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n280), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n237), .A2(new_n284), .B1(new_n281), .B2(new_n282), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n315), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n381), .A2(new_n297), .A3(new_n382), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT18), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n377), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n371), .A2(new_n376), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G200), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n381), .B2(new_n382), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n367), .A4(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n367), .A2(new_n397), .A3(new_n371), .A4(new_n376), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n389), .A2(new_n391), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n258), .B1(KEYINPUT68), .B2(new_n256), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(KEYINPUT68), .B2(new_n256), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n216), .B2(new_n229), .C1(new_n257), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n261), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n330), .A2(G77), .A3(new_n331), .A4(new_n332), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(G77), .C2(new_n263), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n271), .A2(G232), .A3(new_n273), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n271), .A2(G238), .A3(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n218), .C2(new_n271), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n277), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n283), .B1(G244), .B2(new_n285), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n393), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n415), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n395), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n297), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n315), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NOR4_X1   g0223(.A1(new_n304), .A2(new_n343), .A3(new_n402), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n211), .A2(new_n273), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n217), .A2(G1698), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n345), .C2(new_n346), .ZN(new_n427));
  INV_X1    g0227(.A(G116), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n255), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n277), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT76), .ZN(new_n433));
  INV_X1    g0233(.A(G45), .ZN(new_n434));
  OAI21_X1  g0234(.A(G250), .B1(new_n434), .B2(G1), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n277), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n280), .A3(KEYINPUT76), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n434), .A2(G1), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n280), .A2(G274), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n432), .A2(new_n439), .A3(new_n297), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT77), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n359), .A2(G33), .A3(G97), .A4(new_n360), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT19), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n229), .A2(new_n271), .A3(G68), .ZN(new_n447));
  NAND3_X1  g0247(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n359), .A2(new_n360), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G97), .A2(G107), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n212), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n446), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n261), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n405), .A2(new_n264), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT78), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n405), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n205), .A2(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n405), .A2(new_n456), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n457), .A2(new_n265), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G238), .A2(G1698), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n217), .B2(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n429), .B1(new_n463), .B2(new_n271), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n441), .B1(new_n464), .B2(new_n280), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n436), .A2(new_n438), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n315), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n281), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n431), .A2(new_n277), .B1(new_n468), .B2(new_n440), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT77), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n297), .A4(new_n439), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n443), .A2(new_n461), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n432), .A2(new_n439), .A3(new_n441), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G200), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n453), .A2(new_n261), .B1(new_n264), .B2(new_n405), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n265), .A2(new_n458), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G87), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n469), .A2(G190), .A3(new_n439), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n474), .A2(new_n475), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT79), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n218), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT25), .B1(new_n264), .B2(new_n218), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n476), .A2(new_n218), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n359), .B(new_n360), .C1(new_n345), .C2(new_n346), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT22), .B1(new_n489), .B2(new_n212), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n229), .A2(new_n271), .A3(new_n491), .A4(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n361), .A2(new_n494), .A3(new_n218), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT23), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n206), .B1(new_n429), .B2(KEYINPUT23), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT24), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n493), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n488), .B1(new_n503), .B2(new_n261), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n440), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G264), .A3(new_n280), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT5), .B(G41), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(G274), .A3(new_n280), .A4(new_n440), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G250), .A2(G1698), .ZN(new_n512));
  INV_X1    g0312(.A(G257), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(G1698), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n271), .B1(G33), .B2(G294), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n509), .B(new_n511), .C1(new_n515), .C2(new_n280), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n395), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT81), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT81), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n519), .A3(new_n395), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n518), .B(new_n520), .C1(G190), .C2(new_n516), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n504), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n516), .A2(G179), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n315), .B2(new_n516), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n323), .B1(new_n500), .B2(new_n502), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n488), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  AND2_X1   g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n450), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n218), .A2(KEYINPUT6), .A3(G97), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n229), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT74), .B1(new_n256), .B2(new_n216), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT74), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n325), .A2(new_n534), .A3(G77), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n362), .A2(G107), .A3(new_n363), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n261), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n263), .A2(G97), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G97), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n476), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(new_n273), .C1(new_n345), .C2(new_n346), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G250), .A2(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(KEYINPUT4), .A2(G244), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n271), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n277), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n508), .A2(G257), .A3(new_n280), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n558), .A2(new_n511), .ZN(new_n559));
  AOI21_X1  g0359(.A(G169), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n280), .B1(new_n549), .B2(new_n555), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n558), .A2(new_n511), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n562), .A2(new_n563), .A3(G179), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n546), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n395), .B1(new_n562), .B2(new_n563), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n557), .A2(new_n559), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(G190), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT75), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n544), .B1(new_n539), .B2(new_n261), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n566), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n273), .A2(G264), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G257), .A2(G1698), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(new_n345), .B2(new_n346), .ZN(new_n577));
  OR2_X1    g0377(.A1(KEYINPUT3), .A2(G33), .ZN(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  NAND2_X1  g0379(.A1(KEYINPUT3), .A2(G33), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n577), .A2(KEYINPUT80), .A3(new_n277), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n508), .A2(G270), .A3(new_n280), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(new_n511), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n277), .ZN(new_n586));
  INV_X1    g0386(.A(new_n576), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n219), .A2(G1698), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n578), .B2(new_n580), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n585), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n315), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n428), .B1(new_n205), .B2(G33), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n330), .A2(new_n332), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n264), .A2(new_n428), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n255), .A2(G97), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n359), .A2(new_n595), .A3(new_n360), .A4(new_n550), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n260), .A2(new_n230), .B1(G20), .B2(new_n428), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n593), .B(new_n594), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n590), .A2(new_n511), .A3(new_n582), .A4(new_n583), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n604), .B2(G200), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n393), .B2(new_n604), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n600), .A2(new_n584), .A3(G179), .A4(new_n590), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n600), .A2(new_n604), .A3(KEYINPUT21), .A4(G169), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n603), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n574), .A2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n424), .A2(new_n485), .A3(new_n527), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n300), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n377), .A2(new_n387), .A3(new_n390), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n390), .B1(new_n377), .B2(new_n387), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n342), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n338), .B1(new_n616), .B2(new_n422), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n399), .B(KEYINPUT17), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n617), .A2(new_n618), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n294), .A2(new_n303), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n612), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n461), .A2(new_n467), .A3(new_n442), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n480), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n629), .B2(new_n566), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n571), .A2(new_n560), .A3(new_n564), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n482), .A2(new_n484), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g0432(.A(KEYINPUT82), .B(KEYINPUT26), .Z(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT21), .B1(new_n591), .B2(new_n600), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n608), .A2(new_n607), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n526), .ZN(new_n638));
  AOI21_X1  g0438(.A(G200), .B1(new_n557), .B2(new_n559), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n562), .A2(new_n563), .A3(G190), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT75), .B1(new_n641), .B2(new_n546), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n569), .A2(new_n571), .A3(new_n570), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n631), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n629), .B1(new_n504), .B2(new_n521), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n638), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n634), .A2(new_n628), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n424), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n626), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G13), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G1), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n229), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT84), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n229), .A2(KEYINPUT84), .A3(new_n651), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n654), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT85), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n654), .A2(new_n656), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT85), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(G213), .A4(new_n657), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT86), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT86), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n660), .A2(new_n664), .A3(new_n668), .A4(G343), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n600), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(KEYINPUT87), .A3(new_n600), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n637), .A3(new_n606), .A4(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n637), .ZN(new_n677));
  XNOR2_X1  g0477(.A(KEYINPUT88), .B(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n504), .B1(new_n667), .B2(new_n669), .ZN(new_n680));
  INV_X1    g0480(.A(new_n522), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n526), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n670), .ZN(new_n683));
  INV_X1    g0483(.A(new_n526), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n677), .A2(new_n679), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n670), .A2(new_n637), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n682), .A2(new_n688), .B1(new_n684), .B2(new_n683), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(G41), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n232), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n451), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n226), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n646), .A2(new_n628), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n629), .A2(new_n566), .A3(new_n627), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n632), .B2(new_n633), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n683), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT91), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT91), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n703), .B(new_n683), .C1(new_n698), .C2(new_n700), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n697), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  AOI211_X1 g0507(.A(KEYINPUT92), .B(new_n707), .C1(new_n702), .C2(new_n704), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n647), .A2(KEYINPUT90), .A3(new_n683), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT90), .B1(new_n647), .B2(new_n683), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n707), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n610), .A2(new_n485), .A3(new_n527), .A4(new_n683), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n509), .B1(new_n515), .B2(new_n280), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n473), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n582), .A2(new_n511), .A3(new_n583), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n280), .B1(new_n347), .B2(new_n579), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT80), .B1(new_n720), .B2(new_n577), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n719), .A2(new_n721), .A3(new_n297), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n562), .A2(new_n563), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(KEYINPUT89), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(G179), .B1(new_n469), .B2(new_n439), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n568), .A3(new_n516), .A4(new_n604), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT89), .B1(new_n724), .B2(new_n725), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n716), .B1(new_n732), .B2(new_n683), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n724), .A2(new_n725), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n670), .B(KEYINPUT31), .C1(new_n734), .C2(new_n730), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n715), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n679), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n714), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n696), .B1(new_n738), .B2(new_n205), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT93), .Z(G364));
  NOR2_X1   g0540(.A1(new_n361), .A2(new_n650), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G45), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n692), .A2(new_n742), .A3(G1), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n677), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n230), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT95), .ZN(new_n750));
  OAI21_X1  g0550(.A(G20), .B1(new_n750), .B2(G169), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n315), .A2(KEYINPUT95), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n746), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n248), .A2(G45), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n232), .A2(new_n347), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n759), .B(new_n761), .C1(G45), .C2(new_n226), .ZN(new_n762));
  INV_X1    g0562(.A(new_n232), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n347), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G355), .B1(new_n428), .B2(new_n763), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n758), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n361), .A2(G179), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n393), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n393), .A3(G200), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n266), .B1(new_n210), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n361), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n543), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n361), .A2(new_n393), .A3(new_n774), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  OAI21_X1  g0581(.A(KEYINPUT32), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n395), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n361), .A2(new_n393), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G107), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(G20), .A3(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n347), .B1(new_n788), .B2(G87), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n779), .A2(new_n782), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n780), .A2(KEYINPUT32), .A3(new_n781), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n773), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n767), .A2(KEYINPUT97), .ZN(new_n793));
  AOI21_X1  g0593(.A(G200), .B1(new_n767), .B2(KEYINPUT97), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n793), .A2(G190), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n793), .A2(new_n393), .A3(new_n794), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n792), .B1(new_n351), .B2(new_n795), .C1(new_n216), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n784), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n347), .B1(new_n579), .B2(new_n787), .C1(new_n777), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n780), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n800), .B(new_n802), .C1(G329), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n795), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G322), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n796), .A2(G311), .ZN(new_n807));
  INV_X1    g0607(.A(new_n772), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G326), .A2(new_n770), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n806), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n766), .B1(new_n812), .B2(new_n756), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n743), .B1(new_n748), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n743), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n677), .A2(new_n679), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n677), .A2(new_n679), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(G396));
  NOR2_X1   g0620(.A1(new_n670), .A2(new_n422), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n670), .A2(new_n409), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n419), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n422), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n712), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n821), .B1(new_n823), .B2(new_n422), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n827), .A2(new_n647), .A3(new_n683), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n815), .B1(new_n829), .B2(new_n737), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n737), .B2(new_n829), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n785), .A2(G68), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n347), .B1(new_n788), .B2(G50), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n351), .C2(new_n777), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G137), .A2(new_n770), .B1(new_n808), .B2(G150), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n797), .B2(new_n781), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G143), .B2(new_n805), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n834), .B(new_n838), .C1(G132), .C2(new_n803), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n770), .A2(G303), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n271), .B(new_n778), .C1(G107), .C2(new_n788), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n785), .A2(G87), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n803), .A2(G311), .ZN(new_n843));
  AND4_X1   g0643(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n772), .B(KEYINPUT99), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(KEYINPUT100), .B(G283), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n846), .A2(new_n848), .B1(G116), .B2(new_n796), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n844), .B1(new_n801), .B2(new_n795), .C1(new_n849), .C2(KEYINPUT101), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(KEYINPUT101), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n756), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n756), .A2(new_n744), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n743), .B1(new_n853), .B2(new_n216), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n854), .C1(new_n745), .C2(new_n827), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n831), .A2(new_n855), .ZN(G384));
  OAI211_X1 g0656(.A(new_n424), .B(new_n713), .C1(new_n706), .C2(new_n708), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n626), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT106), .Z(new_n859));
  NAND2_X1  g0659(.A1(new_n350), .A2(new_n365), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT16), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n375), .B1(new_n862), .B2(new_n369), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n665), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n402), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n665), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n377), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n388), .A2(new_n867), .A3(new_n868), .A4(new_n399), .ZN(new_n869));
  AND4_X1   g0669(.A1(new_n367), .A2(new_n397), .A3(new_n371), .A4(new_n376), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n863), .B1(new_n386), .B2(new_n665), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT103), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(new_n864), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n615), .B2(new_n620), .ZN(new_n878));
  INV_X1    g0678(.A(new_n873), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n865), .A2(new_n881), .A3(KEYINPUT38), .A4(new_n873), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n821), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n828), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n338), .B(new_n342), .C1(new_n340), .C2(new_n683), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n337), .B(new_n670), .C1(new_n322), .C2(new_n616), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n665), .B1(new_n613), .B2(new_n614), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n322), .A2(new_n683), .A3(new_n337), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n880), .A2(new_n882), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n402), .A2(new_n864), .B1(new_n869), .B2(new_n872), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n881), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT39), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n402), .A2(new_n377), .A3(new_n866), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n388), .A2(new_n867), .A3(new_n399), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT104), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(new_n869), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n897), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n876), .ZN(new_n904));
  XOR2_X1   g0704(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n874), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n892), .B1(new_n896), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n891), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n859), .B(new_n908), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n888), .A2(new_n827), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n730), .A2(new_n731), .ZN(new_n911));
  OAI211_X1 g0711(.A(KEYINPUT31), .B(new_n670), .C1(new_n911), .C2(new_n727), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n715), .A2(new_n912), .A3(new_n733), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n904), .A2(new_n874), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n914), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n917), .A2(KEYINPUT40), .B1(new_n918), .B2(new_n883), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n424), .A2(new_n913), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n678), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n909), .A2(new_n922), .B1(new_n205), .B2(new_n741), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n909), .B2(new_n922), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n530), .A2(new_n531), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT102), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT35), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(G116), .A3(new_n749), .A4(new_n361), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(KEYINPUT35), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n226), .A2(new_n216), .A3(new_n352), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n266), .A2(G68), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n205), .B(G13), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n924), .A2(new_n931), .A3(new_n934), .ZN(G367));
  NAND2_X1  g0735(.A1(new_n761), .A2(new_n243), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n232), .B2(new_n405), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n815), .B1(new_n937), .B2(new_n758), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n784), .A2(new_n216), .ZN(new_n939));
  XNOR2_X1  g0739(.A(KEYINPUT111), .B(G137), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n271), .B1(new_n351), .B2(new_n787), .C1(new_n780), .C2(new_n940), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(new_n846), .C2(G159), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n266), .B2(new_n797), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n770), .A2(G143), .B1(G68), .B2(new_n776), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n254), .B2(new_n795), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(KEYINPUT110), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(KEYINPUT110), .B2(new_n945), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n846), .A2(G294), .B1(new_n796), .B2(new_n848), .ZN(new_n948));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n543), .A2(new_n784), .B1(new_n780), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n271), .B1(new_n776), .B2(G107), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n787), .B2(new_n428), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n950), .B(new_n955), .C1(G311), .C2(new_n770), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n948), .B(new_n956), .C1(new_n579), .C2(new_n795), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n947), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT47), .ZN(new_n959));
  INV_X1    g0759(.A(new_n756), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n958), .B2(KEYINPUT47), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n938), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n628), .B(new_n683), .C1(new_n475), .C2(new_n478), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n475), .A2(new_n478), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n629), .B1(new_n670), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n962), .B1(new_n747), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT112), .Z(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n571), .B1(new_n667), .B2(new_n669), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n683), .A2(new_n566), .B1(new_n972), .B2(new_n574), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n686), .A2(KEYINPUT42), .A3(new_n688), .A4(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n973), .A2(new_n688), .A3(new_n685), .A4(new_n682), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT42), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n572), .A2(new_n573), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n566), .B1(new_n979), .B2(new_n526), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n683), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n967), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n974), .A2(new_n977), .B1(new_n683), .B2(new_n980), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n966), .B1(new_n985), .B2(KEYINPUT107), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n984), .A2(new_n986), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n971), .B(new_n988), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n990), .B1(new_n984), .B2(new_n986), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT108), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n687), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n973), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n991), .A2(new_n994), .A3(new_n996), .A4(new_n973), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n742), .A2(G1), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n709), .A2(new_n713), .B1(new_n679), .B2(new_n736), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n689), .A2(new_n1004), .A3(new_n973), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n689), .B2(new_n973), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n689), .A2(new_n973), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1003), .B(new_n996), .C1(new_n1007), .C2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1006), .A2(new_n1005), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT109), .B1(new_n1014), .B2(new_n687), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n687), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n686), .B(new_n688), .Z(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(new_n817), .Z(new_n1019));
  OAI21_X1  g0819(.A(new_n1002), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n692), .B(KEYINPUT41), .Z(new_n1021));
  AOI21_X1  g0821(.A(new_n1001), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n970), .B1(new_n1000), .B2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n738), .A2(new_n1019), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1019), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1002), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n692), .B(KEYINPUT116), .Z(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n796), .A2(G68), .B1(new_n372), .B2(new_n808), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT113), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n271), .B1(new_n216), .B2(new_n787), .C1(new_n784), .C2(new_n543), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n457), .A2(new_n459), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1032), .A2(new_n777), .B1(new_n254), .B2(new_n780), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(G159), .C2(new_n770), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1030), .B(new_n1034), .C1(new_n266), .C2(new_n795), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n796), .A2(G303), .B1(new_n770), .B2(G322), .ZN(new_n1036));
  INV_X1    g0836(.A(G311), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1036), .B1(new_n949), .B2(new_n795), .C1(new_n845), .C2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1038), .A2(KEYINPUT114), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(KEYINPUT114), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT48), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT48), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n788), .B1(new_n776), .B2(new_n848), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(KEYINPUT115), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n271), .B1(new_n803), .B2(G326), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n428), .C2(new_n784), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT115), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1035), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n756), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n764), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1054), .A2(new_n693), .B1(G107), .B2(new_n232), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n761), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n693), .B(new_n434), .C1(new_n210), .C2(new_n216), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n258), .B2(G50), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n372), .A2(KEYINPUT50), .A3(new_n266), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n240), .A2(G45), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n815), .B1(new_n1064), .B2(new_n758), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n686), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n746), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1053), .A2(new_n1067), .B1(new_n1001), .B2(new_n1025), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1028), .A2(new_n1068), .ZN(G393));
  XNOR2_X1  g0869(.A(new_n1014), .B(new_n996), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1070), .A2(new_n1001), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n973), .A2(new_n747), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n771), .A2(new_n949), .B1(new_n795), .B2(new_n1037), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n803), .A2(G322), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n776), .A2(G116), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n271), .B1(new_n788), .B2(new_n848), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n786), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n797), .A2(new_n801), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n846), .C2(G303), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n803), .A2(G143), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n776), .A2(G77), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n347), .B1(new_n788), .B2(G68), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n842), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n797), .A2(new_n258), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n846), .C2(G50), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n771), .A2(new_n254), .B1(new_n795), .B2(new_n781), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1074), .A2(new_n1080), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(new_n960), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n761), .A2(new_n251), .B1(G97), .B2(new_n763), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n743), .B1(new_n1091), .B2(new_n757), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1072), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1071), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1027), .B1(new_n1026), .B2(new_n1017), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1070), .B1(new_n1002), .B2(new_n1025), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(G390));
  AOI21_X1  g0897(.A(new_n825), .B1(new_n702), .B2(new_n704), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n888), .B1(new_n1098), .B2(new_n821), .ZN(new_n1099));
  AOI221_X4 g0899(.A(new_n876), .B1(new_n869), .B2(new_n872), .C1(new_n402), .C2(new_n864), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n876), .B2(new_n903), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n892), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n646), .A2(new_n628), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n670), .B1(new_n1105), .B2(new_n634), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n821), .B1(new_n1106), .B2(new_n827), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n886), .A2(new_n887), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n892), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n896), .A3(new_n906), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n888), .A2(new_n736), .A3(new_n679), .A4(new_n827), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1104), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n888), .A2(new_n913), .A3(G330), .A4(new_n827), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1001), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(KEYINPUT39), .A2(new_n883), .B1(new_n1101), .B2(new_n905), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n744), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n853), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n815), .B1(new_n1119), .B2(new_n372), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n788), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n787), .B2(new_n254), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n271), .B1(new_n784), .B2(new_n266), .C1(new_n777), .C2(new_n781), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(G125), .C2(new_n803), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n771), .C1(new_n797), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G132), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n845), .A2(new_n940), .B1(new_n1130), .B2(new_n795), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n271), .B1(new_n788), .B2(G87), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n832), .A2(new_n1082), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G294), .B2(new_n803), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n799), .B2(new_n771), .C1(new_n543), .C2(new_n797), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n845), .A2(new_n218), .B1(new_n428), .B2(new_n795), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1129), .A2(new_n1131), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1120), .B1(new_n1137), .B2(new_n756), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1118), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1116), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n705), .A2(new_n824), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n913), .A2(G330), .A3(new_n827), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1108), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1141), .A2(new_n884), .A3(new_n1111), .A4(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n736), .A2(new_n679), .A3(new_n827), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1108), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1113), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n885), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n424), .A2(G330), .A3(new_n913), .ZN(new_n1150));
  AND4_X1   g0950(.A1(new_n626), .A2(new_n1149), .A3(new_n857), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT117), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1104), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1114), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1117), .A2(new_n1109), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1153), .B1(new_n1156), .B2(new_n1113), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1149), .A2(new_n857), .A3(new_n626), .A4(new_n1150), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT117), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1027), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1140), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G378));
  OAI21_X1  g0964(.A(KEYINPUT121), .B1(new_n908), .B2(KEYINPUT120), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT120), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n891), .C2(new_n907), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n866), .A2(new_n269), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n304), .B(new_n1170), .Z(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n919), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1172), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1171), .B(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n918), .A2(new_n883), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT40), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n915), .B2(new_n916), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(G330), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1175), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1169), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1165), .A2(new_n1168), .A3(new_n1175), .A4(new_n1181), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1001), .A3(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n777), .A2(new_n254), .B1(new_n787), .B2(new_n1128), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n772), .A2(new_n1130), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G125), .C2(new_n770), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n796), .A2(G137), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1127), .C2(new_n795), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n255), .B(new_n691), .C1(new_n784), .C2(new_n781), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G124), .B2(new_n803), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n770), .A2(G116), .B1(G68), .B2(new_n776), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT118), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n218), .B2(new_n795), .C1(new_n1032), .C2(new_n797), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1196), .A2(KEYINPUT118), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n347), .A2(new_n691), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n784), .A2(new_n351), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G77), .C2(new_n788), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n543), .B2(new_n772), .C1(new_n799), .C2(new_n780), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1198), .A2(new_n1199), .A3(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT58), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT58), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1200), .B(new_n266), .C1(G33), .C2(G41), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1195), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n815), .B1(G50), .B2(new_n1119), .C1(new_n1208), .C2(new_n960), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1173), .B2(new_n744), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT119), .Z(new_n1211));
  AND2_X1   g1011(.A1(new_n1185), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n857), .A2(new_n626), .A3(new_n1150), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1152), .B1(new_n1115), .B2(new_n1151), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1157), .A2(KEYINPUT117), .A3(new_n1158), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AND4_X1   g1017(.A1(new_n1165), .A2(new_n1168), .A3(new_n1175), .A4(new_n1181), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1165), .A2(new_n1168), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1175), .A2(new_n1181), .A3(new_n908), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n908), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1027), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1212), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT122), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(G375));
  INV_X1    g1031(.A(new_n1149), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1213), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1021), .B(KEYINPUT123), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1158), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1108), .A2(new_n744), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n815), .B1(new_n1119), .B2(G68), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n846), .A2(G116), .B1(G107), .B2(new_n796), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n799), .B2(new_n795), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n939), .A2(new_n271), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT124), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1032), .A2(new_n777), .B1(new_n543), .B2(new_n787), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G303), .B2(new_n803), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(new_n801), .C2(new_n771), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n271), .B1(new_n781), .B2(new_n787), .C1(new_n777), .C2(new_n266), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1201), .B(new_n1245), .C1(G128), .C2(new_n803), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n1130), .B2(new_n771), .C1(new_n795), .C2(new_n940), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n845), .A2(new_n1128), .B1(new_n797), .B2(new_n254), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1239), .A2(new_n1244), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1237), .B1(new_n1249), .B2(new_n756), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1149), .A2(new_n1001), .B1(new_n1236), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1235), .A2(new_n1251), .ZN(G381));
  INV_X1    g1052(.A(G396), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1028), .A2(new_n1253), .A3(new_n1068), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G384), .A2(G390), .A3(new_n1254), .A4(G381), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(G387), .A3(G378), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1229), .B2(new_n1230), .ZN(G407));
  OAI21_X1  g1057(.A(new_n1163), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G407), .B(G213), .C1(new_n1258), .C2(G343), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1259), .B(new_n1260), .ZN(G409));
  OAI211_X1 g1061(.A(G378), .B(new_n1212), .C1(new_n1221), .C2(new_n1226), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1234), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1222), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1001), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1211), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1163), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n666), .A2(G213), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1233), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1213), .A2(KEYINPUT60), .A3(new_n1232), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1027), .A3(new_n1158), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1251), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n831), .A3(new_n855), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(G384), .A3(new_n1251), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1270), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G2897), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1279), .B(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1262), .B2(new_n1268), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1284), .A2(KEYINPUT62), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT62), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1283), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1254), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G390), .B(new_n970), .C1(new_n1000), .C2(new_n1022), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n999), .B(new_n998), .C1(new_n1293), .C2(new_n1001), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G390), .B1(new_n1294), .B2(new_n970), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1290), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G390), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1290), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1291), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1288), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1279), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1269), .A2(new_n1270), .A3(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1304), .B1(new_n1311), .B2(new_n1283), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1269), .A2(new_n1270), .A3(new_n1285), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1305), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1301), .B1(new_n1284), .B2(new_n1306), .ZN(new_n1315));
  AND4_X1   g1115(.A1(new_n1304), .A2(new_n1283), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1303), .B1(new_n1312), .B2(new_n1316), .ZN(G405));
  INV_X1    g1117(.A(new_n1227), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1258), .B1(new_n1163), .B2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1301), .B(new_n1279), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1319), .B(new_n1320), .ZN(G402));
endmodule


