

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U319 ( .A(n352), .B(n287), .ZN(n353) );
  XNOR2_X1 U320 ( .A(n366), .B(n365), .ZN(n562) );
  AND2_X1 U321 ( .A1(G227GAT), .A2(G233GAT), .ZN(n287) );
  XNOR2_X1 U322 ( .A(n450), .B(n449), .ZN(n452) );
  NOR2_X1 U323 ( .A1(n383), .A2(n382), .ZN(n406) );
  XOR2_X1 U324 ( .A(G120GAT), .B(G71GAT), .Z(n425) );
  XNOR2_X1 U325 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U326 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U327 ( .A(n364), .B(KEYINPUT99), .ZN(n365) );
  XNOR2_X1 U328 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U329 ( .A(n363), .B(n390), .Z(n471) );
  NOR2_X1 U330 ( .A1(n471), .A2(n470), .ZN(n556) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(n495) );
  XNOR2_X1 U332 ( .A(n472), .B(G176GAT), .ZN(n473) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n447) );
  XNOR2_X1 U334 ( .A(n474), .B(n473), .ZN(G1349GAT) );
  XNOR2_X1 U335 ( .A(n448), .B(n447), .ZN(G1330GAT) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U337 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n288) );
  XNOR2_X1 U338 ( .A(n288), .B(KEYINPUT71), .ZN(n416) );
  XOR2_X1 U339 ( .A(n434), .B(n416), .Z(n290) );
  NAND2_X1 U340 ( .A1(G231GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U341 ( .A(n290), .B(n289), .ZN(n306) );
  XOR2_X1 U342 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n292) );
  XNOR2_X1 U343 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n304) );
  XOR2_X1 U345 ( .A(G155GAT), .B(G78GAT), .Z(n294) );
  XNOR2_X1 U346 ( .A(G22GAT), .B(G211GAT), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n296) );
  XNOR2_X1 U349 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U351 ( .A(G64GAT), .B(G71GAT), .Z(n298) );
  XNOR2_X1 U352 ( .A(G127GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n300), .B(n299), .Z(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n304), .B(n303), .Z(n305) );
  XOR2_X1 U357 ( .A(n306), .B(n305), .Z(n475) );
  INV_X1 U358 ( .A(KEYINPUT77), .ZN(n325) );
  XOR2_X1 U359 ( .A(G43GAT), .B(G29GAT), .Z(n308) );
  XNOR2_X1 U360 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(n309), .B(KEYINPUT8), .Z(n311) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(KEYINPUT69), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n444) );
  XOR2_X1 U365 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n313) );
  XNOR2_X1 U366 ( .A(KEYINPUT65), .B(KEYINPUT75), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n444), .B(n314), .ZN(n324) );
  XOR2_X1 U369 ( .A(G85GAT), .B(G92GAT), .Z(n316) );
  XNOR2_X1 U370 ( .A(G99GAT), .B(G106GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n418) );
  XOR2_X1 U372 ( .A(G218GAT), .B(G162GAT), .Z(n327) );
  XOR2_X1 U373 ( .A(n418), .B(n327), .Z(n318) );
  NAND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U376 ( .A(G190GAT), .B(G134GAT), .Z(n347) );
  XNOR2_X1 U377 ( .A(n347), .B(KEYINPUT11), .ZN(n320) );
  INV_X1 U378 ( .A(KEYINPUT10), .ZN(n319) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n550) );
  XNOR2_X1 U380 ( .A(n325), .B(n550), .ZN(n557) );
  XNOR2_X1 U381 ( .A(KEYINPUT36), .B(n557), .ZN(n576) );
  AND2_X1 U382 ( .A1(n475), .A2(n576), .ZN(n414) );
  INV_X1 U383 ( .A(KEYINPUT101), .ZN(n408) );
  XNOR2_X1 U384 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n326), .B(KEYINPUT3), .ZN(n391) );
  XOR2_X1 U386 ( .A(n391), .B(n327), .Z(n333) );
  XOR2_X1 U387 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XNOR2_X1 U388 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n328), .B(G148GAT), .ZN(n419) );
  XOR2_X1 U390 ( .A(n419), .B(KEYINPUT24), .Z(n330) );
  NAND2_X1 U391 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n432), .B(n331), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U395 ( .A(KEYINPUT91), .B(G204GAT), .Z(n335) );
  XNOR2_X1 U396 ( .A(G50GAT), .B(G106GAT), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(n337), .B(n336), .Z(n346) );
  XNOR2_X1 U399 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n338), .B(KEYINPUT90), .ZN(n339) );
  XOR2_X1 U401 ( .A(n339), .B(KEYINPUT21), .Z(n341) );
  XNOR2_X1 U402 ( .A(G197GAT), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n379) );
  XOR2_X1 U404 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT92), .B(KEYINPUT87), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n379), .B(n344), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n467) );
  XOR2_X1 U409 ( .A(G99GAT), .B(n425), .Z(n349) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(n347), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U412 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n351) );
  XNOR2_X1 U413 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(G183GAT), .B(KEYINPUT19), .Z(n356) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n372) );
  XOR2_X1 U418 ( .A(n357), .B(n372), .Z(n359) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G15GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n361) );
  XNOR2_X1 U422 ( .A(KEYINPUT84), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(G113GAT), .B(n362), .Z(n390) );
  INV_X1 U425 ( .A(n471), .ZN(n527) );
  NOR2_X1 U426 ( .A1(n467), .A2(n527), .ZN(n366) );
  XNOR2_X1 U427 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n364) );
  XOR2_X1 U428 ( .A(G92GAT), .B(KEYINPUT97), .Z(n368) );
  NAND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n371) );
  XOR2_X1 U431 ( .A(KEYINPUT73), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U432 ( .A(G176GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n417) );
  XOR2_X1 U434 ( .A(n371), .B(n417), .Z(n374) );
  XNOR2_X1 U435 ( .A(n372), .B(G190GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n375), .B(G218GAT), .Z(n377) );
  XOR2_X1 U438 ( .A(G169GAT), .B(G8GAT), .Z(n439) );
  XNOR2_X1 U439 ( .A(G36GAT), .B(n439), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n515) );
  XOR2_X1 U442 ( .A(KEYINPUT27), .B(n515), .Z(n409) );
  NOR2_X1 U443 ( .A1(n562), .A2(n409), .ZN(n383) );
  NAND2_X1 U444 ( .A1(n527), .A2(n515), .ZN(n380) );
  NAND2_X1 U445 ( .A1(n467), .A2(n380), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n381), .B(KEYINPUT25), .ZN(n382) );
  XOR2_X1 U447 ( .A(KEYINPUT96), .B(KEYINPUT93), .Z(n385) );
  XNOR2_X1 U448 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U450 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n387) );
  XNOR2_X1 U451 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U453 ( .A(n389), .B(n388), .Z(n397) );
  INV_X1 U454 ( .A(n390), .ZN(n395) );
  XOR2_X1 U455 ( .A(n391), .B(KEYINPUT6), .Z(n393) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n395), .B(n394), .Z(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n405) );
  XOR2_X1 U460 ( .A(G148GAT), .B(G120GAT), .Z(n399) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(G1GAT), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G162GAT), .Z(n401) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G134GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U466 ( .A(n403), .B(n402), .Z(n404) );
  XOR2_X1 U467 ( .A(n405), .B(n404), .Z(n560) );
  INV_X1 U468 ( .A(n560), .ZN(n513) );
  NOR2_X1 U469 ( .A1(n406), .A2(n513), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n413) );
  NOR2_X1 U471 ( .A1(n560), .A2(n409), .ZN(n525) );
  XOR2_X1 U472 ( .A(n467), .B(KEYINPUT28), .Z(n520) );
  INV_X1 U473 ( .A(n520), .ZN(n526) );
  NAND2_X1 U474 ( .A1(n525), .A2(n526), .ZN(n410) );
  NOR2_X1 U475 ( .A1(n527), .A2(n410), .ZN(n411) );
  XNOR2_X1 U476 ( .A(KEYINPUT98), .B(n411), .ZN(n412) );
  OR2_X1 U477 ( .A1(n413), .A2(n412), .ZN(n478) );
  NAND2_X1 U478 ( .A1(n414), .A2(n478), .ZN(n415) );
  XOR2_X1 U479 ( .A(KEYINPUT37), .B(n415), .Z(n512) );
  XOR2_X1 U480 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U483 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n423) );
  XNOR2_X1 U484 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U486 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n570) );
  INV_X1 U490 ( .A(n570), .ZN(n451) );
  XOR2_X1 U491 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n431) );
  XNOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U495 ( .A(n434), .B(KEYINPUT67), .Z(n436) );
  NAND2_X1 U496 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n442) );
  XNOR2_X1 U500 ( .A(G197GAT), .B(G113GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n500) );
  XOR2_X1 U503 ( .A(KEYINPUT70), .B(n500), .Z(n552) );
  NAND2_X1 U504 ( .A1(n451), .A2(n552), .ZN(n480) );
  NOR2_X1 U505 ( .A1(n512), .A2(n480), .ZN(n446) );
  XOR2_X1 U506 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n445) );
  NAND2_X1 U507 ( .A1(n495), .A2(n527), .ZN(n448) );
  XOR2_X1 U508 ( .A(KEYINPUT54), .B(KEYINPUT123), .Z(n466) );
  INV_X1 U509 ( .A(n475), .ZN(n574) );
  NAND2_X1 U510 ( .A1(n574), .A2(n576), .ZN(n450) );
  XOR2_X1 U511 ( .A(KEYINPUT45), .B(KEYINPUT116), .Z(n449) );
  NAND2_X1 U512 ( .A1(n452), .A2(n451), .ZN(n453) );
  NOR2_X1 U513 ( .A1(n552), .A2(n453), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n454), .B(KEYINPUT117), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n456) );
  INV_X1 U516 ( .A(n500), .ZN(n566) );
  XOR2_X1 U517 ( .A(n570), .B(KEYINPUT41), .Z(n544) );
  NAND2_X1 U518 ( .A1(n566), .A2(n544), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n574), .A2(n457), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n458), .B(KEYINPUT115), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n550), .A2(n459), .ZN(n460) );
  XNOR2_X1 U523 ( .A(KEYINPUT47), .B(n460), .ZN(n461) );
  NAND2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n464) );
  XNOR2_X1 U525 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(n524) );
  NAND2_X1 U527 ( .A1(n515), .A2(n524), .ZN(n465) );
  XOR2_X1 U528 ( .A(n466), .B(n465), .Z(n561) );
  AND2_X1 U529 ( .A1(n467), .A2(n560), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n561), .A2(n468), .ZN(n469) );
  XOR2_X1 U531 ( .A(KEYINPUT55), .B(n469), .Z(n470) );
  NAND2_X1 U532 ( .A1(n556), .A2(n544), .ZN(n474) );
  XOR2_X1 U533 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n472) );
  NOR2_X1 U534 ( .A1(n557), .A2(n475), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n501) );
  NOR2_X1 U538 ( .A1(n480), .A2(n501), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT102), .B(n481), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n488), .A2(n513), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n488), .A2(n515), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U546 ( .A1(n488), .A2(n527), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U548 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  NAND2_X1 U549 ( .A1(n488), .A2(n520), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n495), .A2(n513), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n491) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n515), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(G50GAT), .B(KEYINPUT107), .Z(n497) );
  NAND2_X1 U559 ( .A1(n520), .A2(n495), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT109), .ZN(n499) );
  XOR2_X1 U563 ( .A(KEYINPUT108), .B(n499), .Z(n503) );
  NAND2_X1 U564 ( .A1(n500), .A2(n544), .ZN(n511) );
  NOR2_X1 U565 ( .A1(n501), .A2(n511), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n507), .A2(n513), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n515), .A2(n507), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(KEYINPUT110), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n527), .A2(n507), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U574 ( .A1(n507), .A2(n520), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n510), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n513), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n521), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT112), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT113), .Z(n519) );
  NAND2_X1 U584 ( .A1(n521), .A2(n527), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(KEYINPUT118), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n539), .A2(n528), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n536), .A2(n552), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n536), .A2(n544), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n574), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n557), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n562), .A2(n539), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n566), .A2(n549), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n542) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(n543), .Z(n546) );
  NAND2_X1 U612 ( .A1(n549), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n574), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT122), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n556), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT124), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n574), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n559), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  AND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n564) );
  INV_X1 U629 ( .A(n562), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT125), .B(n565), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

