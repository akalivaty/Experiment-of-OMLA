//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0011(.A1(new_n206), .A2(new_n207), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(G20), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n216), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n215), .B(new_n219), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT67), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n207), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT70), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(new_n213), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n258), .B2(new_n213), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  INV_X1    g0064(.A(G20), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n264), .A2(new_n265), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n257), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n253), .A2(new_n266), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n258), .A2(new_n213), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n260), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT7), .B1(new_n278), .B2(new_n265), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT7), .ZN(new_n280));
  AOI211_X1 g0080(.A(new_n280), .B(G20), .C1(new_n275), .C2(new_n277), .ZN(new_n281));
  OAI21_X1  g0081(.A(G68), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G58), .A2(G68), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n204), .A2(new_n205), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n284), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT16), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n273), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(KEYINPUT16), .A3(new_n286), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n270), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G232), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G1), .A3(G13), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(G274), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n295), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G179), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n275), .A2(new_n277), .A3(G223), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G87), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n292), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n292), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n303), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n296), .A2(G232), .B1(new_n300), .B2(new_n295), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n309), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT18), .B1(new_n291), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT3), .B(G33), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n280), .B1(new_n320), .B2(G20), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n265), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n203), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n284), .A2(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n285), .A2(G159), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n288), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n290), .A2(new_n327), .A3(new_n263), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n257), .A2(new_n267), .B1(new_n266), .B2(new_n253), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n292), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT74), .B1(new_n308), .B2(new_n292), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(new_n303), .B1(new_n316), .B2(new_n315), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT17), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n302), .A2(G190), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n333), .A2(new_n338), .B1(new_n339), .B2(new_n315), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n311), .A2(new_n342), .A3(new_n312), .A4(new_n314), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n315), .A2(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n345), .A2(KEYINPUT17), .A3(new_n328), .A4(new_n329), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n319), .A2(new_n336), .A3(new_n341), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n266), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n273), .A2(G77), .A3(new_n348), .A4(new_n255), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT71), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n250), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n265), .A2(G33), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G77), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n356), .A2(new_n263), .B1(new_n357), .B2(new_n266), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n320), .A2(G232), .A3(new_n305), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n320), .A2(G238), .A3(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G107), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n320), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n292), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n296), .A2(G244), .B1(new_n300), .B2(new_n295), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n316), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(new_n368), .A3(new_n365), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n359), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(G200), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(G190), .A3(new_n365), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n371), .A2(new_n351), .A3(new_n358), .A4(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n370), .A2(KEYINPUT72), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT72), .B1(new_n370), .B2(new_n373), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n347), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n267), .A2(G68), .A3(new_n255), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n357), .B2(new_n354), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n263), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n266), .A2(new_n203), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT12), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n263), .A2(new_n379), .A3(KEYINPUT11), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n377), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT14), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n275), .A2(new_n277), .A3(G232), .A4(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(new_n305), .ZN(new_n389));
  INV_X1    g0189(.A(G97), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n388), .B(new_n389), .C1(new_n274), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n292), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n296), .A2(G238), .B1(new_n300), .B2(new_n295), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n387), .B(G169), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n393), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(G179), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n387), .B1(new_n403), .B2(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n386), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n386), .ZN(new_n406));
  OAI21_X1  g0206(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(G190), .A3(new_n400), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n376), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n320), .A2(G222), .A3(new_n305), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n278), .A2(G77), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n275), .A2(new_n277), .A3(G223), .A4(G1698), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n292), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT68), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n296), .A2(G226), .B1(new_n300), .B2(new_n295), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n416), .B2(new_n418), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n316), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n208), .A2(G20), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n285), .A2(G150), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(new_n253), .C2(new_n354), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n263), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n256), .A2(new_n207), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n267), .A2(new_n427), .B1(new_n207), .B2(new_n266), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n368), .B1(new_n419), .B2(new_n420), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G190), .B1(new_n419), .B2(new_n420), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT73), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT73), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(G190), .C1(new_n419), .C2(new_n420), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(KEYINPUT9), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT9), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n426), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n437), .A2(new_n439), .B1(new_n421), .B2(G200), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT10), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n436), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n436), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n431), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n411), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(new_n305), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT4), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n320), .A2(KEYINPUT4), .A3(G244), .A4(new_n305), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n320), .A2(G250), .A3(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n292), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT77), .B1(new_n454), .B2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n293), .A3(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n254), .A2(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n292), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n254), .B(G45), .C1(new_n293), .C2(KEYINPUT5), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n455), .B2(new_n457), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n462), .A2(G257), .B1(new_n464), .B2(new_n300), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n453), .A2(G179), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n453), .A2(new_n465), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n316), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n348), .A2(G97), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n279), .B2(new_n281), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n285), .A2(G77), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT6), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n474), .A2(G97), .A3(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n390), .A2(KEYINPUT6), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT75), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n475), .A2(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n390), .A2(new_n362), .A3(KEYINPUT6), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(G107), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(G20), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n472), .A2(new_n473), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n471), .B1(new_n487), .B2(new_n263), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n254), .A2(G33), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n348), .B(new_n489), .C1(new_n261), .C2(new_n262), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT76), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n273), .A2(KEYINPUT76), .A3(new_n348), .A4(new_n489), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(G97), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n470), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n486), .A2(new_n473), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n362), .B1(new_n321), .B2(new_n322), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n263), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n471), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n470), .A2(new_n498), .A3(new_n494), .A4(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n469), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n494), .A3(new_n499), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n453), .A2(G190), .A3(new_n465), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n339), .B1(new_n453), .B2(new_n465), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n355), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n492), .A2(new_n493), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n320), .A2(new_n265), .A3(G68), .ZN(new_n509));
  NAND3_X1  g0309(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n265), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n390), .A3(new_n362), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n265), .A2(G33), .A3(G97), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(KEYINPUT79), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT79), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n509), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n263), .B1(new_n266), .B2(new_n355), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n508), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n299), .A2(new_n254), .A3(G45), .A4(G274), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n299), .A2(G250), .A3(new_n460), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n275), .A2(new_n277), .A3(G238), .A4(new_n305), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n292), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n368), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G169), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(G190), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n339), .B2(new_n529), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n492), .A2(new_n493), .A3(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n520), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n501), .A2(new_n506), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n254), .A2(new_n540), .A3(G13), .A4(G20), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n541), .A2(KEYINPUT80), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(KEYINPUT80), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n258), .A2(new_n213), .B1(G20), .B2(new_n540), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n451), .B(new_n265), .C1(G33), .C2(new_n390), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT20), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n490), .A2(new_n540), .ZN(new_n551));
  OAI21_X1  g0351(.A(G179), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n276), .A2(G33), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n554));
  OAI21_X1  g0354(.A(G303), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n275), .A2(new_n277), .A3(G264), .A4(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(new_n305), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n292), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n462), .A2(G270), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n464), .A2(new_n300), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n540), .A2(G20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n546), .A2(new_n271), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n547), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n273), .A2(G116), .A3(new_n348), .A4(new_n489), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n544), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n562), .A3(G169), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT21), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n567), .A2(new_n547), .B1(new_n543), .B2(new_n542), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n316), .B1(new_n573), .B2(new_n569), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n562), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n563), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n462), .A2(G264), .B1(new_n464), .B2(new_n300), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(new_n305), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G294), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n292), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n368), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n458), .A2(new_n461), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(G264), .A3(new_n299), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n561), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n316), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n275), .A2(new_n277), .A3(new_n265), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n320), .A2(new_n591), .A3(new_n265), .A4(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n527), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n265), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n362), .A2(KEYINPUT23), .A3(G20), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT24), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n593), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n273), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n492), .A2(new_n493), .A3(G107), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n266), .A2(new_n362), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT25), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n584), .B(new_n588), .C1(new_n603), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n587), .A2(new_n339), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(G190), .B2(new_n587), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n600), .A2(new_n602), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n263), .ZN(new_n613));
  INV_X1    g0413(.A(new_n608), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n562), .A2(G200), .ZN(new_n616));
  INV_X1    g0416(.A(new_n570), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n342), .C2(new_n562), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n577), .A2(new_n609), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n539), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n445), .A2(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n532), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n552), .A2(new_n562), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n571), .A2(KEYINPUT21), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n575), .B1(new_n574), .B2(new_n562), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n588), .A2(new_n584), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n613), .B2(new_n614), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n615), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n622), .B1(new_n539), .B2(new_n629), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n521), .A2(new_n531), .B1(new_n534), .B2(new_n536), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT26), .B1(new_n501), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n453), .A2(G179), .A3(new_n465), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n316), .B1(new_n453), .B2(new_n465), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n502), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n631), .A2(new_n635), .A3(KEYINPUT26), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n445), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT81), .Z(new_n640));
  INV_X1    g0440(.A(new_n431), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n442), .A2(new_n443), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n319), .A2(new_n336), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n341), .A2(new_n410), .A3(new_n346), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n359), .A2(new_n367), .A3(new_n369), .ZN(new_n645));
  OAI21_X1  g0445(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n401), .A3(new_n397), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(new_n386), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n643), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n641), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n640), .A2(new_n651), .ZN(G369));
  NAND3_X1  g0452(.A1(new_n254), .A2(new_n265), .A3(G13), .ZN(new_n653));
  OAI21_X1  g0453(.A(G213), .B1(new_n653), .B2(KEYINPUT27), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(KEYINPUT27), .B2(new_n653), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT82), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT82), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n656), .A2(G343), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n617), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n626), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n623), .B(new_n618), .C1(new_n624), .C2(new_n625), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n660), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n615), .A2(new_n609), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n603), .A2(new_n608), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n659), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n609), .B2(new_n659), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n577), .A2(new_n658), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n628), .A2(new_n659), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(G399));
  NOR2_X1   g0477(.A1(new_n513), .A2(G116), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT83), .Z(new_n679));
  INV_X1    g0479(.A(new_n217), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n254), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n679), .A2(new_n682), .B1(new_n212), .B2(new_n681), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  NOR2_X1   g0484(.A1(new_n633), .A2(new_n634), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n502), .A2(KEYINPUT78), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n488), .A2(new_n470), .A3(new_n494), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n688), .A2(new_n631), .A3(new_n505), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n577), .A2(new_n609), .B1(new_n668), .B2(new_n611), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n532), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n538), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n636), .B1(new_n692), .B2(KEYINPUT26), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n658), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT85), .B(KEYINPUT29), .Z(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT86), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT26), .B1(new_n631), .B2(new_n635), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n692), .B2(KEYINPUT26), .ZN(new_n698));
  OAI211_X1 g0498(.A(KEYINPUT29), .B(new_n659), .C1(new_n630), .C2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n659), .B1(new_n630), .B2(new_n638), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT86), .ZN(new_n701));
  INV_X1    g0501(.A(new_n695), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n528), .A2(new_n292), .ZN(new_n705));
  INV_X1    g0505(.A(new_n524), .ZN(new_n706));
  AOI21_X1  g0506(.A(G179), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n467), .A2(new_n587), .A3(new_n562), .A4(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT84), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n292), .A2(new_n558), .B1(new_n462), .B2(G270), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n453), .A2(new_n465), .B1(new_n711), .B2(new_n561), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n707), .A2(new_n587), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT84), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n559), .A2(new_n560), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n705), .A2(new_n706), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n587), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n633), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n711), .A2(new_n529), .A3(new_n583), .A4(new_n578), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n466), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n710), .A2(new_n714), .A3(new_n718), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n658), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n658), .A2(KEYINPUT31), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n718), .A2(new_n721), .A3(new_n708), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n723), .A2(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n666), .A2(new_n662), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n686), .A2(new_n687), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n505), .B1(new_n730), .B2(new_n469), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(new_n731), .A3(new_n538), .A4(new_n659), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n704), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n684), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n213), .B1(G20), .B2(new_n316), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n342), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n265), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n390), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n265), .A2(new_n368), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n342), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n741), .B1(G50), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n265), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(new_n342), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n278), .B1(new_n748), .B2(G107), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n742), .A2(KEYINPUT89), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(KEYINPUT89), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n745), .B(new_n749), .C1(new_n357), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n752), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT91), .B(KEYINPUT32), .Z(new_n758));
  XNOR2_X1  g0558(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n743), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n759), .B1(new_n203), .B2(new_n761), .C1(new_n512), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n342), .A2(G200), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n750), .A2(new_n751), .A3(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT90), .Z(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n754), .B(new_n763), .C1(G58), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n744), .A2(G326), .ZN(new_n769));
  INV_X1    g0569(.A(new_n755), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n320), .B1(new_n770), .B2(G329), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n769), .B(new_n771), .C1(new_n753), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n740), .ZN(new_n774));
  INV_X1    g0574(.A(new_n762), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n774), .A2(G294), .B1(new_n775), .B2(G303), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT33), .B(G317), .Z(new_n778));
  OAI221_X1 g0578(.A(new_n776), .B1(new_n777), .B2(new_n747), .C1(new_n761), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n765), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n773), .B(new_n779), .C1(G322), .C2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n738), .B1(new_n768), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n680), .A2(new_n278), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G355), .B1(new_n540), .B2(new_n680), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n245), .A2(new_n294), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n680), .A2(new_n320), .ZN(new_n786));
  INV_X1    g0586(.A(new_n212), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(G45), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT87), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n738), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n264), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n254), .B1(new_n798), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n681), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n782), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT92), .Z(new_n803));
  INV_X1    g0603(.A(new_n795), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n663), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n665), .A2(new_n801), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G330), .B2(new_n663), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n359), .A2(new_n658), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n373), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n370), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n645), .A2(new_n659), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n700), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n814), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n659), .B(new_n816), .C1(new_n630), .C2(new_n638), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n801), .B1(new_n818), .B2(new_n734), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n734), .B2(new_n818), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n738), .A2(new_n793), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n801), .B1(G77), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT93), .B(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n761), .A2(new_n823), .B1(new_n512), .B2(new_n747), .ZN(new_n824));
  INV_X1    g0624(.A(new_n744), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n826), .B1(new_n762), .B2(new_n362), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n320), .B(new_n741), .C1(G311), .C2(new_n770), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n780), .A2(G294), .ZN(new_n830));
  INV_X1    g0630(.A(new_n753), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G116), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n760), .A2(G150), .B1(new_n744), .B2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n756), .B2(new_n753), .C1(new_n766), .C2(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT94), .Z(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n775), .A2(G50), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n278), .B1(new_n770), .B2(G132), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n774), .A2(G58), .B1(new_n748), .B2(G68), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n833), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n822), .B1(new_n844), .B2(new_n738), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n794), .B2(new_n816), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n820), .A2(new_n846), .ZN(G384));
  NOR3_X1   g0647(.A1(new_n213), .A2(new_n265), .A3(new_n540), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n480), .A2(new_n485), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT35), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n212), .A2(G77), .A3(new_n283), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n241), .B(KEYINPUT95), .Z(new_n855));
  AOI211_X1 g0655(.A(new_n254), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n696), .A2(new_n445), .A3(new_n699), .A4(new_n703), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n651), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT99), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n658), .A2(new_n386), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n405), .A2(new_n410), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n386), .B(new_n658), .C1(new_n648), .C2(new_n409), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n817), .B2(new_n813), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n330), .A2(new_n334), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n656), .A2(new_n657), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n330), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n345), .A2(new_n328), .A3(new_n329), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n867), .A2(new_n869), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n347), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT96), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(KEYINPUT96), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n866), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n643), .B2(new_n868), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n648), .A2(new_n386), .A3(new_n659), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT97), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n871), .A2(new_n890), .A3(KEYINPUT37), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT98), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n874), .B(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n893), .A2(new_n895), .B1(new_n347), .B2(new_n876), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n889), .B(new_n883), .C1(new_n896), .C2(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n887), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n860), .B(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n883), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n872), .A2(KEYINPUT97), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n874), .A2(KEYINPUT98), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n867), .A2(new_n870), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n894), .A3(new_n873), .A4(new_n869), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n871), .A2(new_n890), .A3(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n902), .A2(new_n903), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n877), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n901), .B1(new_n908), .B2(new_n880), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n814), .B1(new_n862), .B2(new_n863), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT100), .B1(new_n723), .B2(new_n724), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT100), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n912), .B(KEYINPUT31), .C1(new_n722), .C2(new_n658), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n722), .A2(new_n726), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n732), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n910), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT40), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n864), .A2(new_n816), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n708), .A2(new_n709), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT84), .B1(new_n712), .B2(new_n713), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT30), .B1(new_n717), .B2(new_n633), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n720), .A2(new_n466), .A3(new_n719), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n659), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n912), .B1(new_n926), .B2(KEYINPUT31), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n723), .A2(KEYINPUT100), .A3(new_n724), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n915), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n620), .B2(new_n659), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n919), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n932), .A2(new_n884), .A3(new_n933), .A4(new_n881), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n931), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n445), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n445), .A2(new_n936), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n918), .A2(new_n938), .A3(new_n934), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(G330), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n900), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n254), .B2(new_n798), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n900), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n857), .B1(new_n942), .B2(new_n943), .ZN(G367));
  NAND3_X1  g0744(.A1(new_n532), .A2(new_n536), .A3(new_n658), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n658), .A2(new_n536), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n945), .B(KEYINPUT101), .C1(new_n631), .C2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT101), .B2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n795), .ZN(new_n949));
  INV_X1    g0749(.A(new_n796), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n680), .B2(new_n507), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n236), .A2(new_n786), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n681), .B(new_n800), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n738), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n761), .A2(new_n756), .B1(new_n825), .B2(new_n835), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n747), .A2(new_n357), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n740), .A2(new_n203), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n780), .A2(G150), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n831), .A2(G50), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT108), .B(G137), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n320), .B1(new_n755), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G58), .B2(new_n775), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(G294), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n761), .A2(new_n965), .B1(new_n362), .B2(new_n740), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G311), .B2(new_n744), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n753), .A2(new_n823), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n747), .A2(new_n390), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n278), .B1(new_n755), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n967), .B(new_n972), .C1(new_n766), .C2(new_n826), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT107), .B1(new_n762), .B2(new_n540), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n964), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  OAI211_X1 g0777(.A(new_n949), .B(new_n953), .C1(new_n954), .C2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n635), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n658), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n502), .A2(new_n658), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n501), .A2(new_n506), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT102), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n983), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n675), .C1(KEYINPUT106), .C2(KEYINPUT44), .ZN(new_n989));
  NOR2_X1   g0789(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT102), .B1(new_n731), .B2(new_n983), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n688), .A2(new_n985), .A3(new_n505), .A4(new_n982), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n980), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n990), .B1(new_n993), .B2(new_n676), .ZN(new_n994));
  NAND2_X1  g0794(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n988), .B2(new_n675), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(KEYINPUT45), .A3(new_n676), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n996), .A2(new_n671), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n671), .B1(new_n996), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n673), .B1(new_n670), .B2(new_n672), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n665), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n735), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n681), .B(KEYINPUT41), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n799), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n948), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT104), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT42), .B1(new_n988), .B2(new_n673), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n688), .B1(new_n993), .B2(new_n628), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n658), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT103), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(KEYINPUT103), .B(new_n1012), .C1(new_n1013), .C2(new_n658), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n993), .A2(new_n667), .A3(new_n672), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1011), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(KEYINPUT104), .B(new_n1020), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1010), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1017), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n501), .B1(new_n988), .B2(new_n609), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n659), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT103), .B1(new_n1027), .B2(new_n1012), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1021), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT104), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1018), .A2(new_n1011), .A3(new_n1021), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n948), .B(new_n1009), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n993), .A2(new_n665), .A3(new_n670), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1024), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1024), .B2(new_n1033), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT105), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1008), .B(new_n1035), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n978), .B1(new_n1038), .B2(new_n1039), .ZN(G387));
  OR2_X1    g0840(.A1(new_n670), .A2(new_n804), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n786), .B1(new_n233), .B2(new_n294), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n783), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n679), .B2(new_n1043), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n250), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n250), .B2(G50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n679), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1044), .A2(new_n1048), .B1(new_n362), .B2(new_n680), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n801), .B1(new_n1049), .B2(new_n950), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n774), .A2(new_n507), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n765), .B2(new_n207), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT110), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT109), .B(G150), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n278), .B(new_n969), .C1(new_n770), .C2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n744), .A2(G159), .B1(new_n775), .B2(G77), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n253), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n831), .A2(G68), .B1(new_n1057), .B2(new_n760), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT111), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n760), .A2(G311), .B1(new_n744), .B2(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n826), .B2(new_n753), .C1(new_n766), .C2(new_n970), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n740), .A2(new_n823), .B1(new_n762), .B2(new_n965), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n320), .B1(new_n770), .B2(G326), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n540), .C2(new_n747), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT49), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1060), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1050), .B1(new_n1071), .B2(new_n738), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1005), .A2(new_n800), .B1(new_n1041), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n736), .A2(new_n1005), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n681), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n736), .A2(new_n1005), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1003), .A2(new_n736), .A3(new_n1005), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n681), .A3(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n240), .A2(new_n680), .A3(new_n320), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n796), .B1(new_n390), .B2(new_n217), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n761), .A2(new_n826), .B1(new_n540), .B2(new_n740), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n780), .A2(G311), .B1(G317), .B2(new_n744), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(G294), .C2(new_n831), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n320), .B1(new_n770), .B2(G322), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n362), .B2(new_n747), .C1(new_n762), .C2(new_n823), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT112), .Z(new_n1089));
  INV_X1    g0889(.A(G150), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n756), .A2(new_n765), .B1(new_n825), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n320), .B1(new_n755), .B2(new_n835), .C1(new_n512), .C2(new_n747), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n760), .A2(G50), .B1(new_n775), .B2(G68), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n357), .B2(new_n740), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n352), .C2(new_n831), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1086), .A2(new_n1089), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n801), .B1(new_n1081), .B2(new_n1082), .C1(new_n1097), .C2(new_n954), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n988), .B2(new_n795), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1003), .B2(new_n800), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1080), .A2(new_n1100), .ZN(G390));
  NAND3_X1  g0901(.A1(new_n936), .A2(G330), .A3(new_n816), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n865), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n733), .A2(G330), .A3(new_n816), .A4(new_n864), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n659), .B(new_n812), .C1(new_n630), .C2(new_n698), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1104), .A2(new_n813), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n727), .A2(new_n726), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n926), .B2(KEYINPUT31), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n539), .A2(new_n619), .A3(new_n658), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n816), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n865), .ZN(new_n1111));
  OAI211_X1 g0911(.A(G330), .B(new_n910), .C1(new_n914), .C2(new_n916), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n817), .A2(new_n813), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1103), .A2(new_n1106), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n445), .A2(G330), .A3(new_n936), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n858), .A2(new_n651), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n887), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n888), .B(new_n897), .C1(new_n866), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1105), .A2(new_n813), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n864), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n883), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n887), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1125), .A3(new_n1104), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1112), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n888), .A2(new_n897), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n866), .A2(new_n1120), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1112), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1135), .A3(new_n681), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1130), .A2(new_n794), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n801), .B1(new_n1057), .B2(new_n821), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n761), .A2(new_n961), .B1(new_n756), .B2(new_n740), .ZN(new_n1140));
  XOR2_X1   g0940(.A(KEYINPUT54), .B(G143), .Z(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n831), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT113), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n320), .B1(new_n747), .B2(new_n207), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT114), .Z(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n825), .A2(new_n1146), .B1(new_n755), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n775), .A2(new_n1054), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(G132), .C2(new_n780), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1143), .A2(new_n1145), .A3(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n390), .A2(new_n753), .B1(new_n761), .B2(new_n362), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT115), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1153), .A2(new_n1154), .B1(new_n777), .B2(new_n825), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1154), .B2(new_n1153), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT116), .Z(new_n1157));
  OAI21_X1  g0957(.A(new_n278), .B1(new_n755), .B2(new_n965), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G87), .B2(new_n775), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n774), .A2(G77), .B1(new_n748), .B2(G68), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n540), .C2(new_n765), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1152), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1139), .B1(new_n1162), .B2(new_n738), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1137), .A2(new_n800), .B1(new_n1138), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1136), .A2(new_n1164), .ZN(G378));
  OR2_X1    g0965(.A1(new_n886), .A2(new_n898), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n429), .A2(new_n868), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n444), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n431), .B(new_n1167), .C1(new_n442), .C2(new_n443), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n935), .B2(G330), .ZN(new_n1176));
  INV_X1    g0976(.A(G330), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1177), .B(new_n1174), .C1(new_n918), .C2(new_n934), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1166), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n884), .A2(new_n933), .A3(new_n881), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT38), .B1(new_n907), .B2(new_n877), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n932), .B1(new_n901), .B2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1180), .A2(new_n932), .B1(new_n1182), .B2(KEYINPUT40), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1174), .B1(new_n1183), .B2(new_n1177), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n935), .A2(G330), .A3(new_n1175), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n899), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1175), .A2(new_n794), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n801), .B1(G50), .B2(new_n821), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n756), .B2(new_n747), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n765), .A2(new_n1146), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n760), .A2(G132), .B1(new_n775), .B2(new_n1141), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n1147), .B2(new_n825), .C1(new_n1090), .C2(new_n740), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(G137), .C2(new_n831), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT59), .Z(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1196), .B2(KEYINPUT119), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(KEYINPUT119), .B2(new_n1196), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n278), .A2(new_n293), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G283), .B2(new_n770), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n957), .B(new_n1201), .C1(G107), .C2(new_n780), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n355), .B2(new_n753), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n761), .A2(new_n390), .B1(new_n762), .B2(new_n357), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n825), .A2(new_n540), .B1(new_n747), .B2(new_n202), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1199), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT117), .Z(new_n1212));
  NAND4_X1  g1012(.A1(new_n1198), .A2(new_n1209), .A3(new_n1210), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1189), .B1(new_n1213), .B2(new_n738), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1188), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT120), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1187), .A2(new_n800), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1117), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1135), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1187), .A2(KEYINPUT57), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n681), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1222), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(G375));
  NAND2_X1  g1026(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1007), .B(KEYINPUT121), .Z(new_n1228));
  NAND3_X1  g1028(.A1(new_n1119), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n865), .A2(new_n793), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n801), .B1(G68), .B2(new_n821), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n320), .B(new_n956), .C1(G303), .C2(new_n770), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n362), .B2(new_n753), .C1(new_n777), .C2(new_n765), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n760), .A2(G116), .B1(new_n775), .B2(G97), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n1051), .C1(new_n965), .C2(new_n825), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n766), .A2(new_n961), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n831), .A2(G150), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n744), .A2(G132), .B1(new_n775), .B2(G159), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G50), .A2(new_n774), .B1(new_n760), .B2(new_n1141), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n320), .B1(new_n755), .B2(new_n1146), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G58), .B2(new_n748), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1233), .A2(new_n1235), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1231), .B1(new_n1243), .B2(new_n738), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1230), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1115), .B2(new_n799), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1229), .A2(new_n1247), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT122), .Z(G381));
  OR2_X1    g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G384), .A2(G378), .A3(new_n1250), .A4(G390), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1251), .A2(G375), .A3(G387), .A4(G381), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT123), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1252), .B(new_n1253), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n1187), .A2(new_n800), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1225), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n681), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT57), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1261), .B2(new_n1222), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1257), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G378), .ZN(new_n1264));
  INV_X1    g1064(.A(G343), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(G213), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(G213), .B1(new_n1268), .B2(KEYINPUT124), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(KEYINPUT124), .B2(new_n1268), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G407), .A2(new_n1270), .ZN(G409));
  OAI211_X1 g1071(.A(new_n978), .B(G390), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(G393), .B(new_n808), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G390), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1272), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1280), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1220), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1216), .B1(new_n1187), .B2(new_n800), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1187), .A2(new_n1222), .A3(new_n1228), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1264), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT60), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(new_n681), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1227), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1293), .B2(new_n1247), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(new_n1246), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  AND4_X1   g1097(.A1(KEYINPUT62), .A2(new_n1288), .A3(new_n1266), .A4(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1267), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1297), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1267), .A2(G2897), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1297), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1294), .A2(new_n1296), .A3(KEYINPUT125), .A4(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1297), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1306), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G378), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1263), .B2(G378), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1308), .B(new_n1310), .C1(new_n1312), .C2(new_n1267), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1282), .B1(new_n1302), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1281), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1273), .A2(new_n1274), .B1(new_n1277), .B2(new_n1272), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1288), .A2(new_n1266), .B1(new_n1309), .B2(new_n1306), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1308), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1300), .A2(new_n1297), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1316), .A2(new_n1326), .ZN(G405));
  NAND2_X1  g1127(.A1(G375), .A2(new_n1264), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1283), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1297), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1328), .A2(new_n1309), .A3(new_n1283), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1282), .B(new_n1332), .ZN(G402));
endmodule


