

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  XNOR2_X1 U369 ( .A(n412), .B(n411), .ZN(n392) );
  XNOR2_X1 U370 ( .A(KEYINPUT78), .B(G110), .ZN(n420) );
  XNOR2_X1 U371 ( .A(KEYINPUT4), .B(KEYINPUT68), .ZN(n410) );
  AND2_X1 U372 ( .A1(n526), .A2(n739), .ZN(n405) );
  NOR2_X2 U373 ( .A1(n524), .A2(n632), .ZN(n526) );
  XNOR2_X2 U374 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n475) );
  OR2_X2 U375 ( .A1(n688), .A2(n598), .ZN(n605) );
  NAND2_X2 U376 ( .A1(n357), .A2(n655), .ZN(n373) );
  XNOR2_X2 U377 ( .A(n370), .B(n358), .ZN(n357) );
  AND2_X2 U378 ( .A1(n523), .A2(n522), .ZN(n632) );
  XNOR2_X2 U379 ( .A(n434), .B(G902), .ZN(n596) );
  XOR2_X2 U380 ( .A(n463), .B(n462), .Z(n358) );
  XOR2_X2 U381 ( .A(n614), .B(n613), .Z(n348) );
  XOR2_X2 U382 ( .A(KEYINPUT71), .B(KEYINPUT48), .Z(n364) );
  NOR2_X1 U383 ( .A1(n511), .A2(n678), .ZN(n510) );
  XNOR2_X2 U384 ( .A(n372), .B(n475), .ZN(n511) );
  XOR2_X1 U385 ( .A(G131), .B(G137), .Z(n412) );
  XNOR2_X1 U386 ( .A(n426), .B(n417), .ZN(n625) );
  BUF_X1 U387 ( .A(n501), .Z(n670) );
  BUF_X1 U388 ( .A(G143), .Z(n353) );
  NOR2_X1 U389 ( .A1(n612), .A2(n693), .ZN(n360) );
  INV_X1 U390 ( .A(n550), .ZN(n656) );
  NAND2_X2 U391 ( .A1(n520), .A2(n554), .ZN(n669) );
  NAND2_X1 U392 ( .A1(n647), .A2(n645), .ZN(n578) );
  NAND2_X1 U393 ( .A1(n360), .A2(G475), .ZN(n352) );
  NOR2_X1 U394 ( .A1(n641), .A2(n582), .ZN(n583) );
  AND2_X1 U395 ( .A1(n383), .A2(n382), .ZN(n363) );
  NOR2_X1 U396 ( .A1(n543), .A2(n552), .ZN(n544) );
  BUF_X1 U397 ( .A(n536), .Z(n674) );
  XNOR2_X1 U398 ( .A(G478), .B(n496), .ZN(n517) );
  NOR2_X1 U399 ( .A1(G902), .A2(n712), .ZN(n496) );
  XNOR2_X1 U400 ( .A(n376), .B(n374), .ZN(n614) );
  XNOR2_X1 U401 ( .A(n729), .B(n377), .ZN(n376) );
  XNOR2_X1 U402 ( .A(n483), .B(n375), .ZN(n374) );
  XNOR2_X1 U403 ( .A(G134), .B(KEYINPUT70), .ZN(n411) );
  XNOR2_X1 U404 ( .A(G119), .B(G128), .ZN(n431) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(G60) );
  INV_X1 U406 ( .A(KEYINPUT60), .ZN(n349) );
  NAND2_X1 U407 ( .A1(n351), .A2(n628), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n352), .B(n348), .ZN(n351) );
  NOR2_X2 U409 ( .A1(n355), .A2(n622), .ZN(n529) );
  XNOR2_X2 U410 ( .A(n400), .B(KEYINPUT35), .ZN(n355) );
  BUF_X1 U411 ( .A(n569), .Z(n354) );
  INV_X2 U412 ( .A(G143), .ZN(n365) );
  XNOR2_X2 U413 ( .A(n556), .B(KEYINPUT1), .ZN(n501) );
  BUF_X1 U414 ( .A(n663), .Z(n356) );
  XNOR2_X1 U415 ( .A(n448), .B(n447), .ZN(n663) );
  NOR2_X2 U416 ( .A1(n567), .A2(n670), .ZN(n650) );
  XNOR2_X2 U417 ( .A(n444), .B(KEYINPUT76), .ZN(n509) );
  NOR2_X2 U418 ( .A1(n501), .A2(n669), .ZN(n444) );
  INV_X1 U419 ( .A(n357), .ZN(n546) );
  NOR2_X1 U420 ( .A1(n612), .A2(n693), .ZN(n359) );
  BUF_X1 U421 ( .A(n450), .Z(n361) );
  NOR2_X2 U422 ( .A1(n612), .A2(n693), .ZN(n711) );
  XNOR2_X2 U423 ( .A(n611), .B(n610), .ZN(n693) );
  INV_X1 U424 ( .A(G237), .ZN(n460) );
  NOR2_X1 U425 ( .A1(n704), .A2(G902), .ZN(n428) );
  NOR2_X1 U426 ( .A1(n658), .A2(n465), .ZN(n384) );
  XOR2_X1 U427 ( .A(KEYINPUT104), .B(G107), .Z(n489) );
  AND2_X1 U428 ( .A1(n384), .A2(n551), .ZN(n381) );
  OR2_X1 U429 ( .A1(n384), .A2(n551), .ZN(n382) );
  INV_X1 U430 ( .A(KEYINPUT73), .ZN(n413) );
  XNOR2_X1 U431 ( .A(n729), .B(KEYINPUT24), .ZN(n396) );
  XNOR2_X1 U432 ( .A(n446), .B(KEYINPUT105), .ZN(n447) );
  NAND2_X1 U433 ( .A1(n394), .A2(n557), .ZN(n568) );
  XNOR2_X1 U434 ( .A(n555), .B(n395), .ZN(n394) );
  XNOR2_X1 U435 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n395) );
  XNOR2_X1 U436 ( .A(n516), .B(KEYINPUT103), .ZN(n518) );
  NOR2_X1 U437 ( .A1(G953), .A2(G237), .ZN(n480) );
  NAND2_X1 U438 ( .A1(G234), .A2(G237), .ZN(n466) );
  NAND2_X1 U439 ( .A1(n656), .A2(n655), .ZN(n659) );
  XNOR2_X1 U440 ( .A(n430), .B(n429), .ZN(n486) );
  XNOR2_X1 U441 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n429) );
  XNOR2_X1 U442 ( .A(G116), .B(G122), .ZN(n488) );
  XOR2_X1 U443 ( .A(G131), .B(KEYINPUT11), .Z(n482) );
  XNOR2_X1 U444 ( .A(n476), .B(n478), .ZN(n377) );
  XNOR2_X1 U445 ( .A(G113), .B(n353), .ZN(n476) );
  XNOR2_X1 U446 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n478) );
  XNOR2_X1 U447 ( .A(n477), .B(n479), .ZN(n375) );
  XNOR2_X1 U448 ( .A(G140), .B(KEYINPUT10), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n426), .B(n406), .ZN(n704) );
  XNOR2_X1 U450 ( .A(n425), .B(n457), .ZN(n406) );
  XOR2_X1 U451 ( .A(G101), .B(G140), .Z(n424) );
  XOR2_X1 U452 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n452) );
  NAND2_X1 U453 ( .A1(n363), .A2(n380), .ZN(n681) );
  NAND2_X1 U454 ( .A1(n656), .A2(n381), .ZN(n380) );
  NOR2_X1 U455 ( .A1(n561), .A2(n379), .ZN(n562) );
  XNOR2_X1 U456 ( .A(KEYINPUT16), .B(G122), .ZN(n449) );
  XNOR2_X1 U457 ( .A(n615), .B(KEYINPUT124), .ZN(n616) );
  INV_X1 U458 ( .A(n575), .ZN(n497) );
  INV_X1 U459 ( .A(n568), .ZN(n570) );
  INV_X1 U460 ( .A(KEYINPUT99), .ZN(n512) );
  INV_X1 U461 ( .A(n368), .ZN(n648) );
  INV_X1 U462 ( .A(n369), .ZN(n646) );
  AND2_X1 U463 ( .A1(n741), .A2(n652), .ZN(n362) );
  INV_X1 U464 ( .A(n551), .ZN(n385) );
  NAND2_X1 U465 ( .A1(n699), .A2(n435), .ZN(n370) );
  NAND2_X1 U466 ( .A1(n711), .A2(G210), .ZN(n702) );
  XNOR2_X2 U467 ( .A(n487), .B(n410), .ZN(n458) );
  XNOR2_X2 U468 ( .A(n365), .B(G128), .ZN(n487) );
  XNOR2_X2 U469 ( .A(n366), .B(n440), .ZN(n665) );
  NOR2_X2 U470 ( .A1(n615), .A2(G902), .ZN(n366) );
  INV_X2 U471 ( .A(KEYINPUT64), .ZN(n422) );
  NOR2_X2 U472 ( .A1(n577), .A2(n550), .ZN(n548) );
  OR2_X2 U473 ( .A1(n556), .A2(n669), .ZN(n535) );
  NAND2_X1 U474 ( .A1(n403), .A2(n386), .ZN(n519) );
  NAND2_X1 U475 ( .A1(n515), .A2(n514), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n367), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U477 ( .A1(n703), .A2(n715), .ZN(n367) );
  NAND2_X1 U478 ( .A1(n405), .A2(n529), .ZN(n404) );
  OR2_X1 U479 ( .A1(n386), .A2(n647), .ZN(n368) );
  OR2_X1 U480 ( .A1(n386), .A2(n645), .ZN(n369) );
  XNOR2_X1 U481 ( .A(n510), .B(KEYINPUT31), .ZN(n386) );
  XNOR2_X2 U482 ( .A(n371), .B(n459), .ZN(n699) );
  XNOR2_X2 U483 ( .A(n723), .B(n456), .ZN(n371) );
  NAND2_X1 U484 ( .A1(n569), .A2(n474), .ZN(n372) );
  XNOR2_X2 U485 ( .A(n373), .B(KEYINPUT19), .ZN(n569) );
  NAND2_X1 U486 ( .A1(n518), .A2(n517), .ZN(n645) );
  NAND2_X1 U487 ( .A1(n518), .A2(n378), .ZN(n379) );
  AND2_X1 U488 ( .A1(n517), .A2(n655), .ZN(n378) );
  NAND2_X1 U489 ( .A1(n550), .A2(n385), .ZN(n383) );
  AND2_X2 U490 ( .A1(n519), .A2(n578), .ZN(n524) );
  NOR2_X2 U491 ( .A1(n618), .A2(n715), .ZN(n620) );
  XNOR2_X2 U492 ( .A(n450), .B(n449), .ZN(n723) );
  XNOR2_X2 U493 ( .A(n388), .B(n387), .ZN(n450) );
  XNOR2_X2 U494 ( .A(n389), .B(n413), .ZN(n387) );
  XNOR2_X2 U495 ( .A(n391), .B(n390), .ZN(n388) );
  XNOR2_X2 U496 ( .A(G119), .B(KEYINPUT3), .ZN(n389) );
  XNOR2_X2 U497 ( .A(G101), .B(KEYINPUT74), .ZN(n390) );
  XNOR2_X2 U498 ( .A(G116), .B(G113), .ZN(n391) );
  XNOR2_X2 U499 ( .A(n728), .B(G146), .ZN(n426) );
  XNOR2_X2 U500 ( .A(n458), .B(n392), .ZN(n728) );
  INV_X1 U501 ( .A(n690), .ZN(n597) );
  XNOR2_X1 U502 ( .A(n607), .B(KEYINPUT85), .ZN(n690) );
  AND2_X2 U503 ( .A1(n393), .A2(n362), .ZN(n607) );
  XNOR2_X1 U504 ( .A(n588), .B(n364), .ZN(n393) );
  XNOR2_X2 U505 ( .A(n398), .B(n396), .ZN(n615) );
  XNOR2_X2 U506 ( .A(n453), .B(n397), .ZN(n729) );
  XNOR2_X2 U507 ( .A(n399), .B(n407), .ZN(n398) );
  NAND2_X1 U508 ( .A1(n486), .A2(G221), .ZN(n399) );
  NAND2_X1 U509 ( .A1(n401), .A2(n497), .ZN(n400) );
  XNOR2_X1 U510 ( .A(n402), .B(KEYINPUT34), .ZN(n401) );
  NOR2_X2 U511 ( .A1(n663), .A2(n511), .ZN(n402) );
  NOR2_X1 U512 ( .A1(n403), .A2(n645), .ZN(n633) );
  NOR2_X1 U513 ( .A1(n403), .A2(n647), .ZN(n638) );
  XNOR2_X2 U514 ( .A(n508), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U515 ( .A1(n404), .A2(n527), .ZN(n528) );
  XNOR2_X1 U516 ( .A(n722), .B(KEYINPUT75), .ZN(n457) );
  XNOR2_X2 U517 ( .A(n606), .B(KEYINPUT65), .ZN(n612) );
  OR2_X2 U518 ( .A1(n511), .A2(n498), .ZN(n500) );
  XNOR2_X1 U519 ( .A(n433), .B(KEYINPUT23), .ZN(n407) );
  NOR2_X1 U520 ( .A1(n689), .A2(n730), .ZN(n408) );
  AND2_X1 U521 ( .A1(n554), .A2(n553), .ZN(n409) );
  INV_X1 U522 ( .A(n552), .ZN(n553) );
  INV_X1 U523 ( .A(KEYINPUT38), .ZN(n547) );
  BUF_X1 U524 ( .A(n690), .Z(n730) );
  OR2_X1 U525 ( .A1(n731), .A2(G952), .ZN(n628) );
  INV_X1 U526 ( .A(KEYINPUT125), .ZN(n619) );
  XNOR2_X1 U527 ( .A(n558), .B(KEYINPUT42), .ZN(n742) );
  XOR2_X1 U528 ( .A(KEYINPUT5), .B(KEYINPUT77), .Z(n415) );
  AND2_X1 U529 ( .A1(n480), .A2(G210), .ZN(n414) );
  XNOR2_X1 U530 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U531 ( .A(n361), .B(n416), .ZN(n417) );
  INV_X1 U532 ( .A(G902), .ZN(n461) );
  NAND2_X1 U533 ( .A1(n625), .A2(n461), .ZN(n418) );
  XNOR2_X2 U534 ( .A(n418), .B(G472), .ZN(n536) );
  XNOR2_X1 U535 ( .A(n536), .B(KEYINPUT6), .ZN(n561) );
  INV_X1 U536 ( .A(n561), .ZN(n445) );
  XNOR2_X2 U537 ( .A(G104), .B(G107), .ZN(n419) );
  INV_X1 U538 ( .A(n419), .ZN(n421) );
  XNOR2_X1 U539 ( .A(n421), .B(n420), .ZN(n722) );
  XNOR2_X2 U540 ( .A(n422), .B(G953), .ZN(n731) );
  NAND2_X1 U541 ( .A1(G227), .A2(n731), .ZN(n423) );
  XNOR2_X1 U542 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U543 ( .A(KEYINPUT72), .B(G469), .ZN(n427) );
  XNOR2_X2 U544 ( .A(n428), .B(n427), .ZN(n556) );
  XOR2_X2 U545 ( .A(G146), .B(G125), .Z(n453) );
  NAND2_X1 U546 ( .A1(n731), .A2(G234), .ZN(n430) );
  XOR2_X1 U547 ( .A(G110), .B(G137), .Z(n432) );
  XNOR2_X1 U548 ( .A(n432), .B(n431), .ZN(n433) );
  INV_X1 U549 ( .A(KEYINPUT15), .ZN(n434) );
  INV_X1 U550 ( .A(n596), .ZN(n435) );
  NAND2_X1 U551 ( .A1(n435), .A2(G234), .ZN(n437) );
  XNOR2_X1 U552 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n436) );
  XNOR2_X1 U553 ( .A(n437), .B(n436), .ZN(n441) );
  NAND2_X1 U554 ( .A1(G217), .A2(n441), .ZN(n439) );
  INV_X1 U555 ( .A(KEYINPUT25), .ZN(n438) );
  XNOR2_X1 U556 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X2 U557 ( .A(n665), .ZN(n520) );
  NAND2_X1 U558 ( .A1(n441), .A2(G221), .ZN(n443) );
  INV_X1 U559 ( .A(KEYINPUT21), .ZN(n442) );
  XNOR2_X1 U560 ( .A(n443), .B(n442), .ZN(n554) );
  NAND2_X1 U561 ( .A1(n509), .A2(n445), .ZN(n448) );
  XOR2_X1 U562 ( .A(KEYINPUT33), .B(KEYINPUT91), .Z(n446) );
  NAND2_X1 U563 ( .A1(G224), .A2(n731), .ZN(n451) );
  XNOR2_X1 U564 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U565 ( .A(n453), .B(KEYINPUT92), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n459) );
  NAND2_X1 U568 ( .A1(n461), .A2(n460), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n464), .A2(G210), .ZN(n463) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n462) );
  NAND2_X1 U571 ( .A1(n464), .A2(G214), .ZN(n655) );
  INV_X1 U572 ( .A(n655), .ZN(n465) );
  XNOR2_X1 U573 ( .A(n466), .B(KEYINPUT14), .ZN(n468) );
  NAND2_X1 U574 ( .A1(G952), .A2(n468), .ZN(n467) );
  XNOR2_X1 U575 ( .A(KEYINPUT94), .B(n467), .ZN(n687) );
  NOR2_X1 U576 ( .A1(G953), .A2(n687), .ZN(n542) );
  NAND2_X1 U577 ( .A1(G902), .A2(n468), .ZN(n539) );
  INV_X1 U578 ( .A(G953), .ZN(n716) );
  NOR2_X1 U579 ( .A1(n716), .A2(G898), .ZN(n469) );
  XNOR2_X1 U580 ( .A(n469), .B(KEYINPUT95), .ZN(n724) );
  NOR2_X1 U581 ( .A1(n539), .A2(n724), .ZN(n470) );
  XNOR2_X1 U582 ( .A(n470), .B(KEYINPUT96), .ZN(n471) );
  OR2_X1 U583 ( .A1(n542), .A2(n471), .ZN(n473) );
  INV_X1 U584 ( .A(KEYINPUT97), .ZN(n472) );
  XNOR2_X1 U585 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U586 ( .A(G104), .B(G122), .Z(n477) );
  XOR2_X1 U587 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n479) );
  NAND2_X1 U588 ( .A1(G214), .A2(n480), .ZN(n481) );
  XNOR2_X1 U589 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U590 ( .A1(G902), .A2(n614), .ZN(n485) );
  XOR2_X1 U591 ( .A(KEYINPUT13), .B(G475), .Z(n484) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n516) );
  NAND2_X1 U593 ( .A1(n486), .A2(G217), .ZN(n495) );
  XNOR2_X1 U594 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n487), .B(G134), .ZN(n491) );
  XNOR2_X1 U596 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U597 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U599 ( .A(n495), .B(n494), .ZN(n712) );
  OR2_X1 U600 ( .A1(n516), .A2(n517), .ZN(n575) );
  NAND2_X1 U601 ( .A1(n516), .A2(n517), .ZN(n658) );
  INV_X1 U602 ( .A(n554), .ZN(n666) );
  OR2_X1 U603 ( .A1(n658), .A2(n666), .ZN(n498) );
  INV_X1 U604 ( .A(KEYINPUT22), .ZN(n499) );
  XNOR2_X2 U605 ( .A(n500), .B(n499), .ZN(n523) );
  INV_X1 U606 ( .A(n523), .ZN(n504) );
  NOR2_X1 U607 ( .A1(n674), .A2(n520), .ZN(n502) );
  NAND2_X1 U608 ( .A1(n670), .A2(n502), .ZN(n503) );
  NOR2_X1 U609 ( .A1(n504), .A2(n503), .ZN(n622) );
  INV_X1 U610 ( .A(n670), .ZN(n593) );
  NAND2_X1 U611 ( .A1(n593), .A2(n561), .ZN(n505) );
  NOR2_X1 U612 ( .A1(n520), .A2(n505), .ZN(n506) );
  XNOR2_X1 U613 ( .A(KEYINPUT80), .B(n506), .ZN(n507) );
  NAND2_X1 U614 ( .A1(n523), .A2(n507), .ZN(n508) );
  NAND2_X1 U615 ( .A1(n509), .A2(n674), .ZN(n678) );
  NOR2_X1 U616 ( .A1(n511), .A2(n535), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n515) );
  INV_X1 U618 ( .A(n674), .ZN(n514) );
  OR2_X1 U619 ( .A1(n518), .A2(n517), .ZN(n647) );
  AND2_X1 U620 ( .A1(n670), .A2(n520), .ZN(n521) );
  AND2_X1 U621 ( .A1(n521), .A2(n561), .ZN(n522) );
  INV_X1 U622 ( .A(KEYINPUT44), .ZN(n525) );
  NAND2_X1 U623 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n528), .B(KEYINPUT89), .ZN(n532) );
  NAND2_X1 U625 ( .A1(n529), .A2(n739), .ZN(n530) );
  NOR2_X1 U626 ( .A1(n530), .A2(KEYINPUT44), .ZN(n531) );
  NOR2_X1 U627 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U628 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n533) );
  XNOR2_X1 U629 ( .A(n534), .B(n533), .ZN(n688) );
  INV_X1 U630 ( .A(n535), .ZN(n545) );
  NAND2_X1 U631 ( .A1(n536), .A2(n655), .ZN(n538) );
  XOR2_X1 U632 ( .A(KEYINPUT30), .B(KEYINPUT107), .Z(n537) );
  XNOR2_X1 U633 ( .A(n538), .B(n537), .ZN(n543) );
  OR2_X1 U634 ( .A1(n731), .A2(n539), .ZN(n540) );
  NOR2_X1 U635 ( .A1(G900), .A2(n540), .ZN(n541) );
  NOR2_X1 U636 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n545), .A2(n544), .ZN(n577) );
  XNOR2_X2 U638 ( .A(n546), .B(n547), .ZN(n550) );
  XNOR2_X1 U639 ( .A(n548), .B(KEYINPUT39), .ZN(n589) );
  NOR2_X1 U640 ( .A1(n645), .A2(n589), .ZN(n549) );
  XNOR2_X1 U641 ( .A(n549), .B(KEYINPUT40), .ZN(n740) );
  XNOR2_X1 U642 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n551) );
  AND2_X1 U643 ( .A1(n665), .A2(n409), .ZN(n563) );
  NAND2_X1 U644 ( .A1(n563), .A2(n674), .ZN(n555) );
  XOR2_X1 U645 ( .A(n556), .B(KEYINPUT108), .Z(n557) );
  NOR2_X1 U646 ( .A1(n681), .A2(n568), .ZN(n558) );
  NOR2_X1 U647 ( .A1(n740), .A2(n742), .ZN(n560) );
  XNOR2_X1 U648 ( .A(KEYINPUT46), .B(KEYINPUT87), .ZN(n559) );
  XNOR2_X1 U649 ( .A(n560), .B(n559), .ZN(n587) );
  AND2_X1 U650 ( .A1(n563), .A2(n562), .ZN(n591) );
  INV_X1 U651 ( .A(n546), .ZN(n564) );
  NAND2_X1 U652 ( .A1(n591), .A2(n564), .ZN(n566) );
  XOR2_X1 U653 ( .A(KEYINPUT111), .B(KEYINPUT36), .Z(n565) );
  XNOR2_X1 U654 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U655 ( .A(n650), .B(KEYINPUT88), .ZN(n574) );
  NAND2_X1 U656 ( .A1(n570), .A2(n354), .ZN(n643) );
  XNOR2_X1 U657 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n571) );
  NAND2_X1 U658 ( .A1(n578), .A2(n571), .ZN(n572) );
  NOR2_X1 U659 ( .A1(n643), .A2(n572), .ZN(n573) );
  NOR2_X1 U660 ( .A1(n574), .A2(n573), .ZN(n585) );
  OR2_X1 U661 ( .A1(n546), .A2(n575), .ZN(n576) );
  NOR2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n641) );
  INV_X1 U663 ( .A(n578), .ZN(n660) );
  NAND2_X1 U664 ( .A1(n660), .A2(KEYINPUT47), .ZN(n579) );
  XOR2_X1 U665 ( .A(n579), .B(KEYINPUT83), .Z(n581) );
  NAND2_X1 U666 ( .A1(n643), .A2(KEYINPUT47), .ZN(n580) );
  NAND2_X1 U667 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U668 ( .A(n583), .B(KEYINPUT82), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n588) );
  OR2_X1 U671 ( .A1(n589), .A2(n647), .ZN(n590) );
  XNOR2_X1 U672 ( .A(KEYINPUT112), .B(n590), .ZN(n741) );
  XOR2_X1 U673 ( .A(KEYINPUT106), .B(n591), .Z(n592) );
  NOR2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U675 ( .A(n594), .B(KEYINPUT43), .Z(n595) );
  NAND2_X1 U676 ( .A1(n595), .A2(n546), .ZN(n652) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U678 ( .A(KEYINPUT2), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n599), .A2(KEYINPUT84), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n435), .A2(n600), .ZN(n603) );
  NAND2_X1 U681 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n601) );
  OR2_X1 U682 ( .A1(n435), .A2(n601), .ZN(n602) );
  AND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U685 ( .A(KEYINPUT79), .ZN(n611) );
  BUF_X1 U686 ( .A(n607), .Z(n608) );
  NAND2_X1 U687 ( .A1(n608), .A2(KEYINPUT2), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n688), .A2(n609), .ZN(n610) );
  INV_X1 U689 ( .A(KEYINPUT59), .ZN(n613) );
  INV_X1 U690 ( .A(n628), .ZN(n715) );
  NAND2_X1 U691 ( .A1(n711), .A2(G217), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(G66) );
  XOR2_X1 U694 ( .A(G110), .B(KEYINPUT116), .Z(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(G12) );
  XNOR2_X1 U696 ( .A(G122), .B(KEYINPUT127), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n355), .B(n623), .ZN(G24) );
  NAND2_X1 U698 ( .A1(n359), .A2(G472), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n624) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n631) );
  XNOR2_X1 U703 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n631), .B(n630), .ZN(G57) );
  XOR2_X1 U705 ( .A(G101), .B(n632), .Z(G3) );
  XOR2_X1 U706 ( .A(G104), .B(n633), .Z(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n635) );
  XNOR2_X1 U708 ( .A(G107), .B(KEYINPUT26), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(KEYINPUT27), .B(n636), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G9) );
  NOR2_X1 U712 ( .A1(n643), .A2(n647), .ZN(n640) );
  XNOR2_X1 U713 ( .A(G128), .B(KEYINPUT29), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(G30) );
  XNOR2_X1 U715 ( .A(n353), .B(n641), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n642), .B(KEYINPUT117), .ZN(G45) );
  NOR2_X1 U717 ( .A1(n643), .A2(n645), .ZN(n644) );
  XOR2_X1 U718 ( .A(G146), .B(n644), .Z(G48) );
  XOR2_X1 U719 ( .A(G113), .B(n646), .Z(G15) );
  XOR2_X1 U720 ( .A(KEYINPUT118), .B(n648), .Z(n649) );
  XNOR2_X1 U721 ( .A(G116), .B(n649), .ZN(G18) );
  XNOR2_X1 U722 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U724 ( .A(G140), .B(n652), .Z(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT119), .ZN(G42) );
  NOR2_X1 U726 ( .A1(n681), .A2(n356), .ZN(n654) );
  NOR2_X1 U727 ( .A1(G953), .A2(n654), .ZN(n697) );
  NOR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U729 ( .A1(n658), .A2(n657), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n664), .A2(n356), .ZN(n683) );
  XOR2_X1 U733 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n668) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n676) );
  NAND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT50), .ZN(n672) );
  XNOR2_X1 U738 ( .A(KEYINPUT121), .B(n672), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U742 ( .A(KEYINPUT51), .B(n679), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n684), .B(KEYINPUT122), .ZN(n685) );
  XNOR2_X1 U746 ( .A(KEYINPUT52), .B(n685), .ZN(n686) );
  NOR2_X1 U747 ( .A1(n687), .A2(n686), .ZN(n695) );
  BUF_X1 U748 ( .A(n688), .Z(n689) );
  XOR2_X1 U749 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n691) );
  NOR2_X1 U750 ( .A1(n408), .A2(n691), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U754 ( .A(KEYINPUT53), .B(n698), .Z(G75) );
  XOR2_X1 U755 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n700) );
  XOR2_X1 U756 ( .A(n700), .B(n699), .Z(n701) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n359), .A2(G469), .ZN(n709) );
  XNOR2_X1 U759 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n707) );
  BUF_X1 U760 ( .A(n704), .Z(n705) );
  XNOR2_X1 U761 ( .A(n705), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n715), .A2(n710), .ZN(G54) );
  NAND2_X1 U765 ( .A1(n360), .A2(G478), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(G63) );
  INV_X1 U768 ( .A(n689), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n718) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n719), .A2(G898), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n727) );
  XNOR2_X1 U774 ( .A(n723), .B(n722), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U776 ( .A(n727), .B(n726), .Z(G69) );
  XNOR2_X1 U777 ( .A(n728), .B(n729), .ZN(n733) );
  XNOR2_X1 U778 ( .A(n730), .B(n733), .ZN(n732) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(n737) );
  XNOR2_X1 U780 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U783 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U784 ( .A(KEYINPUT126), .B(n738), .ZN(G72) );
  XNOR2_X1 U785 ( .A(n739), .B(G119), .ZN(G21) );
  XOR2_X1 U786 ( .A(n740), .B(G131), .Z(G33) );
  XNOR2_X1 U787 ( .A(G134), .B(n741), .ZN(G36) );
  XOR2_X1 U788 ( .A(G137), .B(n742), .Z(G39) );
endmodule

