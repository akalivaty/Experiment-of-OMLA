//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G113), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OR3_X1    g036(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT67), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT67), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(new_n462), .B(new_n463), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n468), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n461), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G112), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  NOR3_X1   g053(.A1(new_n477), .A2(new_n461), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n468), .B2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT69), .B1(new_n483), .B2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n468), .A2(new_n476), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n479), .B(new_n484), .C1(G124), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(KEYINPUT69), .A3(G136), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(new_n471), .A2(G138), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT4), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n476), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n485), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT70), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT70), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT6), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n509), .A2(G543), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT71), .B1(new_n512), .B2(G50), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n502), .A2(new_n511), .A3(new_n509), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI211_X1 g090(.A(new_n508), .B(new_n513), .C1(G88), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(KEYINPUT71), .A3(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n515), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI211_X1 g100(.A(new_n523), .B(new_n524), .C1(new_n502), .C2(new_n525), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT72), .B(G51), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n512), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(new_n526), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G52), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(G90), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  XNOR2_X1  g112(.A(KEYINPUT75), .B(G81), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n515), .A2(new_n539), .B1(new_n512), .B2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n499), .A2(new_n501), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  INV_X1    g117(.A(G68), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n498), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  OAI221_X1 g121(.A(new_n546), .B1(new_n543), .B2(new_n498), .C1(new_n541), .C2(new_n542), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n506), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n514), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT79), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT79), .B1(new_n499), .B2(new_n501), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n561), .B1(new_n564), .B2(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n559), .B1(new_n565), .B2(new_n510), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n541), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT79), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(G65), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n510), .B1(new_n570), .B2(new_n560), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n558), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n509), .A2(G53), .A3(G543), .A4(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT76), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n512), .A2(new_n580), .A3(new_n581), .A4(G53), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT77), .B1(new_n574), .B2(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT78), .B1(new_n579), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n573), .B1(new_n585), .B2(new_n586), .ZN(G299));
  NAND2_X1  g162(.A1(new_n515), .A2(G87), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n512), .A2(G49), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n502), .A2(G61), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n592), .A2(KEYINPUT81), .B1(G73), .B2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n507), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n509), .A2(G543), .A3(new_n511), .ZN(new_n597));
  INV_X1    g172(.A(G48), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n514), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n515), .A2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n512), .A2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(new_n507), .C2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT82), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n515), .A2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n564), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(new_n510), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n512), .A2(G54), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n608), .B1(new_n616), .B2(G868), .ZN(G284));
  XNOR2_X1  g192(.A(G284), .B(KEYINPUT83), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G168), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n622));
  AOI211_X1 g197(.A(new_n559), .B(new_n510), .C1(new_n570), .C2(new_n560), .ZN(new_n623));
  OAI22_X1  g198(.A1(new_n622), .A2(new_n623), .B1(new_n557), .B2(new_n514), .ZN(new_n624));
  INV_X1    g199(.A(new_n583), .ZN(new_n625));
  NOR3_X1   g200(.A1(new_n574), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT9), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n577), .B1(new_n574), .B2(KEYINPUT9), .ZN(new_n628));
  OAI22_X1  g203(.A1(new_n625), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n579), .A2(new_n584), .A3(KEYINPUT78), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n621), .B1(new_n633), .B2(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT84), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(KEYINPUT84), .B2(new_n620), .ZN(G297));
  OAI21_X1  g211(.A(new_n635), .B1(KEYINPUT84), .B2(new_n620), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n616), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n549), .A2(new_n619), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n615), .A2(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g218(.A1(new_n465), .A2(new_n467), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n472), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n485), .A2(G123), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n476), .A2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n483), .B2(G135), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2096), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n662), .A2(KEYINPUT87), .A3(KEYINPUT14), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT87), .B1(new_n662), .B2(KEYINPUT14), .ZN(new_n664));
  OAI22_X1  g239(.A1(new_n663), .A2(new_n664), .B1(new_n658), .B2(new_n661), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT16), .Z(new_n666));
  XOR2_X1   g241(.A(G2451), .B(G2454), .Z(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n667), .B(new_n668), .Z(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1341), .B(G1348), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n669), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n670), .A2(KEYINPUT88), .A3(new_n672), .A4(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G14), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n670), .A2(new_n673), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n671), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G401));
  XNOR2_X1  g258(.A(KEYINPUT92), .B(G2096), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  XNOR2_X1  g261(.A(G2067), .B(G2678), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2072), .B(G2078), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT89), .Z(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(KEYINPUT18), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(KEYINPUT18), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(KEYINPUT17), .ZN(new_n693));
  INV_X1    g268(.A(new_n686), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n693), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n686), .B1(new_n693), .B2(new_n687), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n688), .B(KEYINPUT90), .Z(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n687), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  INV_X1    g275(.A(G2100), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n701), .B1(new_n696), .B2(new_n700), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n685), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n702), .A3(new_n684), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(G227));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1971), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT19), .ZN(new_n713));
  XOR2_X1   g288(.A(G1956), .B(G2474), .Z(new_n714));
  XOR2_X1   g289(.A(G1961), .B(G1966), .Z(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n715), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT19), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n712), .B(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n722), .A2(KEYINPUT20), .A3(new_n714), .A4(new_n715), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n713), .A2(new_n716), .A3(new_n719), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n717), .A2(new_n720), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G1991), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(G1991), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(G1996), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(G1996), .B1(new_n726), .B2(new_n727), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n711), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n729), .A2(new_n711), .A3(new_n730), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n710), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n733), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n735), .A2(new_n709), .A3(new_n731), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(G229));
  XNOR2_X1  g313(.A(KEYINPUT94), .B(G16), .ZN(new_n739));
  MUX2_X1   g314(.A(G22), .B(G303), .S(new_n739), .Z(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G6), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n600), .B2(new_n743), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT32), .B(G1981), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G23), .B(G288), .S(G16), .Z(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT33), .B(G1976), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n742), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT34), .Z(new_n752));
  MUX2_X1   g327(.A(G24), .B(G290), .S(new_n739), .Z(new_n753));
  INV_X1    g328(.A(G1986), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(KEYINPUT93), .A2(G29), .ZN(new_n756));
  NOR2_X1   g331(.A1(KEYINPUT93), .A2(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G25), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n485), .A2(G119), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n476), .A2(G107), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n483), .B2(G131), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n760), .B1(new_n765), .B2(new_n759), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT35), .B(G1991), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n752), .A2(new_n755), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT36), .ZN(new_n771));
  INV_X1    g346(.A(G20), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n739), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n633), .B2(new_n743), .ZN(new_n776));
  INV_X1    g351(.A(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G32), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n483), .A2(G141), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n472), .A2(G105), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT103), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n485), .A2(G129), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT26), .Z(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n779), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT27), .B(G1996), .Z(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NOR2_X1   g366(.A1(G164), .A2(new_n759), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G27), .B2(new_n759), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n791), .B1(new_n794), .B2(G2078), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n790), .B(new_n795), .C1(G2078), .C2(new_n794), .ZN(new_n796));
  NOR2_X1   g371(.A1(G5), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G171), .B2(G16), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G1961), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(G1961), .ZN(new_n800));
  NOR2_X1   g375(.A1(G168), .A2(new_n743), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n743), .B2(G21), .ZN(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n799), .B(new_n804), .C1(new_n803), .C2(new_n802), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT31), .B(G11), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT30), .B(G28), .Z(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G29), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n653), .B2(new_n758), .ZN(new_n809));
  INV_X1    g384(.A(G2084), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT24), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(G34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(G34), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n759), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G29), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n474), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n809), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n759), .A2(G26), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT99), .B(KEYINPUT28), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n483), .A2(G140), .ZN(new_n821));
  OR2_X1    g396(.A1(G104), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT98), .ZN(new_n824));
  INV_X1    g399(.A(G128), .ZN(new_n825));
  INV_X1    g400(.A(new_n485), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n820), .B1(new_n828), .B2(new_n815), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT100), .B(G2067), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AOI211_X1 g406(.A(new_n817), .B(new_n831), .C1(new_n810), .C2(new_n816), .ZN(new_n832));
  MUX2_X1   g407(.A(G19), .B(new_n549), .S(new_n739), .Z(new_n833));
  XOR2_X1   g408(.A(KEYINPUT97), .B(G1341), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n796), .A2(new_n805), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n759), .A2(G35), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G162), .B2(new_n759), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT29), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2090), .ZN(new_n840));
  NOR2_X1   g415(.A1(G4), .A2(G16), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT95), .Z(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n615), .B2(new_n743), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT96), .Z(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(G1348), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n815), .A2(G33), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n472), .A2(G103), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT25), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n483), .B2(G139), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n644), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n476), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n846), .B1(new_n855), .B2(new_n815), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT102), .B(G2072), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G1348), .ZN(new_n859));
  INV_X1    g434(.A(new_n844), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR4_X1   g436(.A1(new_n836), .A2(new_n840), .A3(new_n845), .A4(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n771), .A2(new_n778), .A3(new_n862), .ZN(G311));
  NAND3_X1  g438(.A1(new_n771), .A2(new_n778), .A3(new_n862), .ZN(G150));
  NAND2_X1  g439(.A1(new_n616), .A2(G559), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n549), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n540), .A2(new_n548), .A3(KEYINPUT106), .ZN(new_n868));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  INV_X1    g444(.A(G55), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n514), .A2(new_n869), .B1(new_n597), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(G80), .A2(G543), .ZN(new_n872));
  INV_X1    g447(.A(G67), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n541), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(new_n506), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n874), .B2(new_n506), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n867), .A2(new_n868), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n866), .A3(new_n549), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n865), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g460(.A(G860), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n880), .A2(G860), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT37), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(G145));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n485), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n476), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n483), .B2(G142), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n646), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n765), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n854), .A2(KEYINPUT107), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n851), .B2(new_n853), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n828), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G164), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n828), .A2(new_n496), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n787), .ZN(new_n908));
  INV_X1    g483(.A(new_n787), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n900), .A2(new_n903), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n910), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n912), .A2(new_n902), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n898), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n653), .B(new_n474), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n488), .B(new_n916), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n912), .A2(new_n913), .B1(new_n899), .B2(new_n902), .ZN(new_n918));
  INV_X1    g493(.A(new_n898), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n908), .A2(new_n903), .A3(new_n910), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n915), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n891), .B(new_n922), .C1(new_n923), .C2(KEYINPUT108), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n926), .B(new_n927), .Z(G395));
  NAND2_X1  g503(.A1(new_n880), .A2(new_n619), .ZN(new_n929));
  XOR2_X1   g504(.A(G288), .B(KEYINPUT112), .Z(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G290), .A2(G303), .ZN(new_n932));
  NAND2_X1  g507(.A1(G166), .A2(new_n606), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n933), .A3(G305), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G305), .B1(new_n932), .B2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n930), .A3(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT113), .A3(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT113), .B(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n641), .B(new_n882), .ZN(new_n944));
  NAND3_X1  g519(.A1(G299), .A2(KEYINPUT110), .A3(new_n615), .ZN(new_n945));
  NAND2_X1  g520(.A1(G299), .A2(KEYINPUT110), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n573), .C1(new_n585), .C2(new_n586), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n616), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n944), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n616), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n631), .A2(new_n632), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(new_n953), .B2(new_n573), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n945), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT41), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n958), .A3(new_n945), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n951), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n951), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n950), .B1(new_n962), .B2(new_n944), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n943), .B(new_n963), .Z(new_n964));
  OAI21_X1  g539(.A(new_n929), .B1(new_n964), .B2(new_n619), .ZN(G295));
  OAI21_X1  g540(.A(new_n929), .B1(new_n964), .B2(new_n619), .ZN(G331));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n937), .A2(new_n939), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n879), .A2(new_n881), .A3(G301), .ZN(new_n969));
  AOI21_X1  g544(.A(G301), .B1(new_n879), .B2(new_n881), .ZN(new_n970));
  OAI21_X1  g545(.A(G286), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n882), .A2(G171), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n879), .A2(new_n881), .A3(G301), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(G168), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n960), .B2(new_n961), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n974), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n945), .A3(new_n949), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n968), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n968), .A3(new_n978), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n980), .A2(new_n891), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n959), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n958), .B1(new_n949), .B2(new_n945), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n975), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n978), .ZN(new_n988));
  AOI21_X1  g563(.A(G37), .B1(new_n988), .B2(new_n940), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n967), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n989), .A2(new_n981), .A3(new_n983), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n980), .A2(new_n891), .A3(new_n981), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n982), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n967), .B2(new_n995), .ZN(G397));
  OR2_X1    g571(.A1(G305), .A2(G1981), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(G305), .A2(G1981), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  AND2_X1   g578(.A1(G160), .A2(G40), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n491), .B2(new_n495), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1002), .B(new_n1003), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT116), .B1(new_n1007), .B2(G8), .ZN(new_n1008));
  OAI22_X1  g583(.A1(new_n1000), .A2(new_n1001), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g586(.A(new_n1011), .B1(new_n1010), .B2(G288), .C1(new_n1008), .C2(new_n1006), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1013));
  INV_X1    g588(.A(G288), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(G1976), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1009), .B(new_n1012), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n496), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1004), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n741), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1005), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1005), .A2(KEYINPUT117), .A3(new_n1026), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(new_n1004), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1025), .B1(new_n1032), .B2(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  AOI22_X1  g610(.A1(G303), .A2(G8), .B1(new_n1035), .B2(KEYINPUT55), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(KEYINPUT55), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1036), .B(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1030), .A2(new_n1042), .A3(new_n1004), .A4(new_n1027), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1003), .B1(new_n1025), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1018), .A2(new_n1040), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G168), .A2(new_n1003), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1030), .A2(new_n1004), .A3(new_n1027), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1050), .A2(new_n810), .B1(new_n1024), .B2(new_n803), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT51), .B(new_n1048), .C1(new_n1051), .C2(new_n1003), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1024), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1054), .A2(G1966), .B1(G2084), .B2(new_n1049), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1053), .B(G8), .C1(new_n1055), .C2(G286), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1047), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1050), .A2(G1961), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1024), .B2(G2078), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT123), .B(new_n1061), .C1(new_n1024), .C2(G2078), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1024), .A2(new_n1061), .A3(G2078), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1060), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1052), .A2(new_n1056), .A3(new_n1069), .A4(new_n1057), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1059), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1051), .A2(new_n1003), .A3(G286), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1046), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n997), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G288), .A2(G1976), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1009), .B2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1017), .A2(new_n1045), .B1(new_n1078), .B2(new_n1013), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1044), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1039), .B1(new_n1044), .B2(new_n1080), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT119), .B1(new_n1084), .B2(new_n1017), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1044), .A2(new_n1080), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n1039), .A3(new_n1081), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1018), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1045), .A2(new_n1072), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1079), .B1(new_n1091), .B2(KEYINPUT63), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1054), .A2(new_n1093), .B1(new_n1032), .B2(new_n777), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n573), .A2(new_n1096), .A3(new_n629), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT120), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1049), .A2(new_n859), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1007), .A2(G2067), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n616), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1105), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n616), .C1(new_n1108), .C2(KEYINPUT60), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT60), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n615), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1109), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1110), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1007), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT58), .B(G1341), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1024), .A2(G1996), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n550), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT59), .Z(new_n1120));
  NOR3_X1   g695(.A1(new_n1114), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1094), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n1098), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT61), .B1(new_n1123), .B2(new_n1102), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1102), .A2(KEYINPUT121), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1124), .B1(new_n1101), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1107), .B1(new_n1121), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT124), .B(G2078), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1060), .A2(new_n1064), .A3(new_n1065), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(G171), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1067), .A2(G171), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(KEYINPUT125), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1067), .A2(new_n1139), .A3(G171), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1135), .A2(G171), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1132), .B1(new_n1068), .B2(new_n1142), .ZN(new_n1143));
  AND4_X1   g718(.A1(new_n1058), .A2(new_n1018), .A3(new_n1040), .A4(new_n1045), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1075), .B(new_n1092), .C1(new_n1131), .C2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1020), .A2(new_n1021), .A3(new_n1004), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n828), .B(G2067), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n787), .B(G1996), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n765), .B(new_n768), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n606), .B(new_n754), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1146), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1147), .B1(new_n1149), .B2(new_n787), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT46), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1147), .A2(G1996), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n765), .A2(new_n768), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1151), .A2(new_n1164), .B1(G2067), .B2(new_n904), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1148), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT48), .ZN(new_n1167));
  NOR2_X1   g742(.A1(G290), .A2(G1986), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1169), .B2(new_n1147), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(KEYINPUT48), .A3(new_n1148), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1170), .B(new_n1171), .C1(new_n1147), .C2(new_n1153), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1163), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1157), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g749(.A1(new_n981), .A2(new_n891), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n982), .B1(new_n1176), .B2(new_n979), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n989), .A2(new_n981), .A3(new_n983), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g753(.A1(new_n705), .A2(new_n707), .A3(G319), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n1180), .A2(new_n736), .A3(new_n734), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1181), .B1(new_n678), .B2(new_n681), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1182), .B1(new_n924), .B2(new_n925), .ZN(new_n1183));
  INV_X1    g757(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g758(.A(KEYINPUT126), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1186));
  AOI211_X1 g760(.A(new_n1186), .B(new_n1183), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1187), .ZN(G308));
  OAI21_X1  g762(.A(new_n1186), .B1(new_n995), .B2(new_n1183), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n1179), .A2(KEYINPUT126), .A3(new_n1184), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1190), .ZN(G225));
endmodule


