//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G134), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT66), .ZN(new_n193));
  OAI21_X1  g007(.A(G137), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(G137), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n189), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(KEYINPUT66), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n189), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n197), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(new_n199), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n195), .B1(new_n207), .B2(G137), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n206), .B(new_n202), .C1(new_n208), .C2(new_n189), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(KEYINPUT67), .B(G131), .C1(new_n197), .C2(new_n203), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT0), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  AOI211_X1 g033(.A(new_n212), .B(new_n215), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n216), .B2(G143), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(KEYINPUT64), .A3(G146), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n222), .A2(new_n223), .B1(G143), .B2(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n215), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n227), .A3(new_n215), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n220), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n210), .A2(new_n211), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n217), .A2(new_n219), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n214), .A2(KEYINPUT68), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(G143), .B2(new_n216), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n231), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n222), .A2(new_n223), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(new_n236), .A3(G128), .A4(new_n217), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n201), .B1(G134), .B2(new_n200), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n238), .A2(new_n240), .B1(new_n241), .B2(G131), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n209), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n245), .A3(new_n209), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT30), .B1(new_n230), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(G116), .B(G119), .Z(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  XOR2_X1   g064(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n210), .A2(new_n211), .A3(new_n229), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n243), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n242), .A2(new_n245), .A3(new_n209), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n245), .B1(new_n242), .B2(new_n209), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n253), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n251), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  INV_X1    g078(.A(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n266), .B(new_n267), .Z(new_n268));
  AOI21_X1  g082(.A(new_n188), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  AOI211_X1 g084(.A(KEYINPUT31), .B(new_n270), .C1(new_n256), .C2(new_n261), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n260), .B2(new_n251), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n253), .A2(new_n243), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n252), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n251), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n272), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n268), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n269), .A2(new_n271), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n256), .A2(new_n261), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT31), .B1(new_n284), .B2(new_n270), .ZN(new_n285));
  INV_X1    g099(.A(new_n279), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n270), .B1(new_n256), .B2(new_n261), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n188), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT32), .A3(new_n281), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n278), .A3(new_n268), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n256), .A2(new_n261), .A3(new_n270), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n259), .A2(new_n252), .A3(new_n253), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n273), .A2(new_n296), .B1(new_n277), .B2(new_n272), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n270), .A2(new_n292), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G472), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n283), .A2(new_n290), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n214), .A3(G119), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n214), .A2(G119), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT68), .B(G128), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n304), .B1(new_n309), .B2(new_n303), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n311));
  INV_X1    g125(.A(G110), .ZN(new_n312));
  OR3_X1    g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G125), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G140), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n314), .A2(KEYINPUT73), .A3(G140), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n319), .B2(G125), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT16), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n317), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G146), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n319), .A3(G125), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT73), .B1(new_n314), .B2(G140), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n315), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n316), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n216), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n309), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n313), .A2(new_n332), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n310), .A2(new_n312), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n333), .A2(new_n334), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT74), .B1(new_n310), .B2(new_n312), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n325), .A2(KEYINPUT75), .A3(G146), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n330), .B2(new_n216), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n314), .A2(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n320), .A2(new_n348), .A3(new_n216), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n337), .B1(new_n343), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n337), .C1(new_n343), .C2(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G953), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(G221), .A3(G234), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT77), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G137), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n295), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n351), .A2(new_n360), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n355), .B2(new_n360), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT25), .A3(new_n362), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n362), .B2(G234), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT71), .Z(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(G902), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n370), .A2(new_n373), .B1(new_n374), .B2(new_n368), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n302), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n356), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT88), .A2(G143), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n218), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n263), .A2(new_n382), .A3(new_n218), .A4(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n206), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT17), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(G131), .A3(new_n385), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n389), .A2(new_n388), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n326), .A2(new_n390), .A3(new_n391), .A4(new_n331), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n329), .A2(G146), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n349), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n384), .A2(KEYINPUT18), .A3(G131), .A4(new_n385), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT89), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n396), .A2(new_n349), .B1(new_n386), .B2(new_n398), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT89), .B1(new_n404), .B2(new_n400), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n392), .B(new_n395), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n401), .A2(new_n402), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(KEYINPUT89), .A3(new_n400), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n320), .A2(new_n348), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT19), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(KEYINPUT19), .B2(new_n329), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n413), .A2(new_n216), .B1(new_n387), .B2(new_n389), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n347), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n395), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT90), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n408), .A2(new_n409), .B1(new_n347), .B2(new_n414), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n406), .B(new_n418), .C1(new_n419), .C2(new_n395), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n425));
  INV_X1    g239(.A(new_n422), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n417), .B2(new_n420), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n428), .B(new_n422), .C1(new_n407), .C2(new_n416), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n410), .A2(new_n392), .ZN(new_n433));
  INV_X1    g247(.A(new_n395), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT92), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT93), .B(new_n432), .C1(new_n439), .C2(new_n407), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n407), .B1(new_n436), .B2(new_n438), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(G902), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n443), .A3(G475), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G952), .ZN(new_n446));
  AOI211_X1 g260(.A(G953), .B(new_n446), .C1(G234), .C2(G237), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT21), .B(G898), .Z(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT96), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI211_X1 g264(.A(new_n356), .B(new_n362), .C1(G234), .C2(G237), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n207), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n218), .B1(new_n232), .B2(new_n234), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n214), .A2(G143), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n218), .A2(G128), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n207), .B(new_n457), .C1(new_n307), .C2(new_n218), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G116), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT94), .B(G122), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n462), .B2(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(G107), .ZN(new_n465));
  INV_X1    g279(.A(G107), .ZN(new_n466));
  OAI221_X1 g280(.A(new_n461), .B1(KEYINPUT14), .B2(new_n466), .C1(new_n462), .C2(new_n460), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n457), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n471), .C1(new_n307), .C2(new_n218), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G134), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n463), .A2(new_n466), .ZN(new_n474));
  OAI211_X1 g288(.A(G107), .B(new_n461), .C1(new_n462), .C2(new_n460), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n458), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT9), .B(G234), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n478), .A2(new_n371), .A3(G953), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n468), .A2(new_n476), .A3(new_n479), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n362), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n484), .B(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT95), .Z(new_n488));
  NOR3_X1   g302(.A1(new_n445), .A2(new_n452), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G469), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n432), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n466), .A4(G104), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n394), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n394), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n498), .A2(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(KEYINPUT82), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(G101), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(G101), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n265), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT81), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT81), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n503), .A2(new_n507), .A3(KEYINPUT4), .A4(new_n504), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n502), .A2(new_n229), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n237), .A2(new_n214), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n240), .B1(new_n224), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n466), .A2(G104), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n394), .A2(G107), .ZN(new_n513));
  OAI21_X1  g327(.A(G101), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT10), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n240), .A2(new_n238), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n515), .A3(KEYINPUT10), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n509), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n210), .A2(new_n211), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n509), .A2(new_n522), .A3(new_n518), .A4(new_n520), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n356), .A2(G227), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n319), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT79), .B(G110), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n516), .B1(new_n519), .B2(new_n515), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n523), .A2(KEYINPUT12), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n211), .A3(new_n210), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n529), .B1(new_n537), .B2(new_n525), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n491), .B1(new_n539), .B2(G469), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n525), .A2(new_n529), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n533), .B2(new_n536), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n529), .B1(new_n524), .B2(new_n525), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n490), .B(new_n362), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT5), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n308), .A3(G116), .ZN(new_n547));
  OAI211_X1 g361(.A(G113), .B(new_n547), .C1(new_n249), .C2(new_n546), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n249), .A2(new_n250), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n515), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n506), .B(new_n508), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n555), .B2(new_n251), .ZN(new_n556));
  XOR2_X1   g370(.A(G110), .B(G122), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n502), .A2(new_n252), .A3(new_n506), .A4(new_n508), .ZN(new_n559));
  INV_X1    g373(.A(new_n557), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(KEYINPUT6), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n559), .B2(new_n552), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT84), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n558), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n561), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n240), .A2(new_n314), .A3(new_n238), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n229), .B2(new_n314), .ZN(new_n570));
  INV_X1    g384(.A(G224), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G953), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n570), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n577), .B2(new_n572), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n515), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n551), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n550), .A2(new_n581), .A3(new_n515), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n557), .B(KEYINPUT8), .Z(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n570), .B1(new_n576), .B2(new_n572), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n561), .A2(new_n580), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n575), .A2(new_n432), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT87), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n573), .B1(new_n566), .B2(new_n567), .ZN(new_n594));
  INV_X1    g408(.A(new_n588), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n594), .A2(G902), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n590), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G221), .B1(new_n478), .B2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(G214), .B1(G237), .B2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND4_X1   g417(.A1(new_n489), .A2(new_n545), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n302), .A2(KEYINPUT78), .A3(new_n375), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n378), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  AOI21_X1  g421(.A(G902), .B1(new_n568), .B2(new_n574), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n590), .B1(new_n608), .B2(new_n588), .ZN(new_n609));
  INV_X1    g423(.A(new_n590), .ZN(new_n610));
  NOR4_X1   g424(.A1(new_n594), .A2(G902), .A3(new_n610), .A4(new_n595), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n601), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n613));
  INV_X1    g427(.A(new_n452), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(new_n601), .C1(new_n609), .C2(new_n611), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n468), .A2(new_n476), .A3(new_n479), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n479), .B1(new_n468), .B2(new_n476), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT99), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n619), .A2(KEYINPUT99), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT33), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n295), .A2(new_n485), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT98), .B1(new_n483), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(KEYINPUT98), .B(new_n624), .C1(new_n618), .C2(new_n619), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n622), .B(new_n623), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n484), .A2(new_n485), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n624), .B1(new_n618), .B2(new_n619), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n626), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(KEYINPUT100), .A3(new_n623), .A4(new_n622), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n630), .A2(KEYINPUT101), .A3(new_n631), .A4(new_n636), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n445), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n617), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n289), .A2(new_n281), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n600), .B1(new_n540), .B2(new_n544), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n280), .B2(new_n295), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n375), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT34), .B(G104), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  INV_X1    g464(.A(new_n617), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n424), .B(new_n429), .C1(KEYINPUT20), .C2(new_n423), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n652), .A2(new_n444), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n488), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n651), .A2(new_n647), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT35), .B(G107), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT25), .B1(new_n368), .B2(new_n362), .ZN(new_n659));
  INV_X1    g473(.A(new_n360), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n352), .B2(new_n354), .ZN(new_n661));
  NOR4_X1   g475(.A1(new_n661), .A2(new_n366), .A3(new_n295), .A4(new_n363), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n373), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n355), .B(new_n664), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n374), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n646), .A2(new_n644), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n658), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n646), .A3(KEYINPUT102), .A4(new_n644), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n604), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AND3_X1   g488(.A1(new_n302), .A2(new_n645), .A3(new_n667), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n447), .B1(new_n451), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n653), .A2(new_n488), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n675), .A2(new_n616), .A3(new_n613), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XNOR2_X1  g496(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT104), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n598), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n593), .A2(new_n597), .A3(new_n684), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n645), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n677), .B(KEYINPUT39), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n601), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n445), .ZN(new_n694));
  INV_X1    g508(.A(new_n488), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n688), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n261), .A2(new_n270), .A3(new_n296), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n432), .B1(new_n287), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n283), .A2(new_n290), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n283), .A2(new_n290), .A3(new_n702), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n691), .A2(new_n692), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n696), .A2(new_n668), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  AND3_X1   g521(.A1(new_n641), .A2(new_n445), .A3(new_n678), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n613), .A2(new_n708), .A3(new_n616), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n613), .A2(new_n708), .A3(KEYINPUT106), .A4(new_n616), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n675), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  INV_X1    g528(.A(new_n376), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n362), .B1(new_n542), .B2(new_n543), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n717), .A2(new_n544), .A3(new_n599), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n617), .A2(new_n715), .A3(new_n642), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  AND3_X1   g535(.A1(new_n613), .A2(new_n616), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n368), .A2(new_n374), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n663), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n654), .A2(new_n724), .A3(new_n452), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n302), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND4_X1  g541(.A1(new_n722), .A2(new_n302), .A3(new_n489), .A4(new_n667), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n724), .A2(new_n452), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n285), .B(new_n732), .C1(new_n268), .C2(new_n297), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n287), .A2(new_n188), .B1(new_n297), .B2(new_n268), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n271), .B1(new_n734), .B2(KEYINPUT107), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n282), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(G472), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n289), .B2(new_n362), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n736), .A2(new_n694), .A3(new_n738), .A4(new_n695), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n722), .A2(new_n730), .A3(new_n731), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n613), .A2(new_n731), .A3(new_n616), .A4(new_n718), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n694), .A2(new_n695), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n733), .A2(new_n735), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n281), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n744), .A3(new_n646), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT108), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n646), .A3(new_n667), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n722), .A2(new_n708), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NAND2_X1  g566(.A1(new_n283), .A2(new_n290), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n283), .A2(KEYINPUT109), .B1(G472), .B2(new_n300), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n375), .A4(new_n708), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n611), .B1(new_n592), .B2(new_n589), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n601), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n689), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT109), .B1(new_n283), .B2(new_n290), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT32), .B1(new_n289), .B2(new_n281), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n301), .B1(new_n765), .B2(new_n754), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n375), .B(new_n708), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT42), .A4(new_n761), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n715), .A2(new_n708), .A3(new_n761), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n763), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  XNOR2_X1  g589(.A(new_n679), .B(KEYINPUT111), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n715), .A3(new_n761), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n531), .B2(new_n538), .ZN(new_n780));
  INV_X1    g594(.A(new_n521), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n781), .A2(new_n522), .B1(new_n533), .B2(new_n536), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n530), .B(KEYINPUT45), .C1(new_n782), .C2(new_n529), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(G469), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(KEYINPUT112), .A3(G469), .A4(new_n783), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n491), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(KEYINPUT46), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n544), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT46), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n599), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n690), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n639), .A2(new_n640), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT43), .B1(new_n795), .B2(new_n445), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n694), .A2(new_n797), .A3(new_n641), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n798), .A3(new_n669), .A4(new_n667), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n760), .B1(new_n799), .B2(new_n800), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  INV_X1    g619(.A(new_n708), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n793), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT47), .B(new_n599), .C1(new_n791), .C2(new_n792), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n302), .B(new_n806), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n760), .A2(new_n375), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n719), .A2(new_n747), .A3(new_n726), .A4(new_n728), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n647), .A2(new_n759), .A3(new_n602), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n445), .A2(KEYINPUT113), .A3(new_n487), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n445), .A2(new_n487), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n641), .B2(new_n445), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n614), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n302), .A2(new_n487), .A3(new_n653), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n642), .A2(new_n744), .A3(new_n646), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n760), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n689), .A2(new_n677), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n667), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n823), .A2(new_n829), .A3(new_n606), .A4(new_n672), .ZN(new_n830));
  INV_X1    g644(.A(new_n777), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n816), .A2(new_n832), .A3(new_n774), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n613), .A2(new_n742), .A3(new_n616), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n704), .A3(new_n668), .A4(new_n828), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n713), .A2(new_n835), .A3(new_n681), .A4(new_n751), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n815), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n836), .B(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n763), .A2(new_n770), .A3(new_n773), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n606), .A2(new_n672), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n777), .A3(new_n823), .A4(new_n829), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n844), .A3(KEYINPUT53), .A4(new_n816), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT54), .B1(new_n838), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n796), .A2(new_n798), .A3(new_n447), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n593), .A2(new_n718), .A3(new_n597), .A4(new_n601), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n750), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n796), .A3(new_n798), .A4(new_n447), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT116), .B1(new_n853), .B2(new_n749), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n375), .A2(new_n447), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n703), .A2(new_n701), .A3(new_n855), .A4(new_n851), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n641), .A2(new_n445), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n852), .A2(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT117), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n686), .A2(new_n687), .A3(new_n718), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n744), .A2(new_n375), .A3(new_n646), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n849), .A2(new_n860), .A3(new_n602), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n796), .A2(new_n798), .A3(new_n447), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n861), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(KEYINPUT50), .A3(new_n602), .A4(new_n860), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n717), .A2(new_n544), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n600), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n808), .A2(new_n809), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n827), .A3(new_n867), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(KEYINPUT51), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n446), .A2(G953), .ZN(new_n877));
  XNOR2_X1  g691(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n865), .A2(new_n868), .A3(KEYINPUT115), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n874), .A2(new_n879), .A3(new_n858), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT115), .B1(new_n865), .B2(new_n868), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n876), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n724), .B(new_n853), .C1(new_n755), .C2(new_n756), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT48), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n856), .A2(new_n642), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n867), .A2(new_n722), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n883), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n814), .B1(new_n848), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n446), .A2(new_n356), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n876), .A2(new_n882), .A3(new_n877), .A4(new_n888), .ZN(new_n892));
  INV_X1    g706(.A(new_n887), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n885), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(KEYINPUT118), .C1(new_n847), .C2(new_n846), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT49), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n704), .B1(new_n897), .B2(new_n871), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n445), .B(new_n795), .C1(KEYINPUT49), .C2(new_n870), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n688), .A2(new_n375), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n603), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(G75));
  XNOR2_X1  g716(.A(new_n568), .B(new_n574), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n362), .B1(new_n838), .B2(new_n845), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n610), .ZN(new_n908));
  OAI211_X1 g722(.A(KEYINPUT120), .B(new_n906), .C1(new_n908), .C2(KEYINPUT56), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n356), .A2(G952), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n907), .B2(new_n592), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n905), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT56), .B1(new_n907), .B2(new_n610), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n905), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(G51));
  OR2_X1    g730(.A1(new_n789), .A2(KEYINPUT57), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n789), .A2(KEYINPUT57), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n848), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n542), .A2(new_n543), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n907), .A2(new_n786), .A3(new_n787), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n910), .B1(new_n921), .B2(new_n922), .ZN(G54));
  NAND3_X1  g737(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n924));
  INV_X1    g738(.A(new_n421), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n910), .ZN(G60));
  INV_X1    g742(.A(new_n847), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n838), .A2(new_n845), .A3(KEYINPUT54), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n635), .A2(new_n622), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n910), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n838), .B2(new_n845), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(new_n368), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n910), .B1(new_n940), .B2(new_n665), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(KEYINPUT61), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(G66));
  NAND3_X1  g761(.A1(new_n816), .A2(new_n842), .A3(new_n823), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n356), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n450), .B2(new_n571), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT122), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n566), .B(new_n567), .C1(G898), .C2(new_n356), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(new_n955), .Z(G69));
  AND2_X1   g770(.A1(new_n713), .A2(new_n681), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n706), .A2(new_n751), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n822), .A2(KEYINPUT124), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n961), .A2(new_n378), .A3(new_n605), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n762), .A2(new_n690), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n962), .B(new_n963), .C1(KEYINPUT124), .C2(new_n822), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n810), .A2(new_n811), .B1(new_n802), .B2(new_n803), .ZN(new_n965));
  XNOR2_X1  g779(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n958), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n960), .A2(new_n964), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n356), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n248), .A2(new_n255), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n413), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n356), .B1(G227), .B2(G900), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n676), .B2(G227), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n794), .A2(new_n375), .A3(new_n757), .A4(new_n834), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n957), .A2(new_n976), .A3(new_n751), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n965), .A2(new_n977), .A3(new_n774), .A4(new_n777), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n971), .B(new_n975), .C1(new_n978), .C2(G953), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT125), .ZN(G72));
  XNOR2_X1  g795(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n968), .B2(new_n948), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n268), .A3(new_n284), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n838), .A2(new_n845), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n293), .B1(new_n284), .B2(new_n270), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n984), .B1(new_n978), .B2(new_n948), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n284), .A2(new_n268), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n910), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n986), .B(new_n989), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(G57));
endmodule


