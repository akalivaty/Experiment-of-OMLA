//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n213), .B(new_n214), .C1(new_n201), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G58), .C2(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT0), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n219), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n226), .A2(new_n227), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n228), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT64), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n222), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n211), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G226), .B(G232), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G358));
  NAND2_X1  g0049(.A1(G68), .A2(G77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT67), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(G107), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(new_n210), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  NAND3_X1  g0058(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n233), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n218), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n268));
  INV_X1    g0068(.A(G150), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n219), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n219), .A2(G33), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n268), .B1(new_n269), .B2(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n260), .B(new_n267), .C1(new_n279), .C2(new_n262), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(KEYINPUT9), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G223), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n284), .B1(new_n202), .B2(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n288), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(G226), .A3(new_n290), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n280), .A2(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(G200), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n281), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(new_n281), .A4(new_n298), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n280), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT70), .B(G179), .Z(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n296), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n296), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  OAI211_X1 g0116(.A(G226), .B(new_n283), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(G232), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n292), .B1(new_n320), .B2(new_n288), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n294), .A2(G238), .A3(new_n290), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n325));
  OAI21_X1  g0125(.A(G169), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(G169), .C1(new_n324), .C2(new_n325), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n321), .A2(KEYINPUT72), .A3(new_n323), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n321), .A2(KEYINPUT72), .A3(new_n323), .A4(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n331), .A2(new_n334), .A3(G179), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n327), .A2(new_n329), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n201), .A2(G20), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n339), .B1(new_n202), .B2(new_n278), .C1(new_n275), .C2(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n262), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n259), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n201), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(KEYINPUT11), .A3(new_n262), .ZN(new_n347));
  INV_X1    g0147(.A(new_n265), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G68), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n343), .A2(new_n346), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n338), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n350), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n331), .A2(new_n334), .A3(G190), .A4(new_n336), .ZN(new_n353));
  OAI21_X1  g0153(.A(G200), .B1(new_n324), .B2(new_n325), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n276), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n274), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT15), .B(G87), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n357), .B1(new_n219), .B2(new_n202), .C1(new_n278), .C2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n262), .B1(new_n202), .B2(new_n344), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n348), .A2(G77), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n364), .B1(new_n206), .B2(new_n282), .C1(new_n285), .C2(new_n215), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n288), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n294), .A2(G244), .A3(new_n290), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n293), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n363), .B1(G200), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n366), .A2(new_n293), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G190), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n351), .A2(new_n355), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(G226), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n374));
  OAI211_X1 g0174(.A(G223), .B(new_n283), .C1(new_n315), .C2(new_n316), .ZN(new_n375));
  INV_X1    g0175(.A(G87), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n271), .A2(new_n376), .A3(KEYINPUT75), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT75), .B1(new_n271), .B2(new_n376), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n374), .A2(new_n375), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n288), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n294), .A2(G232), .A3(new_n290), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n293), .A3(new_n381), .A4(new_n308), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n293), .A3(new_n381), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n311), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n292), .B1(new_n379), .B2(new_n288), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n381), .A4(new_n308), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n315), .A2(new_n316), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(new_n219), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR4_X1   g0192(.A1(new_n315), .A2(new_n316), .A3(new_n392), .A4(G20), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n274), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n230), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT73), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G159), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n272), .B2(new_n273), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n219), .B1(new_n230), .B2(new_n396), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n394), .B(KEYINPUT16), .C1(new_n399), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n392), .B1(new_n282), .B2(G20), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n201), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n395), .A2(new_n398), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n262), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT68), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n276), .B(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n259), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n348), .B2(new_n415), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n412), .B2(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n389), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n384), .A2(G200), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT77), .B(G190), .Z(new_n423));
  NAND3_X1  g0223(.A1(new_n386), .A2(new_n381), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n412), .A2(new_n417), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT17), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n389), .C1(new_n418), .C2(new_n419), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n370), .A2(new_n308), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n368), .A2(new_n311), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n363), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n314), .A2(new_n373), .A3(new_n429), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(KEYINPUT6), .A2(G97), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT78), .B1(new_n435), .B2(G107), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT78), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(new_n206), .A3(KEYINPUT6), .A4(G97), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT6), .ZN(new_n440));
  XNOR2_X1  g0240(.A(G97), .B(G107), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n442), .A2(new_n219), .B1(new_n202), .B2(new_n275), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n206), .B1(new_n407), .B2(new_n408), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n262), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n259), .A2(G97), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n218), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n259), .A2(new_n448), .A3(new_n233), .A4(new_n261), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n205), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n445), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(G244), .B(new_n283), .C1(new_n315), .C2(new_n316), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n453), .A2(new_n454), .B1(G33), .B2(G283), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n458), .A4(new_n456), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n288), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT5), .B(G41), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n218), .A2(G45), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n465), .A2(G274), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n288), .B1(new_n467), .B2(new_n465), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(G257), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n464), .A2(G190), .A3(new_n470), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n452), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n311), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n464), .A2(new_n308), .A3(new_n470), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n445), .A2(new_n447), .A3(new_n451), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G257), .B(new_n283), .C1(new_n315), .C2(new_n316), .ZN(new_n480));
  INV_X1    g0280(.A(new_n316), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT3), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(G303), .A3(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G264), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n468), .B1(new_n485), .B2(new_n288), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n469), .A2(G270), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n486), .A2(KEYINPUT80), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT80), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g0289(.A(G200), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n288), .ZN(new_n491));
  INV_X1    g0291(.A(new_n468), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(KEYINPUT80), .A3(new_n487), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n423), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n457), .B(new_n219), .C1(G33), .C2(new_n205), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n210), .A2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n262), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n262), .A4(new_n499), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(new_n210), .B2(new_n344), .ZN(new_n504));
  INV_X1    g0304(.A(new_n449), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n490), .A2(new_n497), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n311), .B1(new_n504), .B2(new_n506), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n488), .B2(new_n489), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n486), .A2(G179), .A3(new_n487), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n495), .A2(new_n496), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT21), .A3(new_n510), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n509), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n479), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G257), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n520));
  OAI211_X1 g0320(.A(G250), .B(new_n283), .C1(new_n315), .C2(new_n316), .ZN(new_n521));
  OR2_X1    g0321(.A1(KEYINPUT81), .A2(G294), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT81), .A2(G294), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G33), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT82), .A4(new_n524), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n288), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n469), .A2(G264), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n297), .A4(new_n492), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n492), .A3(new_n530), .ZN(new_n534));
  INV_X1    g0334(.A(G200), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT83), .B1(new_n534), .B2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n219), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n282), .A2(new_n542), .A3(new_n219), .A4(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(G20), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n219), .A2(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT23), .ZN(new_n549));
  AND4_X1   g0349(.A1(new_n539), .A2(new_n544), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n546), .B1(new_n541), .B2(new_n543), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n539), .B1(new_n551), .B2(new_n549), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n262), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n449), .A2(new_n206), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n259), .A2(G107), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n556), .B(KEYINPUT25), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n538), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n534), .A2(new_n311), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n534), .A2(G179), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G41), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n271), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G250), .B(new_n466), .C1(new_n565), .C2(new_n233), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n467), .A2(G274), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G244), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n569));
  OAI211_X1 g0369(.A(G238), .B(new_n283), .C1(new_n315), .C2(new_n316), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n545), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n288), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G190), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n219), .B1(new_n319), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n376), .A2(new_n205), .A3(new_n206), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n219), .A2(G33), .A3(G97), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n219), .B(G68), .C1(new_n315), .C2(new_n316), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n263), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n449), .A2(new_n376), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n358), .A2(new_n259), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n573), .B(new_n583), .C1(new_n535), .C2(new_n572), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n572), .A2(new_n308), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n575), .A2(new_n576), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n577), .A2(new_n574), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n579), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n262), .ZN(new_n589));
  INV_X1    g0389(.A(new_n582), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n359), .C2(new_n449), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n585), .B(new_n591), .C1(G169), .C2(new_n572), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n563), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n434), .A2(new_n519), .A3(new_n560), .A4(new_n594), .ZN(new_n595));
  XOR2_X1   g0395(.A(new_n595), .B(KEYINPUT84), .Z(G372));
  INV_X1    g0396(.A(new_n313), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n370), .A2(new_n308), .B1(new_n361), .B2(new_n362), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n598), .A2(KEYINPUT87), .A3(new_n431), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT87), .B1(new_n598), .B2(new_n431), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n355), .B1(new_n350), .B2(new_n338), .ZN(new_n602));
  INV_X1    g0402(.A(new_n426), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n412), .A2(new_n417), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT18), .B1(new_n389), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n412), .A2(new_n417), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n606), .A2(new_n427), .A3(new_n607), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n602), .A2(new_n603), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n597), .B1(new_n609), .B2(new_n306), .ZN(new_n610));
  INV_X1    g0410(.A(new_n434), .ZN(new_n611));
  INV_X1    g0411(.A(new_n592), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n593), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(KEYINPUT26), .ZN(new_n614));
  INV_X1    g0414(.A(new_n478), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n583), .B(KEYINPUT85), .C1(new_n535), .C2(new_n572), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n571), .A2(new_n288), .ZN(new_n619));
  INV_X1    g0419(.A(new_n568), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n535), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n581), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n589), .A2(new_n622), .A3(new_n590), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n618), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n617), .A2(new_n624), .A3(new_n573), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n625), .A2(KEYINPUT86), .A3(new_n592), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT86), .B1(new_n625), .B2(new_n592), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n615), .B(new_n616), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n478), .B(new_n474), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n560), .B1(new_n626), .B2(new_n627), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n614), .B(new_n628), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n610), .B1(new_n611), .B2(new_n634), .ZN(G369));
  NOR2_X1   g0435(.A1(new_n223), .A2(G20), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT27), .B1(new_n637), .B2(G1), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT27), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n639), .A3(new_n218), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n638), .A2(G213), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G343), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT88), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n558), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n560), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n563), .ZN(new_n646));
  INV_X1    g0446(.A(new_n643), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n629), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT90), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n647), .A2(new_n508), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n518), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n630), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT89), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT89), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n650), .B1(new_n658), .B2(G330), .ZN(new_n659));
  INV_X1    g0459(.A(G330), .ZN(new_n660));
  AOI211_X1 g0460(.A(KEYINPUT90), .B(new_n660), .C1(new_n655), .C2(new_n657), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n649), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n630), .A2(new_n647), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n646), .A2(new_n648), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n648), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(G399));
  NOR2_X1   g0466(.A1(new_n224), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n576), .A2(G116), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n231), .B2(new_n668), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  INV_X1    g0472(.A(new_n627), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n625), .A2(KEYINPUT86), .A3(new_n592), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n563), .A2(new_n515), .A3(new_n517), .A4(new_n513), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n474), .A2(new_n478), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n560), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n615), .B1(new_n626), .B2(new_n627), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n615), .A2(new_n616), .A3(new_n593), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n678), .A2(new_n680), .A3(new_n592), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .A3(new_n647), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n633), .A2(new_n647), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n682), .A2(KEYINPUT92), .A3(KEYINPUT29), .A4(new_n647), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n471), .A2(new_n534), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n309), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n572), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n471), .A2(KEYINPUT91), .A3(new_n534), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n693), .A2(new_n516), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n471), .A2(new_n514), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n529), .A2(new_n530), .A3(new_n572), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT30), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n471), .A2(new_n701), .A3(new_n698), .A4(new_n514), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n647), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n519), .A2(new_n560), .A3(new_n594), .A4(new_n647), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n696), .A2(new_n703), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n690), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n672), .B1(new_n713), .B2(G1), .ZN(G364));
  NAND2_X1  g0514(.A1(new_n658), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT90), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n658), .A2(new_n650), .A3(G330), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n218), .B1(new_n636), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI221_X1 g0521(.A(new_n719), .B1(G330), .B2(new_n658), .C1(new_n667), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n233), .B1(G20), .B2(new_n311), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n219), .A2(G179), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n297), .A3(G200), .ZN(new_n725));
  INV_X1    g0525(.A(G283), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n308), .A2(new_n219), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G200), .ZN(new_n729));
  INV_X1    g0529(.A(new_n423), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n731), .A2(G326), .B1(new_n734), .B2(G311), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n724), .A2(G190), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(G303), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n390), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n219), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n522), .A2(new_n523), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n724), .A2(new_n732), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n738), .B(new_n742), .C1(G329), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n309), .A2(G20), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(G200), .A3(new_n730), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n735), .B(new_n745), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n729), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT96), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n729), .A2(new_n753), .A3(G190), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n727), .B(new_n750), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(new_n201), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n749), .A2(new_n229), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT95), .B(G159), .Z(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n744), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n736), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(G87), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n725), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G107), .ZN(new_n767));
  INV_X1    g0567(.A(new_n740), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n390), .B1(new_n768), .B2(G97), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n744), .A2(new_n761), .A3(new_n762), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n765), .A2(new_n767), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n731), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n772), .A2(new_n266), .B1(new_n733), .B2(new_n202), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n759), .A2(new_n760), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n723), .B1(new_n758), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n667), .A2(new_n721), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n224), .A2(new_n282), .ZN(new_n778));
  INV_X1    g0578(.A(G45), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n232), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(new_n254), .C2(new_n779), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n225), .A2(G355), .A3(new_n282), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n781), .B(new_n782), .C1(G116), .C2(new_n225), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n723), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n777), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT94), .Z(new_n789));
  INV_X1    g0589(.A(new_n786), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n775), .B(new_n789), .C1(new_n658), .C2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n722), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  AND2_X1   g0593(.A1(new_n643), .A2(new_n363), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n369), .B2(new_n371), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n432), .A2(KEYINPUT99), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n432), .A2(KEYINPUT99), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n794), .B1(new_n599), .B2(new_n600), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n686), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n633), .A2(new_n647), .A3(new_n800), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n711), .B(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(new_n776), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n734), .A2(new_n762), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G137), .A2(new_n731), .B1(new_n748), .B2(G143), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n755), .C2(new_n269), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT34), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n764), .A2(G50), .B1(new_n766), .B2(G68), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n282), .B1(new_n229), .B2(new_n740), .C1(new_n813), .C2(KEYINPUT98), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(KEYINPUT98), .B2(new_n813), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n811), .B(new_n816), .C1(G132), .C2(new_n744), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n390), .B1(new_n743), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n766), .A2(G87), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n820), .B1(new_n206), .B2(new_n736), .C1(new_n205), .C2(new_n740), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G116), .C2(new_n734), .ZN(new_n822));
  INV_X1    g0622(.A(G294), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n823), .B2(new_n749), .C1(new_n755), .C2(new_n726), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G303), .B2(new_n731), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n723), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n777), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n723), .A2(new_n784), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(G77), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n826), .B(new_n831), .C1(new_n785), .C2(new_n800), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n806), .A2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(KEYINPUT40), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n351), .A2(new_n835), .A3(new_n355), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n350), .A2(new_n643), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n338), .A2(new_n837), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n839), .A2(new_n351), .A3(new_n835), .A4(new_n355), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n709), .A2(new_n707), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n800), .C1(new_n842), .C2(new_n705), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  INV_X1    g0644(.A(new_n641), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n394), .B1(new_n399), .B2(new_n404), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n406), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n262), .A3(new_n405), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n607), .A2(new_n845), .B1(new_n848), .B2(new_n417), .ZN(new_n849));
  AND4_X1   g0649(.A1(new_n412), .A2(new_n417), .A3(new_n422), .A4(new_n424), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n418), .A2(new_n419), .B1(new_n389), .B2(new_n641), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n425), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n845), .B1(new_n848), .B2(new_n417), .ZN(new_n857));
  AOI221_X4 g0657(.A(new_n844), .B1(new_n851), .B2(new_n856), .C1(new_n429), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n429), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n851), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n834), .B1(new_n843), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n860), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n604), .A2(KEYINPUT74), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n866), .A2(new_n867), .B1(new_n607), .B2(new_n845), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n868), .B2(new_n854), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n845), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n425), .B1(new_n606), .B2(new_n607), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n852), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n608), .A2(new_n605), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n870), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n864), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n838), .A2(new_n840), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n801), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n880), .A2(new_n710), .A3(KEYINPUT40), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n863), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n434), .A2(new_n710), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n885), .B(new_n886), .Z(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(G330), .ZN(new_n888));
  OR3_X1    g0688(.A1(new_n608), .A2(new_n605), .A3(new_n641), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n796), .A2(new_n797), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n643), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n803), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n841), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n859), .A2(new_n860), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n844), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n895), .B1(new_n897), .B2(new_n864), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n874), .B2(new_n878), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n858), .A2(new_n899), .A3(KEYINPUT39), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n351), .A2(new_n643), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI221_X1 g0703(.A(new_n889), .B1(new_n862), .B2(new_n894), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n685), .A2(new_n434), .A3(new_n688), .A4(new_n689), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n610), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n904), .B(new_n906), .Z(new_n907));
  XNOR2_X1  g0707(.A(new_n888), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n218), .B2(new_n636), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT35), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n219), .B(new_n233), .C1(new_n442), .C2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(G116), .C1(new_n910), .C2(new_n442), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n396), .A2(G77), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n231), .A2(new_n914), .B1(G50), .B2(new_n201), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(G1), .A3(new_n223), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n913), .A3(new_n916), .ZN(G367));
  OAI22_X1  g0717(.A1(new_n749), .A2(new_n737), .B1(new_n726), .B2(new_n733), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n282), .B1(new_n744), .B2(G317), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n766), .A2(G97), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(new_n206), .C2(new_n740), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n736), .A2(new_n210), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT46), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n918), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n924), .B1(new_n818), .B2(new_n772), .C1(new_n741), .C2(new_n755), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n768), .A2(G68), .B1(new_n764), .B2(G58), .ZN(new_n926));
  INV_X1    g0726(.A(G137), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n926), .B1(new_n202), .B2(new_n725), .C1(new_n927), .C2(new_n743), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n390), .B(new_n928), .C1(G143), .C2(new_n731), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n756), .A2(new_n762), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(new_n266), .C2(new_n733), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n749), .A2(new_n269), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n777), .B1(new_n934), .B2(new_n723), .ZN(new_n935));
  INV_X1    g0735(.A(new_n778), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n787), .B1(new_n225), .B2(new_n359), .C1(new_n243), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n647), .A2(new_n583), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n673), .B2(new_n674), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT103), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n612), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n940), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n935), .B(new_n937), .C1(new_n790), .C2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n677), .B1(new_n452), .B2(new_n647), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n615), .A2(new_n643), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT105), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n478), .B1(new_n951), .B2(new_n563), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n647), .ZN(new_n953));
  INV_X1    g0753(.A(new_n950), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n664), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT42), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n947), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n947), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n662), .A2(new_n951), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n649), .A2(new_n663), .ZN(new_n965));
  INV_X1    g0765(.A(new_n664), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT106), .B1(new_n716), .B2(new_n717), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT106), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n659), .A2(new_n661), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n718), .A2(new_n969), .ZN(new_n972));
  INV_X1    g0772(.A(new_n967), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n974), .A3(new_n713), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n665), .B2(new_n950), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n664), .A2(new_n648), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n665), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n978), .B2(new_n954), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n977), .A2(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n662), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n662), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n713), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n667), .B(KEYINPUT41), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n721), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n945), .B1(new_n964), .B2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n356), .A2(new_n266), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n992));
  INV_X1    g0792(.A(new_n669), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n994));
  AND4_X1   g0794(.A1(new_n779), .A2(new_n992), .A3(new_n994), .A4(new_n250), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n778), .B1(new_n248), .B2(new_n779), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n225), .A3(new_n282), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n225), .A2(G107), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n787), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G322), .A2(new_n731), .B1(new_n748), .B2(G317), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n737), .B2(new_n733), .C1(new_n755), .C2(new_n818), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT48), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n726), .B2(new_n740), .C1(new_n741), .C2(new_n736), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n744), .A2(G326), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n282), .B1(new_n766), .B2(G116), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n749), .A2(new_n266), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n768), .A2(new_n358), .B1(new_n764), .B2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n269), .B2(new_n743), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n733), .A2(new_n201), .ZN(new_n1014));
  NOR4_X1   g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n390), .A4(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT107), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n772), .B2(new_n400), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n731), .A2(KEYINPUT107), .A3(G159), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n1017), .A2(new_n920), .A3(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1015), .B(new_n1019), .C1(new_n277), .C2(new_n755), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1010), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n723), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n827), .B(new_n1000), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT108), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n649), .A2(new_n790), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(KEYINPUT108), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n716), .A2(KEYINPUT106), .A3(new_n717), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n973), .B1(new_n972), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n968), .A2(new_n967), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n712), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n667), .A3(new_n975), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n721), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1027), .A2(new_n1032), .A3(new_n1034), .ZN(G393));
  NAND3_X1  g0835(.A1(new_n984), .A2(new_n721), .A3(new_n985), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G150), .A2(new_n731), .B1(new_n748), .B2(G159), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT51), .Z(new_n1038));
  AOI22_X1  g0838(.A1(new_n768), .A2(G77), .B1(new_n764), .B2(G68), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n744), .A2(G143), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n276), .C2(new_n733), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n756), .B2(G50), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1042), .A3(new_n282), .A4(new_n820), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G317), .A2(new_n731), .B1(new_n748), .B2(G311), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n282), .B1(new_n768), .B2(G116), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n736), .A2(new_n726), .B1(new_n743), .B2(new_n746), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n767), .C1(KEYINPUT109), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(KEYINPUT109), .B2(new_n1047), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1045), .B(new_n1049), .C1(new_n737), .C2(new_n755), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n733), .A2(new_n823), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n723), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n787), .B1(new_n205), .B2(new_n225), .C1(new_n257), .C2(new_n936), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n827), .A3(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT110), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n951), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n790), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1036), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT111), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1036), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n668), .B1(new_n975), .B2(new_n986), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n986), .B2(new_n975), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(G390));
  NAND3_X1  g0866(.A1(new_n710), .A2(G330), .A3(new_n882), .ZN(new_n1067));
  OAI211_X1 g0867(.A(G330), .B(new_n800), .C1(new_n842), .C2(new_n705), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n881), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n893), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n682), .A2(new_n647), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n891), .B1(new_n1072), .B2(new_n800), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n434), .A2(new_n710), .A3(G330), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n905), .A2(new_n610), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT112), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n894), .A2(new_n1080), .A3(new_n903), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n881), .B1(new_n803), .B2(new_n892), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT112), .B1(new_n1082), .B2(new_n902), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n901), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n903), .B(new_n880), .C1(new_n1073), .C2(new_n881), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n1067), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1067), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1079), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1067), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1084), .A2(new_n1085), .A3(new_n1067), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1077), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1088), .A2(new_n1094), .A3(new_n667), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT113), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1088), .A2(new_n1094), .A3(KEYINPUT113), .A4(new_n667), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n755), .A2(new_n206), .B1(new_n205), .B2(new_n733), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT117), .Z(new_n1101));
  AOI22_X1  g0901(.A1(new_n768), .A2(G77), .B1(new_n766), .B2(G68), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n376), .B2(new_n736), .C1(new_n749), .C2(new_n210), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n390), .B1(new_n823), .B2(new_n743), .C1(new_n772), .C2(new_n726), .ZN(new_n1104));
  OR3_X1    g0904(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  AOI22_X1  g0906(.A1(new_n756), .A2(G137), .B1(new_n734), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT115), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n731), .A2(G128), .B1(G132), .B2(new_n748), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n282), .B1(new_n725), .B2(new_n266), .C1(new_n740), .C2(new_n400), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G125), .B2(new_n744), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n736), .A2(new_n269), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1022), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n827), .B1(new_n415), .B2(new_n829), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT114), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(new_n901), .C2(new_n784), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n721), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1099), .A2(new_n1121), .ZN(G378));
  INV_X1    g0922(.A(KEYINPUT57), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1077), .B1(new_n1120), .B2(new_n1075), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n863), .A2(G330), .A3(new_n883), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT55), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n306), .B2(new_n313), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n306), .A2(new_n1127), .A3(new_n313), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(new_n280), .C2(new_n845), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n280), .A2(new_n845), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1130), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n1128), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1126), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT39), .B1(new_n858), .B2(new_n861), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n880), .B2(KEYINPUT39), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n862), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(new_n902), .B1(new_n1144), .B2(new_n1082), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT122), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n863), .A2(new_n883), .A3(new_n1146), .A4(G330), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1147), .A3(new_n889), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n889), .B2(new_n1145), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1141), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1147), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n904), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1145), .A2(new_n1147), .A3(new_n889), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n1126), .A4(new_n1140), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1123), .B1(new_n1124), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1094), .A2(new_n1078), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1157), .A2(KEYINPUT57), .A3(new_n1154), .A4(new_n1150), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n667), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1155), .A2(new_n720), .ZN(new_n1160));
  INV_X1    g0960(.A(G132), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n755), .A2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G125), .A2(new_n731), .B1(new_n748), .B2(G128), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n927), .B2(new_n733), .C1(new_n269), .C2(new_n740), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(new_n764), .C2(new_n1106), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT59), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G41), .B1(new_n766), .B2(new_n762), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G33), .B1(new_n744), .B2(G124), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n755), .A2(new_n205), .B1(new_n359), .B2(new_n733), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT119), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n768), .A2(G68), .B1(G283), .B2(new_n744), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G116), .A2(new_n731), .B1(new_n748), .B2(G107), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G41), .B(new_n282), .C1(new_n764), .C2(G77), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT118), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n766), .A2(G58), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1171), .B(new_n1178), .C1(KEYINPUT118), .C2(new_n1175), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT58), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n266), .B1(new_n315), .B2(G41), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1169), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1184), .A2(new_n723), .B1(new_n266), .B2(new_n828), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n776), .B(new_n1185), .C1(new_n1140), .C2(new_n785), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT121), .Z(new_n1187));
  NOR2_X1   g0987(.A1(new_n1160), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1159), .A2(new_n1188), .ZN(G375));
  NOR2_X1   g0989(.A1(new_n755), .A2(new_n210), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n359), .A2(new_n740), .B1(new_n205), .B2(new_n736), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n390), .B1(new_n737), .B2(new_n743), .C1(new_n733), .C2(new_n206), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G77), .C2(new_n766), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n726), .B2(new_n749), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1190), .B(new_n1194), .C1(G294), .C2(new_n731), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n748), .A2(G137), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n744), .A2(G128), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n768), .A2(G50), .B1(new_n764), .B2(G159), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1196), .A2(new_n282), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1177), .B1(new_n269), .B2(new_n733), .C1(new_n772), .C2(new_n1161), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n756), .C2(new_n1106), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n723), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n827), .B(new_n1202), .C1(new_n841), .C2(new_n785), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n201), .B2(new_n828), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1075), .B2(new_n721), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1071), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n988), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1207), .B2(new_n1093), .ZN(G381));
  AND2_X1   g1008(.A1(new_n1095), .A2(new_n1121), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1159), .A2(new_n1188), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G384), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1027), .A2(new_n1032), .A3(new_n792), .A4(new_n1034), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G387), .A2(G381), .A3(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1214), .ZN(G407));
  INV_X1    g1015(.A(G213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(G343), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1210), .A2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT123), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1020(.A1(G387), .A2(new_n1212), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n662), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(new_n983), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n712), .B1(new_n1033), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n988), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n720), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n961), .B(new_n962), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(G390), .A3(new_n945), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1213), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1221), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1221), .A2(new_n1229), .A3(new_n1231), .A4(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1229), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1228), .A2(G390), .A3(KEYINPUT125), .A4(new_n945), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1221), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1231), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G378), .A2(new_n1159), .A3(new_n1188), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1124), .A2(new_n1155), .A3(new_n1225), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1186), .B1(new_n1155), .B2(new_n720), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1209), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1217), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n668), .B1(new_n1206), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1079), .C1(new_n1249), .C2(new_n1206), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G384), .A3(new_n1205), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1251), .B2(new_n1205), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1217), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1217), .A2(G2897), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT124), .Z(new_n1262));
  OR3_X1    g1062(.A1(new_n1253), .A2(new_n1254), .A3(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1257), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1255), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1260), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1243), .B(new_n1256), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1248), .A2(new_n1271), .A3(new_n1255), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1248), .B2(new_n1265), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1248), .B2(new_n1255), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1270), .B1(new_n1276), .B2(new_n1277), .ZN(G405));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G375), .A2(new_n1209), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1255), .A2(KEYINPUT127), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1244), .A4(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1281), .A2(new_n1244), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1277), .ZN(G402));
endmodule


