//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT68), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  NAND2_X1  g011(.A1(G113gat), .A2(G120gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n208), .B(new_n214), .C1(KEYINPUT68), .C2(new_n205), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  AND2_X1   g015(.A1(G113gat), .A2(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G113gat), .A2(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n211), .A2(KEYINPUT69), .A3(new_n213), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n212), .A4(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n224));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT77), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G155gat), .A3(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G155gat), .ZN(new_n230));
  INV_X1    g029(.A(G162gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G141gat), .B(G148gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n229), .B(new_n232), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G148gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT78), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G148gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n241), .A3(G141gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(G141gat), .B2(new_n238), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT80), .B1(new_n225), .B2(KEYINPUT2), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n225), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248));
  NOR2_X1   g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n248), .B1(new_n233), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n232), .A2(KEYINPUT79), .A3(new_n225), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n243), .A2(new_n247), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n223), .A2(new_n224), .A3(new_n237), .A4(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n225), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n250), .B(new_n251), .C1(new_n254), .C2(new_n244), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n238), .A2(G141gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT78), .B(G148gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(G141gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n237), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n215), .A2(new_n222), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n237), .C1(new_n255), .C2(new_n258), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  AOI211_X1 g065(.A(KEYINPUT39), .B(new_n203), .C1(new_n262), .C2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n202), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n266), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT39), .ZN(new_n274));
  INV_X1    g073(.A(new_n203), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT84), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n275), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n252), .A2(new_n215), .A3(new_n222), .A4(new_n237), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n260), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(new_n275), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(new_n274), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n272), .A2(new_n278), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT85), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT40), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n279), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n267), .A2(new_n202), .A3(new_n271), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT84), .B1(new_n276), .B2(new_n277), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT40), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT85), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(KEYINPUT40), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n282), .B2(new_n275), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(KEYINPUT4), .C1(new_n259), .C2(new_n260), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n266), .A2(new_n299), .A3(new_n203), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n253), .A2(new_n261), .A3(KEYINPUT81), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n262), .A2(new_n296), .A3(new_n203), .A4(new_n266), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n304), .A2(KEYINPUT86), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n277), .B1(new_n304), .B2(KEYINPUT86), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(G218gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n310), .B(new_n311), .C1(new_n317), .C2(KEYINPUT22), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n321));
  OAI21_X1  g120(.A(G218gat), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n311), .B1(new_n324), .B2(new_n310), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n309), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n311), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT73), .B(G211gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT22), .B1(new_n328), .B2(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n310), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(KEYINPUT74), .A3(new_n318), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT23), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT24), .B1(new_n343), .B2(G183gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n342), .A2(G190gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT65), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(G169gat), .A3(G176gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n336), .A2(KEYINPUT23), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n340), .A2(new_n347), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n352), .A2(new_n355), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(new_n357), .A3(new_n340), .A4(new_n347), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n336), .A2(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(KEYINPUT26), .A2(new_n365), .B1(new_n349), .B2(new_n351), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n365), .A2(KEYINPUT26), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n366), .A2(new_n367), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n342), .A2(KEYINPUT27), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G183gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n371), .A3(new_n343), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n362), .A2(new_n363), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n362), .B2(new_n375), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n334), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n375), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n319), .A2(new_n325), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n359), .A2(new_n361), .B1(new_n368), .B2(new_n374), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n377), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  AOI21_X1  g186(.A(new_n308), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  AOI211_X1 g188(.A(KEYINPUT76), .B(new_n389), .C1(new_n379), .C2(new_n383), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n388), .A2(new_n390), .A3(KEYINPUT30), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n387), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n387), .B2(new_n384), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n295), .B(new_n307), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT87), .B1(new_n294), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n286), .B1(new_n285), .B2(KEYINPUT40), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n291), .A2(KEYINPUT85), .A3(new_n292), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n393), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n387), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT76), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n308), .A3(new_n387), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n399), .A2(new_n404), .B1(new_n305), .B2(new_n306), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n398), .A2(new_n405), .A3(new_n406), .A4(new_n295), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n376), .A2(new_n378), .B1(new_n319), .B2(new_n325), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n380), .B(new_n333), .C1(new_n382), .C2(new_n377), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT37), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n408), .A2(KEYINPUT88), .A3(KEYINPUT37), .A4(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT37), .B1(new_n379), .B2(new_n383), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n415), .A2(KEYINPUT38), .A3(new_n387), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n384), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n379), .A2(KEYINPUT37), .A3(new_n383), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n389), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT38), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n388), .A2(new_n390), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n417), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n302), .A2(new_n277), .A3(new_n303), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n277), .B1(new_n302), .B2(new_n303), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n307), .A2(new_n428), .B1(KEYINPUT6), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G228gat), .ZN(new_n431));
  INV_X1    g230(.A(G233gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n331), .B2(new_n318), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n259), .B1(new_n434), .B2(KEYINPUT3), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n265), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n381), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT82), .B1(new_n333), .B2(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n435), .A2(new_n433), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n326), .A2(new_n332), .B1(new_n436), .B2(new_n265), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT82), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n433), .B(new_n435), .C1(new_n445), .C2(KEYINPUT82), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n319), .A2(new_n325), .A3(new_n309), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT74), .B1(new_n331), .B2(new_n318), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n437), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n448), .A2(new_n453), .A3(KEYINPUT83), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n440), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G22gat), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT83), .B1(new_n448), .B2(new_n453), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n435), .A2(new_n433), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n452), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n446), .A4(new_n441), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G22gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n440), .ZN(new_n463));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT31), .B(G50gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n456), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n462), .B1(new_n461), .B2(new_n440), .ZN(new_n469));
  AOI211_X1 g268(.A(G22gat), .B(new_n439), .C1(new_n457), .C2(new_n460), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n424), .A2(new_n430), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n395), .A2(new_n407), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(new_n471), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n304), .A2(KEYINPUT6), .A3(new_n271), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n427), .B2(new_n429), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n402), .B(new_n389), .C1(new_n379), .C2(new_n383), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n384), .A2(new_n387), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n392), .B(KEYINPUT75), .C1(new_n387), .C2(new_n384), .ZN(new_n481));
  AND4_X1   g280(.A1(new_n476), .A2(new_n404), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n382), .A2(new_n260), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n382), .A2(new_n260), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G227gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n432), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT34), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  OAI221_X1 g291(.A(new_n492), .B1(new_n489), .B2(new_n432), .C1(new_n486), .C2(new_n487), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G43gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT71), .ZN(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G99gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n362), .A2(new_n375), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n223), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n490), .A3(new_n485), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(KEYINPUT32), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n500), .B(KEYINPUT32), .C1(new_n501), .C2(new_n497), .ZN(new_n505));
  AOI221_X4 g304(.A(new_n484), .B1(new_n491), .B2(new_n493), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n493), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n505), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(KEYINPUT72), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT36), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n507), .A2(new_n504), .A3(new_n505), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n504), .B2(new_n505), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n483), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n473), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n506), .A2(new_n509), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n474), .A2(new_n482), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n512), .A2(new_n513), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n399), .A2(new_n404), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n430), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n474), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT14), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT90), .B(G36gat), .Z(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(G29gat), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT91), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(KEYINPUT89), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(KEYINPUT89), .B2(new_n536), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n534), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n536), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(G1gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n548), .B(new_n551), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n534), .B(new_n538), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n541), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n552), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n543), .A2(new_n556), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n529), .B(new_n554), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n541), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n552), .A3(new_n557), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n554), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n529), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n554), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n543), .A2(new_n553), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n562), .A2(new_n566), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G197gat), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT11), .B(G169gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n566), .A3(new_n580), .A4(new_n572), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n528), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G64gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(G57gat), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT96), .B(G57gat), .Z(new_n588));
  OAI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  OR2_X1    g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n590), .B(new_n591), .C1(new_n594), .C2(new_n592), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n589), .A2(new_n593), .B1(new_n595), .B2(KEYINPUT95), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(KEYINPUT95), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n552), .B1(new_n599), .B2(new_n598), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT97), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G155gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n608), .B(new_n611), .Z(new_n612));
  OR2_X1    g411(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT103), .ZN(new_n618));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT100), .Z(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n618), .B(new_n622), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G99gat), .B(G106gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT7), .ZN(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n627), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n629), .A2(new_n627), .A3(new_n633), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n634), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(KEYINPUT101), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n557), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT102), .B1(new_n641), .B2(new_n559), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n636), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n543), .B2(new_n556), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n564), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n563), .A2(new_n640), .B1(new_n621), .B2(new_n620), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n626), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n649), .B(new_n625), .C1(new_n642), .C2(new_n647), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n624), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n641), .A2(new_n559), .A3(KEYINPUT102), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n646), .B1(new_n645), .B2(new_n564), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n625), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n648), .A2(new_n650), .A3(new_n626), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n623), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n640), .A2(new_n662), .A3(new_n598), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n598), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n598), .A2(new_n639), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n666), .B2(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT105), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n671));
  INV_X1    g470(.A(new_n669), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT10), .B1(new_n664), .B2(new_n665), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n663), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n666), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n669), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n670), .A2(new_n674), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n667), .A2(new_n669), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n669), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n678), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n616), .A2(new_n661), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n585), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n476), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT106), .B(G1gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1324gat));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n523), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n695), .B(new_n701), .C1(new_n696), .C2(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n696), .A2(G8gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(G1325gat));
  INV_X1    g503(.A(new_n690), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n705), .A2(G15gat), .A3(new_n521), .ZN(new_n706));
  INV_X1    g505(.A(new_n515), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1326gat));
  XNOR2_X1  g508(.A(KEYINPUT43), .B(G22gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  INV_X1    g511(.A(new_n474), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n690), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n712), .B1(new_n690), .B2(new_n713), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n716), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n714), .A3(new_n710), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(G29gat), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n616), .A2(new_n661), .A3(new_n686), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n585), .A2(new_n721), .A3(new_n691), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n520), .A2(new_n725), .A3(new_n526), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n520), .B2(new_n526), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n517), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n729), .A3(new_n660), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n661), .B1(new_n517), .B2(new_n527), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n731), .B2(new_n729), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n473), .A2(new_n516), .B1(new_n520), .B2(new_n526), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n733), .B(KEYINPUT44), .C1(new_n734), .C2(new_n661), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n730), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n615), .B(KEYINPUT109), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n737), .A2(new_n582), .A3(new_n687), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n476), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n740), .ZN(G1328gat));
  NOR2_X1   g540(.A1(new_n524), .A2(new_n532), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n585), .A2(new_n722), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT46), .Z(new_n744));
  OAI21_X1  g543(.A(new_n532), .B1(new_n739), .B2(new_n524), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1329gat));
  AND2_X1   g545(.A1(new_n585), .A2(new_n722), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n521), .A2(G43gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n736), .A2(new_n515), .A3(new_n738), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g550(.A(G50gat), .B1(new_n739), .B2(new_n474), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n474), .A2(G50gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n585), .A2(new_n722), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT48), .B1(new_n755), .B2(KEYINPUT112), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n757), .B(new_n758), .C1(new_n752), .C2(new_n754), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n756), .A2(new_n759), .ZN(G1331gat));
  NOR4_X1   g559(.A1(new_n615), .A2(new_n660), .A3(new_n582), .A4(new_n687), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n728), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n691), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT113), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n588), .ZN(G1332gat));
  NOR2_X1   g565(.A1(new_n762), .A2(new_n524), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n762), .B2(new_n707), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n521), .A2(G71gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n763), .A2(new_n713), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n616), .A2(new_n582), .A3(new_n687), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n736), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n736), .A2(KEYINPUT115), .A3(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n691), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n782), .A2(KEYINPUT116), .A3(new_n691), .A4(new_n783), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(G85gat), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n616), .A2(new_n582), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n728), .A2(new_n660), .A3(new_n789), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT51), .Z(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n631), .A3(new_n691), .A4(new_n686), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n524), .A2(new_n687), .A3(G92gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI21_X1  g595(.A(G92gat), .B1(new_n780), .B2(new_n524), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n523), .A3(new_n783), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(KEYINPUT51), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n790), .B(new_n801), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n799), .A2(G92gat), .B1(new_n802), .B2(new_n794), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n803), .B2(new_n796), .ZN(G1337gat));
  INV_X1    g603(.A(G99gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n521), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n805), .A3(new_n806), .A4(new_n686), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n782), .A2(new_n515), .A3(new_n783), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n805), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n474), .A2(G106gat), .A3(new_n687), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n791), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  OAI21_X1  g611(.A(G106gat), .B1(new_n780), .B2(new_n474), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n782), .A2(new_n713), .A3(new_n783), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n815), .A2(G106gat), .B1(new_n802), .B2(new_n810), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n812), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n667), .B2(new_n669), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n670), .A2(new_n819), .A3(new_n674), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n677), .B1(new_n682), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT55), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n681), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n529), .B1(new_n565), .B2(new_n554), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n570), .A2(new_n571), .A3(new_n569), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n577), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n581), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n653), .B2(new_n659), .ZN(new_n832));
  INV_X1    g631(.A(new_n681), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n822), .B2(new_n823), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n825), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n827), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n827), .A2(new_n832), .A3(new_n839), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n827), .A2(new_n582), .A3(new_n836), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n581), .A2(new_n686), .A3(new_n830), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n661), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n737), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n688), .A2(new_n582), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n713), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n523), .A2(new_n476), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n806), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n582), .A2(G113gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n737), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n841), .B2(new_n845), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n848), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n476), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n474), .A3(new_n518), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n523), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n582), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n854), .B1(new_n861), .B2(new_n209), .ZN(G1340gat));
  NOR3_X1   g661(.A1(new_n852), .A2(new_n210), .A3(new_n687), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n686), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n210), .ZN(G1341gat));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n206), .A3(new_n616), .ZN(new_n866));
  OAI21_X1  g665(.A(G127gat), .B1(new_n852), .B2(new_n737), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1342gat));
  NAND2_X1  g667(.A1(new_n660), .A2(new_n524), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT120), .Z(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n204), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n859), .A2(KEYINPUT56), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n852), .B2(new_n661), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT56), .B1(new_n859), .B2(new_n872), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NAND3_X1  g675(.A1(new_n582), .A2(new_n825), .A3(new_n834), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n660), .B1(new_n877), .B2(new_n843), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AND4_X1   g678(.A1(new_n835), .A2(new_n824), .A3(new_n681), .A4(new_n825), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n835), .B1(new_n834), .B2(new_n825), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n839), .B1(new_n882), .B2(new_n832), .ZN(new_n883));
  INV_X1    g682(.A(new_n840), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n848), .B1(new_n885), .B2(new_n615), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n474), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n888), .B(new_n713), .C1(new_n856), .C2(new_n848), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n515), .A2(new_n476), .A3(new_n523), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n582), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n515), .A2(new_n474), .ZN(new_n893));
  INV_X1    g692(.A(G141gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n582), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n858), .A2(new_n524), .A3(new_n893), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n892), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1344gat));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n687), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n257), .A2(KEYINPUT59), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n857), .B2(new_n474), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n661), .A2(new_n831), .A3(new_n826), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n615), .B1(new_n909), .B2(new_n878), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n849), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n888), .A3(new_n713), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n686), .B1(new_n890), .B2(KEYINPUT121), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(KEYINPUT121), .B2(new_n890), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n907), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n858), .A2(new_n524), .A3(new_n893), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n686), .A2(new_n257), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n906), .A2(new_n916), .B1(new_n917), .B2(new_n918), .ZN(G1345gat));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n230), .A3(new_n737), .ZN(new_n920));
  AND4_X1   g719(.A1(new_n524), .A2(new_n858), .A3(new_n616), .A4(new_n893), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  AOI21_X1  g721(.A(G155gat), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT122), .B1(new_n917), .B2(new_n615), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1346gat));
  NAND4_X1  g724(.A1(new_n858), .A2(new_n231), .A3(new_n871), .A4(new_n893), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  OAI21_X1  g726(.A(G162gat), .B1(new_n903), .B2(new_n661), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  NAND4_X1  g728(.A1(new_n474), .A2(new_n476), .A3(new_n518), .A4(new_n523), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n857), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n582), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n524), .A2(new_n521), .A3(new_n691), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n474), .B(new_n933), .C1(new_n856), .C2(new_n848), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n582), .A2(G169gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  INV_X1    g736(.A(G176gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n931), .A2(new_n938), .A3(new_n686), .ZN(new_n939));
  OAI21_X1  g738(.A(G176gat), .B1(new_n934), .B2(new_n687), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n931), .A2(new_n369), .A3(new_n371), .A4(new_n616), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n934), .B2(new_n737), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G183gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n934), .A2(new_n943), .A3(new_n737), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n949), .B(new_n942), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n343), .A3(new_n660), .ZN(new_n952));
  OAI21_X1  g751(.A(G190gat), .B1(new_n934), .B2(new_n661), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n956), .B(G190gat), .C1(new_n934), .C2(new_n661), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n954), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n515), .A2(new_n691), .A3(new_n524), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n713), .B(new_n961), .C1(new_n856), .C2(new_n848), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n582), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n908), .A2(new_n912), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n961), .B(KEYINPUT126), .Z(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n582), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  OR2_X1    g769(.A1(new_n687), .A2(G204gat), .ZN(new_n971));
  OR3_X1    g770(.A1(new_n962), .A2(KEYINPUT127), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT127), .B1(new_n962), .B2(new_n971), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n908), .A2(new_n686), .A3(new_n912), .A4(new_n967), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G204gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n972), .A2(KEYINPUT62), .A3(new_n973), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(G1353gat));
  OR3_X1    g779(.A1(new_n962), .A2(new_n328), .A3(new_n615), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n908), .A2(new_n616), .A3(new_n912), .A4(new_n967), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  NAND3_X1  g784(.A1(new_n965), .A2(new_n660), .A3(new_n967), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G218gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n963), .A2(new_n312), .A3(new_n660), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1355gat));
endmodule


