//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n192), .B1(new_n190), .B2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n199), .A3(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n188), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(new_n196), .A3(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n191), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n201), .B1(new_n190), .B2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n206), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n212), .A2(KEYINPUT81), .A3(G125), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT81), .B1(new_n212), .B2(G125), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G224), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G953), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n215), .B(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT6), .ZN(new_n219));
  XNOR2_X1  g033(.A(G110), .B(G122), .ZN(new_n220));
  XOR2_X1   g034(.A(new_n220), .B(KEYINPUT80), .Z(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n223), .A2(KEYINPUT3), .A3(G107), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(KEYINPUT3), .C1(new_n223), .C2(G107), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(G104), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(G101), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n227), .B(new_n236), .C1(new_n230), .C2(new_n232), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n223), .A2(G107), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n223), .B2(G107), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT77), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n229), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(new_n236), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n235), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT2), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G113), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT68), .A2(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT68), .A2(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(G116), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G119), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G116), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n250), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT68), .A2(G119), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT68), .A2(G119), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n255), .B1(new_n261), .B2(G116), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT69), .B1(new_n262), .B2(new_n250), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n253), .A2(new_n250), .A3(KEYINPUT69), .A4(new_n256), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(new_n256), .A3(new_n250), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n264), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n258), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n245), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(G113), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n236), .B1(new_n231), .B2(new_n239), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n243), .B2(new_n236), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n279), .A3(new_n271), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n222), .B1(new_n274), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n234), .B1(new_n243), .B2(new_n236), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n233), .A2(G101), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n272), .B1(new_n271), .B2(new_n258), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT70), .B(new_n257), .C1(new_n270), .C2(new_n264), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n235), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n280), .A3(new_n220), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n219), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n221), .B1(new_n288), .B2(new_n280), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(KEYINPUT6), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n218), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G210), .B1(G237), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n217), .A2(KEYINPUT84), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n217), .A2(KEYINPUT84), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n205), .B(new_n298), .C1(new_n213), .C2(new_n214), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n217), .A2(new_n295), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT83), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n205), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n195), .A2(KEYINPUT83), .A3(new_n196), .A4(new_n204), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n212), .A2(G125), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n220), .B(KEYINPUT82), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT8), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n277), .A2(new_n271), .ZN(new_n311));
  INV_X1    g125(.A(new_n278), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n237), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n310), .B1(new_n314), .B2(new_n280), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n300), .A2(new_n307), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n316), .B2(new_n289), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n293), .A2(new_n294), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n294), .B1(new_n293), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n187), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT9), .B(G234), .ZN(new_n321));
  OAI21_X1  g135(.A(G221), .B1(new_n321), .B2(G902), .ZN(new_n322));
  XOR2_X1   g136(.A(new_n322), .B(KEYINPUT76), .Z(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n191), .A2(new_n208), .B1(new_n210), .B2(new_n206), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n325), .B(new_n235), .C1(new_n238), .C2(new_n244), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n194), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n204), .B1(new_n210), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n237), .A3(new_n312), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT11), .ZN(new_n332));
  INV_X1    g146(.A(G134), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G137), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT11), .A3(G134), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(G137), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G131), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT65), .B(G131), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(new_n336), .A3(new_n337), .A4(new_n334), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n194), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n344));
  INV_X1    g158(.A(new_n189), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n197), .A2(new_n199), .ZN(new_n346));
  INV_X1    g160(.A(G143), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n204), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n279), .A2(KEYINPUT10), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n326), .A2(new_n331), .A3(new_n343), .A4(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G140), .ZN(new_n352));
  INV_X1    g166(.A(G953), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(G227), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n352), .B(new_n354), .Z(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT79), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n329), .B1(new_n349), .B2(new_n279), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n342), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT12), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(KEYINPUT12), .A3(new_n342), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n313), .A2(new_n195), .A3(new_n204), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n360), .B(new_n343), .C1(new_n365), .C2(new_n329), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT12), .B1(new_n358), .B2(new_n342), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT78), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n351), .A2(new_n369), .A3(new_n355), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n357), .A2(new_n364), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n326), .A2(new_n331), .A3(new_n350), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n342), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n351), .ZN(new_n374));
  INV_X1    g188(.A(new_n355), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI211_X1 g190(.A(G469), .B(G902), .C1(new_n371), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n351), .B1(new_n366), .B2(new_n367), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n375), .ZN(new_n380));
  INV_X1    g194(.A(new_n356), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n373), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G902), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n324), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n320), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G237), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n353), .A3(G210), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT27), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(G101), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n393));
  INV_X1    g207(.A(new_n338), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n335), .A2(KEYINPUT66), .A3(G134), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n333), .B2(G137), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n333), .A2(G137), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n394), .A2(new_n340), .B1(new_n399), .B2(G131), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n342), .A2(new_n325), .B1(new_n349), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n267), .A2(new_n401), .A3(new_n273), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n349), .A2(new_n400), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT67), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n325), .A2(new_n342), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT67), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n349), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n267), .A2(new_n273), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n393), .A2(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n403), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n411), .A2(new_n286), .A3(new_n287), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n392), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT71), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n402), .A2(new_n416), .A3(new_n392), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n402), .B2(new_n392), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n404), .A2(new_n420), .A3(new_n405), .A4(new_n407), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n411), .A2(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n409), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT31), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n392), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT71), .B1(new_n412), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n402), .A2(new_n416), .A3(new_n392), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n427), .A3(KEYINPUT31), .A4(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n415), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G472), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(KEYINPUT32), .A3(new_n432), .A4(new_n384), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT73), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n286), .A2(new_n287), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n401), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n409), .A2(KEYINPUT73), .A3(new_n411), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n402), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT28), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n402), .A2(new_n393), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n439), .A2(KEYINPUT29), .A3(new_n392), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n410), .A2(new_n392), .A3(new_n413), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n412), .B1(new_n423), .B2(new_n409), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n392), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n445), .A3(new_n384), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G472), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT31), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n414), .B1(new_n450), .B2(new_n429), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(G472), .A3(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n433), .B(new_n447), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G125), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n196), .A2(G140), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(KEYINPUT74), .A3(G125), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(KEYINPUT16), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT16), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G146), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n456), .A2(new_n457), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n190), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n261), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G110), .ZN(new_n473));
  NOR2_X1   g287(.A1(G119), .A2(G128), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n261), .B2(new_n194), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G110), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n465), .B(new_n467), .C1(new_n473), .C2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n472), .A2(G110), .B1(new_n476), .B2(new_n478), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n461), .A2(new_n188), .A3(new_n463), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n188), .B1(new_n461), .B2(new_n463), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT22), .B(G137), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n353), .A2(G221), .A3(G234), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n480), .B2(new_n485), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G217), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(G234), .B2(new_n384), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n493), .A2(G902), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n497));
  OAI211_X1 g311(.A(KEYINPUT75), .B(new_n497), .C1(new_n493), .C2(G902), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n480), .A2(new_n485), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n488), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n500), .B2(new_n490), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT75), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT25), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n496), .B1(new_n504), .B2(new_n495), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  INV_X1    g320(.A(G214), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n507), .A2(G237), .A3(G953), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT86), .B1(new_n509), .B2(G143), .ZN(new_n510));
  OR2_X1    g324(.A1(KEYINPUT86), .A2(G143), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n340), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n388), .A2(new_n353), .A3(G214), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(KEYINPUT86), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n512), .A2(new_n513), .A3(new_n516), .A4(KEYINPUT17), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n465), .A2(new_n482), .A3(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n513), .B1(new_n512), .B2(new_n516), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT17), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n523), .A2(KEYINPUT18), .A3(G131), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n512), .A2(new_n524), .A3(new_n516), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n512), .B2(new_n516), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT88), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n459), .A2(new_n528), .A3(new_n460), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n459), .B2(new_n460), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(new_n188), .ZN(new_n531));
  INV_X1    g345(.A(new_n467), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT89), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n522), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT90), .B(G104), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n506), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n540), .B(KEYINPUT91), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  OR3_X1    g358(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT17), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n545), .A2(new_n482), .A3(new_n465), .A4(new_n517), .ZN(new_n546));
  INV_X1    g360(.A(new_n536), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n459), .A2(new_n460), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT88), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n459), .A2(new_n528), .A3(new_n460), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(G146), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n467), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n535), .B1(new_n552), .B2(new_n527), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n546), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT92), .A3(new_n540), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n542), .A2(new_n544), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n384), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(KEYINPUT93), .A3(new_n384), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(G475), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT13), .B1(new_n194), .B2(G143), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n333), .ZN(new_n563));
  XNOR2_X1  g377(.A(G128), .B(G143), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G116), .B(G122), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT94), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n567), .A2(new_n225), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n225), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n225), .ZN(new_n571));
  INV_X1    g385(.A(G116), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G122), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(G122), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(KEYINPUT14), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(KEYINPUT14), .B2(new_n573), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G107), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n564), .B(new_n333), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n321), .A2(new_n494), .A3(G953), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n570), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n570), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n384), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G478), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n466), .A2(KEYINPUT19), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n549), .A2(new_n550), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(KEYINPUT19), .ZN(new_n589));
  OAI221_X1 g403(.A(new_n465), .B1(new_n519), .B2(new_n520), .C1(new_n589), .C2(new_n346), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n547), .B2(new_n553), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n540), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n544), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT20), .ZN(new_n594));
  NOR2_X1   g408(.A1(G475), .A2(G902), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n591), .A2(new_n540), .B1(new_n537), .B2(new_n543), .ZN(new_n597));
  INV_X1    g411(.A(new_n595), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT20), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n586), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n353), .A2(G952), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(G234), .B2(G237), .ZN(new_n602));
  NAND2_X1  g416(.A1(G234), .A2(G237), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(G902), .A3(G953), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(KEYINPUT95), .Z(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT21), .B(G898), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n561), .A2(new_n600), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n387), .A2(new_n454), .A3(new_n505), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  NAND2_X1  g425(.A1(new_n596), .A2(new_n599), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n560), .A2(G475), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT93), .B1(new_n556), .B2(new_n384), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n584), .A2(G902), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n581), .A2(new_n582), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT33), .B1(new_n617), .B2(new_n618), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n583), .A2(new_n584), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n615), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n615), .B2(new_n625), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  INV_X1    g444(.A(new_n294), .ZN(new_n631));
  INV_X1    g445(.A(new_n217), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n215), .B(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n220), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n274), .A2(new_n281), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT6), .B1(new_n635), .B2(new_n291), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n282), .A2(new_n219), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n314), .A2(new_n280), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n309), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n305), .A2(new_n306), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n640), .B(new_n299), .C1(new_n641), .C2(new_n301), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n384), .B1(new_n642), .B2(new_n635), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n631), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n293), .A2(new_n317), .A3(new_n294), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n630), .B1(new_n646), .B2(new_n187), .ZN(new_n647));
  INV_X1    g461(.A(new_n187), .ZN(new_n648));
  AOI211_X1 g462(.A(KEYINPUT96), .B(new_n648), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n608), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n629), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n431), .A2(new_n432), .A3(new_n384), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n451), .B2(G902), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n505), .B(new_n324), .C1(new_n377), .C2(new_n385), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  NAND2_X1  g473(.A1(new_n320), .A2(KEYINPUT96), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n646), .A2(new_n630), .A3(new_n187), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n607), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT99), .B1(new_n613), .B2(new_n614), .ZN(new_n664));
  INV_X1    g478(.A(new_n586), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n599), .B2(new_n596), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n559), .A2(new_n667), .A3(G475), .A4(new_n560), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n662), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n663), .B1(new_n662), .B2(new_n669), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n654), .B(new_n656), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT101), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT35), .B(G107), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  INV_X1    g489(.A(new_n495), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n498), .B2(new_n503), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n499), .B1(KEYINPUT36), .B2(new_n489), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n489), .A2(KEYINPUT36), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n480), .A2(new_n485), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n678), .A2(new_n384), .A3(new_n676), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n652), .A2(new_n653), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n387), .A2(new_n685), .A3(new_n609), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n660), .A2(new_n661), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n605), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n602), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n664), .A2(new_n666), .A3(new_n668), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n677), .A2(new_n683), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n386), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n689), .A2(new_n694), .A3(new_n454), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  AOI21_X1  g512(.A(new_n665), .B1(new_n561), .B2(new_n612), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n187), .A3(new_n695), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n419), .A2(new_n424), .B1(new_n426), .B2(new_n438), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n701), .B2(G902), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n433), .B(new_n702), .C1(new_n452), .C2(new_n453), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n646), .B(KEYINPUT38), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n371), .A2(new_n376), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n378), .A3(new_n384), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n383), .A2(new_n384), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n323), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n693), .B(KEYINPUT39), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT40), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n347), .ZN(G45));
  AND3_X1   g529(.A1(new_n615), .A2(new_n625), .A3(new_n693), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n689), .A2(new_n454), .A3(new_n696), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n615), .A2(new_n625), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT98), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n615), .A2(new_n625), .A3(new_n626), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n662), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n706), .A2(new_n384), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n707), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n323), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n454), .A2(new_n505), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT41), .B(G113), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  INV_X1    g545(.A(new_n728), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n670), .B2(new_n671), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  AOI211_X1 g548(.A(new_n607), .B(new_n586), .C1(new_n599), .C2(new_n596), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n735), .A2(new_n561), .A3(new_n684), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n689), .A2(new_n736), .A3(new_n454), .A4(new_n727), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  AND4_X1   g552(.A1(new_n608), .A2(new_n725), .A3(new_n324), .A4(new_n707), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n699), .B(new_n739), .C1(new_n647), .C2(new_n649), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n653), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT103), .B(G472), .C1(new_n451), .C2(G902), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n425), .A2(new_n430), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n392), .B1(new_n439), .B2(new_n440), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n432), .B(new_n384), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n505), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  AND4_X1   g564(.A1(new_n684), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n689), .A3(new_n716), .A4(new_n727), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  OR2_X1    g567(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n433), .A3(new_n447), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n644), .A2(new_n187), .A3(new_n645), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n756), .A2(new_n386), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n758), .A3(new_n505), .A4(new_n716), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n756), .A2(new_n386), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n716), .A2(new_n454), .A3(new_n505), .A4(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n757), .B1(new_n761), .B2(KEYINPUT104), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n694), .A2(new_n454), .A3(new_n505), .A4(new_n760), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  OR2_X1    g581(.A1(new_n654), .A2(new_n695), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n625), .A2(new_n561), .A3(new_n612), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n769), .A3(new_n773), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(KEYINPUT108), .A3(new_n776), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n768), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT44), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n383), .A2(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n383), .A2(KEYINPUT45), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n378), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n378), .A2(new_n384), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT105), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n790), .B(new_n783), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  INV_X1    g605(.A(new_n786), .ZN(new_n792));
  INV_X1    g606(.A(new_n787), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n789), .A2(new_n707), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n324), .A3(new_n711), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n756), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n782), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(KEYINPUT109), .B(G137), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G39));
  INV_X1    g617(.A(new_n716), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n804), .A2(new_n454), .A3(new_n505), .A4(new_n756), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n324), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT47), .B1(new_n795), .B2(new_n324), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND2_X1  g624(.A1(new_n795), .A2(new_n324), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n806), .C1(new_n324), .C2(new_n726), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n692), .B1(new_n775), .B2(new_n776), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n748), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n798), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n727), .A2(new_n648), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n704), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n748), .A4(new_n821), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n727), .A2(new_n798), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n692), .B(new_n826), .C1(new_n775), .C2(new_n776), .ZN(new_n827));
  INV_X1    g641(.A(new_n505), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n826), .A2(new_n703), .A3(new_n828), .A4(new_n692), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n615), .A2(new_n625), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n827), .A2(new_n751), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n818), .A2(new_n825), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n827), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n755), .A2(new_n505), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT48), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT48), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n827), .A2(new_n841), .A3(new_n505), .A4(new_n755), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n844));
  OAI211_X1 g658(.A(KEYINPUT116), .B(KEYINPUT48), .C1(new_n836), .C2(new_n837), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n840), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n689), .A2(new_n815), .A3(new_n727), .A4(new_n748), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n601), .B(new_n847), .C1(new_n722), .C2(new_n829), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n835), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n833), .A2(new_n834), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n693), .B(KEYINPUT111), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n710), .A2(new_n695), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n689), .A2(new_n703), .A3(new_n699), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n752), .A2(new_n697), .A3(new_n717), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n454), .A2(new_n696), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n689), .C1(new_n694), .C2(new_n716), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n857), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n607), .B(new_n648), .C1(new_n644), .C2(new_n645), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n612), .B(new_n586), .C1(new_n613), .C2(new_n614), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n654), .A2(new_n866), .A3(new_n656), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n735), .A3(new_n710), .A4(new_n561), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n652), .A2(new_n653), .A3(new_n684), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n865), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n654), .A2(new_n866), .A3(new_n656), .A4(new_n868), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n686), .A2(new_n875), .A3(KEYINPUT110), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n748), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n723), .A2(new_n728), .B1(new_n878), .B2(new_n740), .ZN(new_n879));
  INV_X1    g693(.A(new_n719), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n654), .A3(new_n656), .A4(new_n866), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n737), .A2(new_n610), .A3(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n877), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n743), .A2(new_n744), .A3(new_n747), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n664), .A2(new_n600), .A3(new_n668), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n884), .A2(new_n880), .B1(new_n454), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n760), .A2(new_n684), .A3(new_n693), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n766), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n454), .A2(new_n505), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT104), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n716), .A4(new_n760), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n757), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n893), .B2(new_n759), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n864), .A2(new_n883), .A3(new_n733), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT112), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n686), .A2(KEYINPUT110), .A3(new_n875), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT110), .B1(new_n686), .B2(new_n875), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n651), .A2(new_n732), .B1(new_n741), .B2(new_n748), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n737), .A2(new_n610), .A3(new_n881), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n733), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(KEYINPUT53), .A3(new_n864), .A4(new_n894), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT112), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n899), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n853), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(G952), .A2(G953), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR4_X1    g730(.A1(new_n828), .A2(new_n704), .A3(new_n648), .A4(new_n323), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n726), .B(KEYINPUT49), .ZN(new_n918));
  OR4_X1    g732(.A1(new_n703), .A2(new_n917), .A3(new_n770), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(G75));
  XOR2_X1   g734(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n290), .A2(new_n292), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n633), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n924), .A2(new_n293), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n384), .B1(new_n899), .B2(new_n907), .ZN(new_n926));
  AOI211_X1 g740(.A(KEYINPUT56), .B(new_n925), .C1(new_n926), .C2(G210), .ZN(new_n927));
  INV_X1    g741(.A(new_n925), .ZN(new_n928));
  INV_X1    g742(.A(new_n888), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n764), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n905), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n931), .B2(new_n864), .ZN(new_n932));
  OAI211_X1 g746(.A(G210), .B(G902), .C1(new_n897), .C2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n922), .B1(new_n927), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(G210), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n937), .B(new_n384), .C1(new_n899), .C2(new_n907), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n925), .B1(new_n938), .B2(KEYINPUT56), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n933), .A2(new_n934), .A3(new_n928), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n940), .A3(new_n921), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n353), .A2(G952), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n936), .A2(new_n941), .A3(new_n943), .ZN(G51));
  XOR2_X1   g758(.A(new_n706), .B(KEYINPUT118), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n899), .A2(new_n907), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n912), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n787), .B(KEYINPUT57), .Z(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n926), .A2(new_n786), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n597), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n597), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n942), .ZN(G60));
  OR2_X1    g769(.A1(new_n621), .A2(new_n622), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT119), .Z(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  OR2_X1    g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n943), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n911), .A2(new_n913), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(new_n957), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n899), .B2(new_n907), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n942), .B1(new_n970), .B2(new_n493), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n678), .A2(new_n680), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT120), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n969), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n971), .B(KEYINPUT61), .C1(new_n975), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G66));
  NOR3_X1   g795(.A1(new_n606), .A2(new_n216), .A3(new_n353), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n905), .B(KEYINPUT122), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n353), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n923), .B1(G898), .B2(new_n353), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G69));
  INV_X1    g800(.A(new_n766), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n505), .A2(new_n755), .A3(new_n689), .A4(new_n699), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n797), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n862), .A2(new_n752), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n809), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n801), .A2(new_n764), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT124), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n801), .A2(new_n995), .A3(new_n764), .A4(new_n992), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(new_n353), .A3(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n589), .B(KEYINPUT123), .Z(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n423), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(G900), .B2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n712), .A2(new_n756), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n889), .B(new_n1002), .C1(new_n880), .C2(new_n868), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n809), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n990), .B2(new_n714), .ZN(new_n1006));
  OR3_X1    g820(.A1(new_n990), .A2(new_n714), .A3(new_n1005), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1008), .A2(new_n801), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n999), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT125), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n999), .A2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n353), .B(new_n1013), .C1(G227), .C2(G900), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1014), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1001), .A2(new_n1010), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n1009), .B2(new_n983), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n444), .A2(new_n426), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(KEYINPUT126), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT126), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n983), .A2(new_n801), .A3(new_n1008), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1026), .B(new_n1023), .C1(new_n1027), .C2(new_n1021), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n942), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n994), .A2(new_n983), .A3(new_n996), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n1020), .ZN(new_n1031));
  INV_X1    g845(.A(new_n444), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1032), .A2(new_n392), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n426), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1021), .B1(new_n1034), .B2(new_n448), .ZN(new_n1035));
  AOI22_X1  g849(.A1(new_n1031), .A2(new_n1033), .B1(new_n910), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n1029), .A2(new_n1036), .ZN(G57));
endmodule


