//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n202), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G77), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n212), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G1), .B2(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n206), .A2(G13), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(G257), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n210), .B(new_n236), .C1(new_n237), .C2(new_n215), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n234), .B1(KEYINPUT0), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g0039(.A(new_n225), .B(new_n239), .C1(KEYINPUT0), .C2(new_n238), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G250), .B(G257), .Z(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT66), .ZN(new_n251));
  XOR2_X1   g0051(.A(G50), .B(G58), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  AND2_X1   g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n228), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n264), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT68), .B(G226), .Z(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n265), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G274), .A3(new_n260), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n226), .A2(G1), .A3(G13), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n262), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n284), .C1(G77), .C2(new_n277), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n272), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n271), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(KEYINPUT70), .A3(new_n285), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n289), .A2(new_n292), .A3(G200), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n289), .B2(new_n292), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n282), .A2(new_n283), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G1), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n303), .A2(new_n202), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n203), .A2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(G150), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT71), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(new_n207), .A3(KEYINPUT8), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n231), .A2(G33), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n307), .B1(new_n308), .B2(new_n310), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n306), .B1(new_n298), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n301), .A2(new_n202), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT9), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n296), .B(new_n321), .C1(KEYINPUT74), .C2(KEYINPUT10), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT70), .B1(new_n291), .B2(new_n285), .ZN(new_n323));
  AND4_X1   g0123(.A1(KEYINPUT70), .A2(new_n272), .A3(new_n285), .A4(new_n286), .ZN(new_n324));
  OAI21_X1  g0124(.A(G190), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n289), .A2(new_n292), .A3(G200), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(KEYINPUT74), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n321), .A3(new_n326), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT10), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n323), .A2(new_n324), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(new_n320), .C1(G179), .C2(new_n331), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n322), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n213), .A2(new_n278), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n208), .A2(G1698), .ZN(new_n337));
  AND2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NOR2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(KEYINPUT75), .A3(new_n341), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n284), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n266), .A2(G238), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n270), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .A4(new_n270), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G77), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n310), .A2(new_n202), .B1(new_n316), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n231), .A2(G68), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n298), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g0159(.A(new_n359), .B(KEYINPUT11), .Z(new_n360));
  XNOR2_X1  g0160(.A(new_n300), .B(KEYINPUT72), .ZN(new_n361));
  INV_X1    g0161(.A(new_n298), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n304), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n221), .B1(new_n363), .B2(KEYINPUT12), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n301), .A2(KEYINPUT12), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT72), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n300), .B(new_n366), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n367), .A2(KEYINPUT12), .A3(new_n221), .ZN(new_n368));
  NOR4_X1   g0168(.A1(new_n360), .A2(new_n364), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n294), .B2(new_n352), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n353), .A2(G179), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT14), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n373), .A4(G169), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT76), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n352), .A2(new_n375), .A3(KEYINPUT77), .A4(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n375), .B1(new_n352), .B2(G169), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n372), .B(new_n374), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n369), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n367), .A2(new_n356), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n311), .A2(new_n310), .B1(new_n383), .B2(new_n316), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(G20), .B2(G77), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n382), .B1(new_n363), .B2(new_n356), .C1(new_n385), .C2(new_n362), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G238), .A2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n277), .B(new_n390), .C1(new_n208), .C2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n284), .C1(G107), .C2(new_n277), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n266), .A2(new_n218), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n270), .A3(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n388), .A2(new_n389), .B1(new_n332), .B2(new_n394), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(G179), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n381), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n335), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n338), .A2(new_n339), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n400), .B2(new_n231), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n276), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n309), .A2(G159), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n201), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n405), .A4(new_n408), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n298), .A3(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n303), .A2(new_n315), .A3(new_n305), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n301), .B2(new_n315), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n280), .A2(new_n278), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n213), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n338), .C2(new_n339), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT78), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(KEYINPUT78), .A3(new_n420), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n284), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n266), .A2(G232), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n270), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n354), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n294), .A3(new_n270), .A4(new_n426), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT79), .B1(new_n416), .B2(new_n430), .ZN(new_n431));
  AND4_X1   g0231(.A1(KEYINPUT79), .A2(new_n430), .A3(new_n415), .A4(new_n413), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT17), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT80), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n416), .A2(new_n430), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT17), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n428), .A2(new_n429), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n413), .A2(new_n415), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n430), .A2(KEYINPUT79), .A3(new_n415), .A4(new_n413), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT80), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT17), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n434), .A2(new_n437), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n427), .A2(new_n332), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n440), .B(new_n447), .C1(G179), .C2(new_n427), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n394), .A2(new_n294), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n394), .A2(G200), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n388), .A2(new_n451), .A3(new_n389), .A4(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n446), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n399), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G20), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n231), .C1(G33), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n298), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n298), .A2(KEYINPUT20), .A3(new_n457), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n367), .A2(new_n456), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n299), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n361), .A2(G116), .A3(new_n362), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G264), .A2(G1698), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n470), .B1(new_n237), .B2(G1698), .C1(new_n338), .C2(new_n339), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT84), .B(G303), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n284), .C1(new_n277), .C2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n259), .A2(G1), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G41), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n269), .A2(G274), .A3(new_n478), .A4(new_n260), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n269), .A2(G270), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n469), .A2(G169), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G179), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n469), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n469), .A2(KEYINPUT21), .A3(G169), .A4(new_n482), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n269), .A2(G257), .A3(new_n480), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT81), .ZN(new_n493));
  OAI21_X1  g0293(.A(G244), .B1(new_n338), .B2(new_n339), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(G1698), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(G244), .C1(new_n339), .C2(new_n338), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n458), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n277), .A2(G250), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n278), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n284), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n479), .A2(new_n503), .A3(new_n491), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n493), .A2(new_n502), .A3(new_n486), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n302), .A2(new_n467), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G97), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n300), .A2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n275), .A2(new_n231), .A3(new_n276), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT7), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n214), .B1(new_n513), .B2(new_n402), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n459), .A2(new_n214), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n231), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n310), .A2(new_n356), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n508), .B(new_n510), .C1(new_n522), .C2(new_n362), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n264), .B1(new_n227), .B2(new_n229), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n496), .A2(new_n458), .A3(new_n498), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n332), .B1(new_n528), .B2(new_n492), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n505), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n493), .A2(new_n502), .A3(new_n504), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  INV_X1    g0332(.A(new_n492), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n502), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT82), .B1(new_n534), .B2(new_n294), .ZN(new_n535));
  INV_X1    g0335(.A(new_n523), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n533), .A2(new_n502), .A3(new_n537), .A4(G190), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n532), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n469), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n482), .A2(G200), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n294), .C2(new_n482), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n490), .A2(new_n530), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n231), .B(G87), .C1(new_n338), .C2(new_n339), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n277), .A2(new_n548), .A3(new_n231), .A4(G87), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n231), .A2(G107), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT23), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n550), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT24), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n547), .A2(new_n549), .ZN(new_n557));
  INV_X1    g0357(.A(new_n545), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n553), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT85), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n298), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n277), .B1(G257), .B2(new_n278), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G250), .A2(G1698), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n284), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n269), .A2(G264), .A3(new_n480), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n479), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n354), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G190), .B2(new_n572), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  AOI211_X1 g0376(.A(G107), .B(new_n300), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(new_n507), .B2(G107), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n565), .A2(new_n574), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n572), .A2(new_n332), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n572), .A2(G179), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n362), .B1(new_n556), .B2(new_n563), .ZN(new_n585));
  INV_X1    g0385(.A(new_n581), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n209), .A2(new_n459), .A3(new_n214), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n341), .A2(new_n231), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT19), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n231), .B(G68), .C1(new_n338), .C2(new_n339), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n316), .B2(new_n459), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n298), .B1(new_n367), .B2(new_n383), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n302), .A2(G87), .A3(new_n467), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n222), .A2(new_n278), .ZN(new_n598));
  INV_X1    g0398(.A(G244), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G1698), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n600), .C1(new_n338), .C2(new_n339), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n544), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n284), .ZN(new_n603));
  AOI21_X1  g0403(.A(G250), .B1(new_n299), .B2(G45), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n259), .A2(G1), .A3(G274), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n269), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n354), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT83), .B1(new_n597), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n524), .B1(new_n544), .B2(new_n601), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n604), .B(new_n606), .C1(new_n263), .C2(new_n265), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n595), .A4(new_n596), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n603), .A2(new_n608), .A3(G190), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n332), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n594), .A2(new_n298), .ZN(new_n619));
  INV_X1    g0419(.A(new_n383), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n362), .A2(new_n300), .A3(new_n620), .A4(new_n467), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n367), .A2(new_n383), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n603), .A2(new_n608), .A3(new_n486), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n582), .A2(new_n587), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n455), .A2(new_n543), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n455), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n485), .A2(KEYINPUT88), .A3(new_n488), .A4(new_n489), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n587), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT89), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n586), .B1(new_n564), .B2(new_n298), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n613), .A2(new_n595), .A3(new_n596), .A4(new_n616), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n625), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(KEYINPUT87), .A3(new_n625), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n637), .A2(new_n574), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n539), .A2(new_n530), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n632), .A2(new_n633), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n587), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n636), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n530), .B1(new_n641), .B2(new_n642), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT90), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n505), .A2(new_n523), .A3(new_n529), .ZN(new_n653));
  INV_X1    g0453(.A(new_n642), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT87), .B1(new_n638), .B2(new_n625), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n653), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n652), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n625), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n650), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n629), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n334), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n444), .B1(new_n443), .B2(KEYINPUT17), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT17), .ZN(new_n667));
  AOI211_X1 g0467(.A(KEYINPUT80), .B(new_n667), .C1(new_n441), .C2(new_n442), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n666), .A2(new_n668), .A3(new_n436), .ZN(new_n669));
  INV_X1    g0469(.A(new_n371), .ZN(new_n670));
  INV_X1    g0470(.A(new_n397), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n380), .A2(new_n379), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n450), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n322), .A2(new_n330), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n665), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n664), .A2(new_n675), .ZN(G369));
  INV_X1    g0476(.A(G13), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G20), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n299), .ZN(new_n679));
  XNOR2_X1  g0479(.A(KEYINPUT91), .B(KEYINPUT27), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(KEYINPUT92), .B(G343), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n540), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n634), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n542), .A2(new_n485), .A3(new_n488), .A4(new_n489), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT93), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n582), .A2(new_n587), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n637), .B2(new_n687), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n587), .B2(new_n687), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n490), .A2(new_n686), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n695), .A2(new_n699), .B1(new_n635), .B2(new_n687), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(G399));
  NOR2_X1   g0501(.A1(new_n236), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n588), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n233), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n651), .A2(new_n658), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n653), .A2(new_n617), .A3(new_n658), .A4(new_n625), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n625), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n587), .A2(new_n490), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n643), .A3(new_n645), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n708), .B1(new_n715), .B2(new_n687), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n686), .B1(new_n650), .B2(new_n662), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n708), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n531), .A2(KEYINPUT95), .A3(new_n572), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n720), .A2(new_n486), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n603), .A2(new_n608), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n531), .A2(new_n572), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n721), .A2(new_n482), .A3(new_n722), .A4(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(KEYINPUT94), .A2(KEYINPUT30), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n528), .A2(new_n482), .A3(new_n492), .A4(new_n486), .ZN(new_n728));
  AND4_X1   g0528(.A1(new_n570), .A2(new_n571), .A3(new_n603), .A4(new_n608), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n528), .A2(new_n492), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n731), .A2(new_n729), .A3(new_n487), .A4(new_n727), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n687), .B1(new_n726), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n627), .A2(new_n543), .A3(new_n686), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n725), .A2(new_n482), .A3(new_n722), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n720), .A2(new_n486), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n733), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n719), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n718), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n707), .B1(new_n746), .B2(G1), .ZN(G364));
  NAND2_X1  g0547(.A1(new_n678), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n703), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n231), .A2(G190), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n486), .A3(new_n354), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT98), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT98), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G159), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n294), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n231), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n459), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n354), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n486), .A2(new_n354), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n750), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n277), .B1(new_n762), .B2(new_n214), .C1(new_n221), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n231), .A2(new_n294), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n486), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G50), .A2(new_n768), .B1(new_n771), .B2(G58), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n750), .A2(new_n769), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n766), .A2(new_n761), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n772), .B1(new_n356), .B2(new_n773), .C1(new_n209), .C2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n757), .A2(new_n760), .A3(new_n765), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  INV_X1    g0577(.A(new_n762), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n755), .A2(G329), .B1(G283), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT100), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n768), .A2(G326), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n400), .B1(new_n759), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n773), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G322), .A2(new_n771), .B1(new_n784), .B2(G311), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT33), .B(G317), .Z(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n764), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n774), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n783), .B(new_n787), .C1(G303), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n780), .A2(new_n781), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n230), .B1(G20), .B2(new_n332), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n749), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT97), .Z(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n792), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n236), .A2(new_n277), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n233), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n253), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n277), .A2(new_n235), .ZN(new_n802));
  INV_X1    g0602(.A(G355), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n803), .B1(G116), .B2(new_n235), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n797), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n796), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n793), .B(new_n805), .C1(new_n691), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n693), .A2(new_n749), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n692), .A2(G330), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n397), .A2(new_n686), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n388), .A2(new_n389), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n686), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(new_n453), .B1(new_n395), .B2(new_n396), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n717), .B(new_n815), .ZN(new_n816));
  OR3_X1    g0616(.A1(new_n816), .A2(KEYINPUT103), .A3(new_n744), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT103), .B1(new_n816), .B2(new_n744), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n749), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT104), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n816), .A2(new_n744), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n817), .A2(KEYINPUT104), .A3(new_n749), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n792), .ZN(new_n825));
  INV_X1    g0625(.A(new_n764), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G143), .A2(new_n771), .B1(new_n826), .B2(G150), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n768), .A2(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n773), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n778), .A2(G68), .ZN(new_n832));
  INV_X1    g0632(.A(new_n759), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G58), .B1(new_n788), .B2(G50), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n400), .B1(new_n755), .B2(G132), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n831), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G107), .A2(new_n788), .B1(new_n784), .B2(G116), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n209), .B2(new_n762), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n400), .B1(new_n770), .B2(new_n782), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n768), .A2(G303), .ZN(new_n840));
  NOR4_X1   g0640(.A1(new_n838), .A2(new_n760), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n764), .A2(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n764), .A2(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n841), .B1(new_n842), .B2(new_n845), .C1(new_n846), .C2(new_n754), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n825), .B1(new_n836), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n795), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n792), .A2(new_n849), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n749), .B(new_n848), .C1(new_n356), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT102), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n795), .B2(new_n815), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n824), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(new_n683), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n440), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n446), .B2(new_n450), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n448), .A2(KEYINPUT105), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n448), .A2(KEYINPUT105), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n858), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n441), .B2(new_n442), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n448), .A2(new_n435), .A3(new_n858), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n862), .A2(new_n864), .B1(KEYINPUT37), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n856), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n864), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n443), .A2(new_n448), .A3(new_n858), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n666), .A2(new_n668), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n449), .B1(new_n872), .B2(new_n437), .ZN(new_n873));
  OAI211_X1 g0673(.A(KEYINPUT38), .B(new_n871), .C1(new_n873), .C2(new_n858), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT106), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n742), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n734), .A2(KEYINPUT106), .A3(KEYINPUT31), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n738), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n815), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n369), .A2(new_n687), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n381), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n379), .A2(new_n380), .A3(new_n686), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n875), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n862), .A2(new_n864), .B1(KEYINPUT37), .B2(new_n869), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n856), .B1(new_n859), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n874), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT40), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n629), .A2(new_n879), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(G330), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n863), .B1(new_n669), .B2(new_n449), .ZN(new_n897));
  INV_X1    g0697(.A(new_n866), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n859), .A2(new_n856), .A3(new_n888), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n379), .A2(new_n380), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n686), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n889), .A2(new_n874), .A3(KEYINPUT39), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n450), .A2(new_n857), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n717), .A2(new_n815), .ZN(new_n908));
  INV_X1    g0708(.A(new_n811), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n883), .A2(new_n884), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n890), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n905), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n675), .B1(new_n718), .B2(new_n455), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n913), .B(new_n914), .Z(new_n915));
  XNOR2_X1  g0715(.A(new_n895), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n299), .B2(new_n678), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n518), .A2(new_n519), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n231), .B(new_n230), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(G116), .C1(new_n919), .C2(new_n918), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n406), .A2(G77), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n233), .A2(new_n923), .B1(G50), .B2(new_n221), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n677), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n922), .A3(new_n925), .ZN(G367));
  XNOR2_X1  g0726(.A(new_n702), .B(KEYINPUT41), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n645), .B1(new_n536), .B2(new_n687), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n530), .B2(new_n687), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n700), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT107), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT45), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n930), .A2(new_n700), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(KEYINPUT44), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n934), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n698), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n695), .A2(new_n699), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n697), .B2(new_n699), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n693), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n745), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT108), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n939), .A2(new_n947), .A3(new_n940), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n941), .A2(new_n945), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n928), .B1(new_n949), .B2(new_n746), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT109), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n748), .A2(G1), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n940), .A2(new_n930), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n597), .A2(new_n686), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n654), .B2(new_n655), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n625), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n957), .B(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n942), .A2(new_n929), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT42), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n530), .B1(new_n929), .B2(new_n587), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n687), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n965), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n963), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n956), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n788), .A2(G116), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT46), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n277), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n972), .B2(new_n971), .C1(new_n214), .C2(new_n759), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G311), .B2(new_n768), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n778), .A2(G97), .ZN(new_n976));
  INV_X1    g0776(.A(new_n472), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n976), .B1(new_n977), .B2(new_n770), .C1(new_n845), .C2(new_n782), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G317), .B2(new_n755), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n975), .B(new_n979), .C1(new_n842), .C2(new_n773), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n759), .A2(new_n221), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n768), .A2(G143), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n202), .B2(new_n773), .C1(new_n207), .C2(new_n774), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(G150), .C2(new_n771), .ZN(new_n984));
  INV_X1    g0784(.A(new_n845), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G137), .A2(new_n755), .B1(new_n985), .B2(G159), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n277), .B1(new_n762), .B2(new_n356), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT110), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n980), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n749), .B1(new_n991), .B2(new_n792), .ZN(new_n992));
  INV_X1    g0792(.A(new_n798), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n797), .B1(new_n235), .B2(new_n383), .C1(new_n248), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n959), .A2(new_n796), .A3(new_n960), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n970), .A2(new_n996), .ZN(G387));
  AND2_X1   g0797(.A1(new_n755), .A2(G326), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G322), .A2(new_n768), .B1(new_n771), .B2(G317), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n977), .B2(new_n773), .C1(new_n845), .C2(new_n846), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n842), .B2(new_n759), .C1(new_n782), .C2(new_n774), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n277), .B(new_n998), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .C1(new_n456), .C2(new_n762), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G50), .A2(new_n771), .B1(new_n784), .B2(G68), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n356), .B2(new_n774), .C1(new_n829), .C2(new_n767), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n759), .A2(new_n383), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1007), .A2(new_n400), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n826), .A2(new_n312), .A3(new_n314), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n755), .A2(G150), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1009), .A2(new_n976), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n825), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n798), .B1(new_n245), .B2(new_n259), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n704), .B2(new_n802), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n221), .A2(new_n356), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n311), .A2(G50), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G116), .B(new_n588), .C1(new_n1017), .C2(KEYINPUT50), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n259), .C1(KEYINPUT50), .C2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(G107), .B2(new_n235), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1013), .B1(new_n797), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n749), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n697), .C2(new_n806), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n944), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n702), .B1(new_n1025), .B2(new_n746), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1024), .B1(new_n955), .B2(new_n944), .C1(new_n1026), .C2(new_n945), .ZN(G393));
  XNOR2_X1  g0827(.A(new_n939), .B(new_n940), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n745), .B2(new_n944), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n949), .A3(new_n702), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1028), .A2(new_n955), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n985), .A2(G50), .B1(G77), .B2(new_n833), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n311), .B2(new_n773), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT111), .Z(new_n1034));
  OAI22_X1  g0834(.A1(new_n767), .A2(new_n308), .B1(new_n770), .B2(new_n829), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT51), .Z(new_n1036));
  AOI211_X1 g0836(.A(new_n400), .B(new_n1036), .C1(G68), .C2(new_n788), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n755), .A2(G143), .B1(G87), .B2(new_n778), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT112), .Z(new_n1040));
  AOI22_X1  g0840(.A1(G317), .A2(new_n768), .B1(new_n771), .B2(G311), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1041), .A2(KEYINPUT52), .B1(new_n845), .B2(new_n977), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT52), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n755), .A2(G322), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n774), .A2(new_n842), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n400), .B1(new_n762), .B2(new_n214), .C1(new_n782), .C2(new_n773), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G116), .C2(new_n833), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1040), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n749), .B1(new_n1049), .B2(new_n792), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n797), .B1(new_n459), .B2(new_n235), .C1(new_n256), .C2(new_n993), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n806), .C2(new_n930), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1030), .A2(new_n1031), .A3(new_n1052), .ZN(G390));
  INV_X1    g0853(.A(new_n903), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n811), .B1(new_n717), .B2(new_n815), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n884), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n381), .B2(new_n882), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1054), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n889), .A2(new_n874), .A3(KEYINPUT39), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT39), .B1(new_n867), .B2(new_n874), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n738), .A2(new_n742), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n815), .A2(G330), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n911), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT114), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n686), .B(new_n814), .C1(new_n712), .C2(new_n714), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT113), .B1(new_n1067), .B2(new_n811), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n814), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n715), .A2(new_n687), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT113), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n909), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n911), .A3(new_n1072), .ZN(new_n1073));
  AND4_X1   g0873(.A1(new_n1066), .A2(new_n875), .A3(new_n1073), .A4(new_n1054), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n903), .B1(new_n867), .B2(new_n874), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1066), .B1(new_n1075), .B2(new_n1073), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1061), .B(new_n1065), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n875), .A2(new_n1073), .A3(new_n1054), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT114), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n901), .A2(new_n904), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1079), .A2(new_n1080), .B1(new_n1081), .B2(new_n1058), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n644), .A2(new_n690), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n695), .A2(new_n1083), .A3(new_n626), .A4(new_n687), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n734), .B1(new_n1084), .B2(KEYINPUT31), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n877), .A2(new_n878), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1087), .A2(new_n1057), .A3(new_n1063), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1077), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n911), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n910), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1057), .B1(new_n1087), .B2(new_n1063), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1065), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n879), .A2(new_n399), .A3(G330), .A4(new_n454), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n675), .C1(new_n718), .C2(new_n455), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT115), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1090), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1077), .C1(new_n1082), .C2(new_n1089), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n702), .A3(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1090), .A2(new_n955), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1081), .A2(new_n849), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n850), .A2(new_n315), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  AOI22_X1  g0909(.A1(G132), .A2(new_n771), .B1(new_n784), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n768), .A2(G128), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n829), .C2(new_n759), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G137), .B2(new_n985), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n774), .A2(new_n308), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n277), .B1(new_n762), .B2(new_n202), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G125), .B2(new_n755), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1113), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT117), .Z(new_n1120));
  OAI21_X1  g0920(.A(new_n832), .B1(new_n754), .B2(new_n782), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT118), .Z(new_n1122));
  AOI22_X1  g0922(.A1(G283), .A2(new_n768), .B1(new_n771), .B2(G116), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n209), .B2(new_n774), .C1(new_n459), .C2(new_n773), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G77), .B2(new_n833), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n277), .B1(new_n985), .B2(G107), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n749), .B1(new_n1128), .B2(new_n792), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1107), .A2(new_n1108), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1105), .A2(new_n1106), .A3(new_n1130), .ZN(G378));
  OAI211_X1 g0931(.A(new_n1077), .B(new_n1096), .C1(new_n1082), .C2(new_n1089), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1099), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT122), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n887), .A2(new_n891), .A3(new_n719), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n913), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n875), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n879), .A2(new_n885), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n874), .B2(new_n889), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(G330), .C1(KEYINPUT40), .C2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n907), .A3(new_n905), .A4(new_n912), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n335), .B(KEYINPUT55), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n320), .A2(new_n857), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1145), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n1144), .A3(new_n1149), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1137), .A2(new_n1142), .A3(new_n1155), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1132), .A2(KEYINPUT122), .A3(new_n1099), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1135), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1135), .A2(new_n1159), .A3(KEYINPUT57), .A4(new_n1160), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n702), .A3(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1137), .A2(new_n1142), .A3(new_n1155), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1155), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n954), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n202), .B1(new_n338), .B2(G41), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n773), .A2(new_n383), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n826), .B1(new_n771), .B2(G107), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n221), .B2(new_n759), .C1(new_n456), .C2(new_n767), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n755), .A2(G283), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n778), .A2(G58), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n788), .B2(G77), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1173), .A2(new_n400), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1170), .B(new_n1172), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1169), .B1(new_n1179), .B2(KEYINPUT58), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n833), .A2(G150), .B1(new_n768), .B2(G125), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G128), .A2(new_n771), .B1(new_n788), .B2(new_n1109), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n826), .A2(G132), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n784), .A2(G137), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G33), .B1(new_n778), .B2(G159), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G41), .B1(new_n755), .B2(G124), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1194), .A2(new_n792), .B1(new_n202), .B2(new_n850), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1023), .B(new_n1195), .C1(new_n1156), .C2(new_n795), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1168), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1165), .A2(new_n1198), .ZN(G375));
  NAND3_X1  g0999(.A1(new_n1098), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1100), .A2(new_n927), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1057), .A2(new_n849), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G132), .A2(new_n768), .B1(new_n771), .B2(G137), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n308), .B2(new_n773), .C1(new_n829), .C2(new_n774), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n400), .B(new_n1204), .C1(G50), .C2(new_n833), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n755), .A2(G128), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n985), .A2(new_n1109), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1205), .A2(new_n1174), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G97), .A2(new_n788), .B1(new_n771), .B2(G283), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n214), .B2(new_n773), .C1(new_n782), .C2(new_n767), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G77), .B2(new_n778), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G303), .A2(new_n755), .B1(new_n985), .B2(G116), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n383), .C2(new_n759), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1208), .B1(new_n277), .B2(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1214), .A2(new_n792), .B1(new_n221), .B2(new_n850), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1202), .A2(new_n1023), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1096), .B2(new_n954), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1201), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n970), .A2(new_n996), .A3(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G378), .A2(new_n1197), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1165), .A2(new_n1221), .ZN(new_n1222));
  OR3_X1    g1022(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1223));
  OR4_X1    g1023(.A1(G381), .A2(new_n1220), .A3(new_n1222), .A4(new_n1223), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n685), .A2(G213), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT123), .Z(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(new_n1222), .C2(new_n1226), .ZN(G409));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1165), .B2(new_n1198), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1132), .A2(KEYINPUT122), .A3(new_n1099), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT122), .B1(new_n1132), .B2(new_n1099), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1232), .A2(KEYINPUT124), .A3(new_n927), .A4(new_n1159), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1135), .A2(new_n1159), .A3(new_n927), .A4(new_n1160), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1221), .A2(new_n1233), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1225), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1200), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1239), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT60), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1098), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1245));
  OAI211_X1 g1045(.A(KEYINPUT125), .B(new_n1200), .C1(new_n1245), .C2(new_n1240), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n702), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT126), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1217), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n854), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1217), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT126), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1250), .B(new_n1252), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1229), .A2(new_n1237), .A3(new_n1238), .A4(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT127), .B1(new_n1254), .B2(KEYINPUT63), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1229), .A2(new_n1237), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1253), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1226), .A4(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1221), .A2(new_n1233), .A3(new_n1236), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1225), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1252), .A2(new_n854), .A3(new_n1249), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1251), .A2(KEYINPUT126), .A3(G384), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1262), .A2(new_n1263), .B1(G2897), .B2(new_n1238), .ZN(new_n1264));
  INV_X1    g1064(.A(G2897), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1226), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1253), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1259), .A2(new_n1225), .A3(new_n1260), .A4(new_n1257), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1255), .A2(new_n1258), .A3(new_n1268), .A4(new_n1272), .ZN(new_n1273));
  XOR2_X1   g1073(.A(G393), .B(G396), .Z(new_n1274));
  AOI21_X1  g1074(.A(new_n1219), .B1(new_n970), .B2(new_n996), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n996), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1276), .B(G390), .C1(new_n956), .C2(new_n969), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n969), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n950), .B(KEYINPUT109), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n955), .ZN(new_n1281));
  OAI21_X1  g1081(.A(G390), .B1(new_n1281), .B2(new_n1276), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1274), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1220), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1256), .A2(new_n1287), .A3(new_n1225), .A4(new_n1257), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1164), .A2(new_n702), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1197), .B1(new_n1289), .B2(new_n1163), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1226), .B(new_n1260), .C1(new_n1290), .C2(new_n1228), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1267), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1288), .A2(new_n1285), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1256), .A2(new_n1226), .A3(new_n1257), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1294), .B2(KEYINPUT62), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1273), .A2(new_n1286), .B1(new_n1293), .B2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(new_n1285), .A2(new_n1253), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1278), .A2(new_n1284), .A3(new_n1257), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1259), .A2(new_n1222), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1222), .A3(new_n1259), .A4(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(G402));
endmodule


