//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n217), .B1(new_n212), .B2(new_n211), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G226), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XNOR2_X1  g0043(.A(KEYINPUT3), .B(G33), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G223), .A3(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G222), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n245), .B1(new_n246), .B2(new_n244), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(G1), .B(G13), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n253), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n255), .B1(new_n260), .B2(G226), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n252), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT66), .B(G200), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT67), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  INV_X1    g0066(.A(new_n264), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n262), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n207), .A2(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n213), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n202), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n206), .B2(G20), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n202), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT9), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n263), .A2(G190), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n265), .A2(new_n268), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT10), .ZN(new_n285));
  INV_X1    g0085(.A(new_n281), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n262), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT65), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n263), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n289), .B2(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n244), .A2(G226), .A3(new_n247), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G97), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n244), .A2(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n230), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n251), .ZN(new_n298));
  INV_X1    g0098(.A(new_n255), .ZN(new_n299));
  INV_X1    g0099(.A(G238), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n259), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n301), .B1(new_n297), .B2(new_n251), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n303), .ZN(new_n306));
  OAI21_X1  g0106(.A(G169), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(KEYINPUT14), .B(G169), .C1(new_n304), .C2(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n298), .A2(new_n302), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n305), .A2(new_n303), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G179), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT70), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(new_n317), .A3(G179), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n269), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n272), .A2(new_n246), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n275), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g0124(.A(new_n324), .B(KEYINPUT11), .Z(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT69), .B1(new_n277), .B2(G68), .ZN(new_n326));
  XOR2_X1   g0126(.A(new_n326), .B(KEYINPUT12), .Z(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  INV_X1    g0128(.A(new_n279), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n320), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G200), .B1(new_n304), .B2(new_n306), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n313), .A2(G190), .A3(new_n314), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n331), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G20), .A2(G77), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n338), .B1(new_n271), .B2(new_n321), .C1(new_n272), .C2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(new_n275), .ZN(new_n341));
  INV_X1    g0141(.A(new_n277), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n246), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n329), .B2(new_n246), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G107), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n350), .B1(new_n296), .B2(new_n300), .C1(new_n230), .C2(new_n248), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n251), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n255), .B1(new_n260), .B2(G244), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n264), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n346), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n354), .A2(G169), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n345), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n293), .A2(new_n337), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n299), .B1(new_n259), .B2(new_n230), .ZN(new_n364));
  OAI211_X1 g0164(.A(G226), .B(G1698), .C1(new_n347), .C2(new_n348), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT72), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n244), .A2(KEYINPUT72), .A3(G226), .A4(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n244), .A2(G223), .A3(new_n247), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n364), .B1(new_n371), .B2(new_n251), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(G169), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n290), .B2(new_n372), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n271), .A2(new_n277), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n279), .B2(new_n271), .ZN(new_n376));
  INV_X1    g0176(.A(new_n275), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n244), .B2(G20), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n328), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G58), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n328), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n269), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT16), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n349), .B2(new_n207), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n347), .A2(new_n348), .A3(new_n378), .A4(G20), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(new_n386), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n377), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n376), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g0196(.A(KEYINPUT71), .B(new_n377), .C1(new_n387), .C2(new_n393), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n374), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT18), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n374), .B(new_n400), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n275), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n394), .A2(new_n395), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n372), .A2(new_n356), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G200), .B2(new_n372), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(new_n409), .A4(new_n376), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n376), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n405), .B2(KEYINPUT71), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT17), .A3(new_n407), .A4(new_n409), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT73), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n402), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n363), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n244), .A2(G257), .A3(G1698), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G294), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n244), .A2(G250), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n251), .ZN(new_n427));
  INV_X1    g0227(.A(G45), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G1), .ZN(new_n429));
  NOR2_X1   g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  AND2_X1   g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(G274), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT5), .B(G41), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n251), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G264), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT86), .B1(new_n436), .B2(G190), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(KEYINPUT86), .A3(new_n438), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT24), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT83), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT22), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT82), .ZN(new_n446));
  OR2_X1    g0246(.A1(KEYINPUT3), .A2(G33), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT3), .A2(G33), .ZN(new_n448));
  AOI21_X1  g0248(.A(G20), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n449), .B2(G87), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n207), .B(G87), .C1(new_n347), .C2(new_n348), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(KEYINPUT82), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n445), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(KEYINPUT82), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n244), .A2(new_n446), .A3(new_n207), .A4(G87), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT22), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  OR3_X1    g0257(.A1(new_n457), .A2(KEYINPUT84), .A3(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT85), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n207), .B2(G107), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT23), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT84), .B1(new_n272), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n459), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n458), .A2(new_n462), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AND4_X1   g0267(.A1(new_n444), .A2(new_n453), .A3(new_n456), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n454), .A2(new_n455), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n469), .B2(new_n445), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n444), .B1(new_n470), .B2(new_n456), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n443), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n453), .A2(new_n456), .A3(new_n467), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT83), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n444), .A3(new_n456), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(KEYINPUT24), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n275), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G13), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(G20), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n481), .A2(KEYINPUT25), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n206), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n277), .A2(new_n484), .A3(new_n213), .A4(new_n274), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n482), .B(new_n483), .C1(new_n480), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n442), .A2(new_n477), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n436), .A2(new_n290), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(G169), .B2(new_n436), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n477), .B2(new_n487), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n244), .A2(G264), .A3(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n349), .A2(G303), .ZN(new_n495));
  OAI211_X1 g0295(.A(G257), .B(new_n247), .C1(new_n347), .C2(new_n348), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n251), .ZN(new_n498));
  INV_X1    g0298(.A(new_n432), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n434), .B2(G270), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n493), .B(new_n287), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n500), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n290), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n207), .A2(new_n463), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G33), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n508), .B2(new_n207), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n504), .B1(new_n509), .B2(new_n377), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n256), .A2(G97), .ZN(new_n511));
  AOI21_X1  g0311(.A(G20), .B1(new_n511), .B2(new_n506), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT20), .B(new_n275), .C1(new_n512), .C2(new_n505), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n485), .A2(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n277), .A2(new_n463), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT78), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT78), .ZN(new_n519));
  AOI221_X4 g0319(.A(new_n519), .B1(new_n515), .B2(new_n516), .C1(new_n510), .C2(new_n513), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n501), .A2(new_n503), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT79), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI221_X1 g0323(.A(KEYINPUT79), .B1(new_n518), .B2(new_n520), .C1(new_n501), .C2(new_n503), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n287), .B1(new_n498), .B2(new_n500), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n520), .B2(new_n518), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n493), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n530), .A3(new_n493), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n520), .A2(new_n518), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n498), .A2(new_n500), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n438), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n520), .A2(new_n518), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n538), .B(KEYINPUT81), .C1(new_n438), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(G190), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n525), .A2(new_n532), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n543), .A2(new_n507), .A3(G107), .ZN(new_n544));
  XNOR2_X1  g0344(.A(G97), .B(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n546), .A2(new_n207), .B1(new_n246), .B2(new_n321), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n480), .B1(new_n379), .B2(new_n380), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n275), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n277), .A2(new_n507), .ZN(new_n550));
  INV_X1    g0350(.A(new_n485), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n507), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n247), .A2(KEYINPUT4), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n244), .A2(G244), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G244), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n349), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n506), .B(new_n555), .C1(new_n557), .C2(KEYINPUT4), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n247), .B1(new_n425), .B2(KEYINPUT4), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n251), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n499), .B1(new_n434), .B2(G257), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n433), .A2(new_n429), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G257), .A3(new_n258), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n432), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n553), .B1(new_n568), .B2(G179), .ZN(new_n569));
  AOI21_X1  g0369(.A(G169), .B1(new_n560), .B2(new_n561), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n560), .A2(G190), .A3(new_n561), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n549), .A3(new_n552), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n565), .A2(new_n562), .A3(new_n432), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n562), .B1(new_n565), .B2(new_n432), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n438), .B1(new_n575), .B2(new_n560), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n569), .A2(new_n570), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n207), .B1(new_n295), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n507), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n579), .B1(G107), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n244), .A2(new_n207), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(new_n328), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT76), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n578), .C1(new_n295), .C2(G20), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(new_n578), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n275), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n339), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n551), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n591), .B(new_n593), .C1(new_n277), .C2(new_n592), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n244), .A2(G238), .A3(new_n247), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n244), .A2(G244), .A3(G1698), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n457), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n251), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n206), .A2(G45), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n254), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n429), .A2(KEYINPUT75), .A3(G274), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n258), .A2(G250), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n290), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n251), .B2(new_n597), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n287), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n594), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n609), .A2(KEYINPUT77), .A3(G190), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT77), .B1(new_n609), .B2(G190), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI221_X1 g0414(.A(new_n582), .B1(new_n587), .B2(new_n589), .C1(new_n328), .C2(new_n583), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n275), .B1(new_n342), .B2(new_n339), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n551), .A2(G87), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n264), .C2(new_n609), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n611), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n577), .A2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n422), .A2(new_n492), .A3(new_n542), .A4(new_n620), .ZN(G372));
  NAND2_X1  g0421(.A1(new_n362), .A2(new_n336), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n418), .A2(new_n419), .B1(new_n333), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n285), .B1(new_n623), .B2(new_n402), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n292), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n560), .A2(new_n561), .ZN(new_n627));
  OAI221_X1 g0427(.A(new_n553), .B1(new_n568), .B2(G179), .C1(new_n627), .C2(G169), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n619), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n569), .A2(new_n570), .ZN(new_n630));
  INV_X1    g0430(.A(new_n613), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n609), .A2(KEYINPUT77), .A3(G190), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n591), .B(new_n617), .C1(new_n277), .C2(new_n592), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n267), .B2(new_n607), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n630), .A2(new_n636), .A3(new_n637), .A4(new_n611), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n611), .B(KEYINPUT87), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n442), .A2(new_n477), .A3(new_n487), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n532), .A2(new_n521), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n643), .B(new_n620), .C1(new_n644), .C2(new_n491), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n629), .A2(new_n638), .A3(new_n639), .A4(KEYINPUT88), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n626), .B1(new_n421), .B2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n479), .A2(new_n207), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n477), .B2(new_n487), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n488), .A2(new_n491), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n491), .A2(new_n655), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT89), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n657), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n477), .A2(new_n487), .ZN(new_n663));
  INV_X1    g0463(.A(new_n490), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n665), .A3(new_n643), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT89), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n659), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n538), .A2(new_n656), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n542), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n532), .A2(new_n521), .A3(new_n671), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G330), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n665), .A2(new_n655), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n655), .B1(new_n525), .B2(new_n532), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n669), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n581), .A2(G107), .A3(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n215), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n542), .A2(new_n492), .A3(new_n620), .A4(new_n656), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n535), .A2(G179), .A3(new_n609), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n436), .A3(new_n568), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n609), .A2(new_n435), .A3(new_n427), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n627), .A3(new_n503), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n692), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n655), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT31), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n688), .B1(new_n689), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n665), .A2(KEYINPUT91), .A3(new_n532), .A4(new_n525), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT91), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n527), .A2(new_n530), .A3(new_n493), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n530), .B1(new_n527), .B2(new_n493), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n523), .B(new_n524), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n701), .B1(new_n704), .B2(new_n491), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n620), .A2(new_n643), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n640), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT92), .B1(new_n709), .B2(new_n656), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n711), .B(new_n655), .C1(new_n707), .C2(new_n708), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT29), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n715), .B(KEYINPUT29), .C1(new_n710), .C2(new_n712), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n647), .A2(new_n656), .ZN(new_n718));
  XOR2_X1   g0518(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n699), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n687), .B1(new_n721), .B2(G1), .ZN(G364));
  NAND3_X1  g0522(.A1(new_n207), .A2(G13), .A3(G45), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n683), .A2(G1), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n672), .A2(new_n673), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n478), .A2(new_n256), .A3(KEYINPUT95), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G13), .B2(G33), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT101), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n681), .A2(new_n349), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G355), .B1(new_n463), .B2(new_n681), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n210), .A2(new_n349), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT94), .Z(new_n738));
  NOR2_X1   g0538(.A1(new_n216), .A2(G45), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n242), .B2(G45), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n736), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n213), .B1(G20), .B2(new_n287), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n207), .A2(new_n356), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n746), .A2(new_n290), .A3(G200), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n349), .B1(new_n747), .B2(G58), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n207), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT98), .B(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n753), .A2(new_n754), .B1(G97), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n748), .B(new_n757), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  INV_X1    g0558(.A(new_n749), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n264), .A2(new_n759), .A3(G179), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n480), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n759), .A2(new_n290), .A3(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT96), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n763), .A2(KEYINPUT96), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n762), .B1(new_n768), .B2(G77), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n746), .A2(new_n264), .A3(G179), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n769), .B1(new_n580), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(G190), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n758), .B(new_n772), .C1(G50), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n774), .A2(new_n356), .A3(new_n775), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT100), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT100), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G68), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n751), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n763), .A2(G311), .B1(G329), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  INV_X1    g0588(.A(new_n747), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n349), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n771), .B1(new_n761), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n776), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n756), .ZN(new_n796));
  INV_X1    g0596(.A(G294), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n790), .A2(new_n793), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n778), .A2(new_n783), .B1(new_n785), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n742), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n744), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n725), .B1(new_n734), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n674), .ZN(new_n804));
  AOI21_X1  g0604(.A(G330), .B1(new_n672), .B2(new_n673), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n724), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT102), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n362), .A2(new_n656), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n345), .A2(new_n656), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n359), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(new_n811), .B2(new_n362), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n718), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n725), .B1(new_n814), .B2(new_n699), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n699), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n730), .A2(new_n742), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n724), .B1(new_n246), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT103), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n349), .B1(new_n789), .B2(new_n797), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G311), .B2(new_n786), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n507), .B2(new_n796), .C1(new_n791), .C2(new_n776), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n768), .A2(G116), .B1(G107), .B2(new_n770), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n580), .B2(new_n761), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(G283), .C2(new_n782), .ZN(new_n825));
  INV_X1    g0625(.A(new_n752), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n768), .A2(new_n826), .B1(G143), .B2(new_n747), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  INV_X1    g0629(.A(new_n782), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n827), .B1(new_n828), .B2(new_n776), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n760), .A2(G68), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n770), .A2(G50), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n756), .A2(G58), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n349), .B1(new_n786), .B2(G132), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n825), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n819), .B1(new_n813), .B2(new_n731), .C1(new_n838), .C2(new_n801), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n816), .A2(new_n839), .ZN(G384));
  INV_X1    g0640(.A(new_n720), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n714), .B2(new_n716), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n625), .B1(new_n842), .B2(new_n422), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n333), .A2(new_n655), .ZN(new_n844));
  INV_X1    g0644(.A(new_n410), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n394), .A2(new_n413), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n372), .A2(new_n290), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(G169), .B2(new_n372), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n848), .B2(new_n653), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT37), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n653), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n396), .B2(new_n397), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n398), .A2(new_n852), .A3(new_n853), .A4(new_n410), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n846), .A2(new_n653), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n420), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT38), .B(new_n855), .C1(new_n420), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n398), .A2(new_n852), .A3(new_n410), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT106), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n854), .ZN(new_n866));
  INV_X1    g0666(.A(new_n852), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n402), .B2(new_n416), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n865), .B1(new_n864), .B2(new_n854), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n859), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n861), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n862), .A2(KEYINPUT39), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(KEYINPUT105), .B(new_n872), .C1(new_n860), .C2(new_n861), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n844), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n647), .A2(new_n656), .A3(new_n813), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n809), .ZN(new_n879));
  INV_X1    g0679(.A(new_n336), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n332), .B(new_n655), .C1(new_n320), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n332), .A2(new_n655), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n309), .A2(new_n310), .B1(new_n316), .B2(new_n318), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n336), .B(new_n882), .C1(new_n883), .C2(new_n331), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n887), .A2(new_n862), .B1(new_n402), .B2(new_n653), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n877), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n843), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n885), .A2(new_n813), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n689), .B2(new_n698), .ZN(new_n892));
  INV_X1    g0692(.A(new_n861), .ZN(new_n893));
  INV_X1    g0693(.A(new_n402), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n415), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT73), .B1(new_n412), .B2(new_n415), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n856), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n898), .B2(new_n855), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n892), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n871), .A2(new_n861), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n689), .A2(new_n698), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n812), .B1(new_n881), .B2(new_n884), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n900), .A2(new_n901), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n422), .A2(new_n903), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n907), .B(new_n908), .Z(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(new_n688), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n890), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT107), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n890), .A2(new_n910), .ZN(new_n915));
  OAI21_X1  g0715(.A(G1), .B1(new_n478), .B2(G20), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(G77), .B1(new_n382), .B2(new_n328), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n918), .A2(new_n215), .B1(G50), .B2(new_n328), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G1), .A3(new_n478), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n214), .A2(G116), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n546), .B(KEYINPUT104), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT35), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT36), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n925), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n917), .A2(new_n928), .ZN(G367));
  NOR3_X1   g0729(.A1(new_n658), .A2(new_n660), .A3(KEYINPUT89), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n667), .B1(new_n666), .B2(new_n659), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n678), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n656), .B1(new_n549), .B2(new_n552), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n577), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n630), .A2(new_n655), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n628), .B1(new_n935), .B2(new_n665), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n656), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n938), .B2(KEYINPUT42), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT43), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n634), .A2(new_n655), .ZN(new_n944));
  MUX2_X1   g0744(.A(new_n639), .B(new_n619), .S(new_n944), .Z(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT108), .Z(new_n946));
  OAI22_X1  g0746(.A1(new_n939), .A2(new_n942), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n943), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n675), .A2(new_n937), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n682), .B(KEYINPUT41), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n717), .A2(new_n720), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n674), .A2(KEYINPUT110), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n669), .A2(new_n678), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n954), .A2(new_n933), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n954), .B1(new_n933), .B2(new_n955), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n699), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT111), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n679), .B2(new_n937), .ZN(new_n964));
  INV_X1    g0764(.A(new_n677), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n932), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n937), .ZN(new_n967));
  INV_X1    g0767(.A(new_n963), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n964), .A2(new_n969), .B1(KEYINPUT109), .B2(new_n962), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT45), .B1(new_n679), .B2(new_n937), .ZN(new_n971));
  AND4_X1   g0771(.A1(KEYINPUT45), .A2(new_n932), .A3(new_n965), .A4(new_n937), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n675), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n679), .A2(new_n937), .A3(new_n963), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n971), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n937), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n981), .A3(new_n676), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n974), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT111), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n721), .A2(new_n984), .A3(new_n958), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n961), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n952), .B1(new_n986), .B2(new_n721), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n723), .A2(G1), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n951), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n946), .A2(new_n733), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n770), .A2(G116), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT46), .Z(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n349), .B1(new_n751), .B2(new_n993), .C1(new_n789), .C2(new_n791), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G107), .B2(new_n756), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n768), .A2(G283), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n777), .A2(G311), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n760), .A2(G97), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n992), .B(new_n999), .C1(G294), .C2(new_n782), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n244), .B1(new_n751), .B2(new_n828), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n770), .B2(G58), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n246), .B2(new_n761), .C1(new_n767), .C2(new_n202), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n756), .A2(G68), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n789), .B2(new_n829), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g0807(.A(G143), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n776), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1003), .B(new_n1009), .C1(new_n782), .C2(new_n826), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1000), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n801), .B1(new_n1011), .B2(KEYINPUT47), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT47), .B2(new_n1011), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n743), .B1(new_n210), .B2(new_n339), .C1(new_n738), .C2(new_n234), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n990), .A2(new_n725), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n989), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n956), .A2(new_n957), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n988), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT113), .Z(new_n1020));
  INV_X1    g0820(.A(new_n684), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n735), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(G107), .B2(new_n210), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n231), .A2(G45), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n271), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n202), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT50), .Z(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1021), .C1(G68), .C2(G77), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n738), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1023), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n743), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n725), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT114), .Z(new_n1033));
  INV_X1    g0833(.A(G159), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n776), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n763), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n789), .A2(new_n202), .B1(new_n1036), .B2(new_n328), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n349), .B(new_n1037), .C1(G150), .C2(new_n786), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n592), .A2(new_n756), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n770), .A2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1038), .A2(new_n998), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1035), .B(new_n1041), .C1(new_n1025), .C2(new_n782), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n768), .A2(G303), .B1(G317), .B2(new_n747), .ZN(new_n1043));
  INV_X1    g0843(.A(G311), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n788), .B2(new_n776), .C1(new_n1044), .C2(new_n830), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT48), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(KEYINPUT48), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n770), .A2(G294), .B1(G283), .B2(new_n756), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n349), .B1(new_n794), .B2(new_n751), .C1(new_n761), .C2(new_n463), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1042), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1033), .B1(new_n1055), .B2(new_n801), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n670), .B2(new_n733), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1020), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n984), .B1(new_n721), .B2(new_n958), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n842), .A2(new_n1017), .A3(KEYINPUT111), .A4(new_n699), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n682), .B1(new_n721), .B2(new_n958), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n983), .A2(new_n988), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n738), .A2(new_n239), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n743), .B1(new_n507), .B2(new_n210), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n725), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n768), .A2(new_n1025), .B1(G68), .B2(new_n770), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n789), .A2(new_n1034), .B1(new_n829), .B2(new_n776), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n782), .A2(G50), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n244), .B1(new_n751), .B2(new_n1008), .C1(new_n796), .C2(new_n246), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G87), .B2(new_n760), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n244), .B1(new_n786), .B2(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n463), .B2(new_n796), .C1(new_n1036), .C2(new_n797), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n762), .B(new_n1075), .C1(G283), .C2(new_n770), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n791), .B2(new_n830), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n777), .A2(G317), .B1(G311), .B2(new_n747), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1066), .B1(new_n1080), .B2(new_n742), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n732), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n937), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n683), .B1(new_n1085), .B2(new_n983), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n983), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(G390));
  NAND2_X1  g0890(.A1(new_n873), .A2(new_n874), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT39), .B1(new_n893), .B2(new_n899), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n862), .A2(new_n874), .A3(KEYINPUT39), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n730), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n817), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n725), .B1(new_n1025), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n776), .A2(new_n792), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n747), .A2(G116), .B1(G294), .B2(new_n786), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n833), .C1(new_n246), .C2(new_n796), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G97), .C2(new_n768), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n244), .B1(new_n770), .B2(G87), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n480), .C2(new_n830), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT118), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n349), .B1(new_n786), .B2(G125), .ZN(new_n1108));
  INV_X1    g0908(.A(G132), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n789), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n767), .A2(new_n1111), .B1(new_n202), .B2(new_n761), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(G159), .C2(new_n756), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n782), .A2(G137), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n770), .A2(G150), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT53), .Z(new_n1116));
  NAND2_X1  g0916(.A1(new_n777), .A2(G128), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1106), .A2(new_n1107), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1097), .B1(new_n1119), .B2(new_n742), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1095), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n699), .A2(new_n904), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n844), .B1(new_n879), .B2(new_n885), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n875), .A2(new_n876), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n844), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n902), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n811), .A2(new_n362), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n710), .B2(new_n712), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n809), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1127), .B1(new_n1131), .B2(new_n885), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1123), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n886), .A2(new_n1126), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1093), .A2(new_n1134), .A3(new_n1094), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n885), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1130), .B2(new_n809), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1122), .C1(new_n1137), .C2(new_n1127), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1121), .B1(new_n1139), .B2(new_n1018), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n717), .A2(new_n422), .A3(new_n720), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n422), .A2(G330), .A3(new_n903), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n699), .A2(new_n813), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1136), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n879), .B1(new_n1145), .B2(new_n1122), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1123), .B1(new_n1136), .B2(new_n1144), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1131), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1142), .A2(new_n626), .A3(new_n1143), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT116), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT116), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n843), .A2(new_n1151), .A3(new_n1143), .A4(new_n1148), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1150), .A2(new_n1139), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n682), .B1(new_n1139), .B2(new_n1149), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1141), .B1(new_n1153), .B2(new_n1154), .ZN(G378));
  NAND3_X1  g0955(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n892), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n903), .A2(new_n904), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n860), .B2(new_n861), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1156), .B(G330), .C1(new_n1158), .C2(KEYINPUT40), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n286), .B(new_n653), .C1(new_n285), .C2(new_n292), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n286), .A2(new_n653), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n293), .A2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  OR3_X1    g0963(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(KEYINPUT121), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n900), .A2(new_n901), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1169), .A2(G330), .A3(new_n1156), .A4(new_n1166), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n877), .A2(new_n1168), .A3(new_n888), .A4(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1170), .A2(new_n1168), .B1(new_n877), .B2(new_n888), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT122), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n889), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT122), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1168), .A2(new_n877), .A3(new_n1170), .A4(new_n888), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1142), .A2(new_n626), .A3(new_n1143), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1148), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1139), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n682), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1164), .A2(new_n730), .A3(new_n1165), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n725), .B1(G50), .B2(new_n1096), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n349), .A2(new_n257), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n789), .A2(new_n480), .B1(new_n1036), .B2(new_n339), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(G283), .C2(new_n786), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n760), .A2(G58), .ZN(new_n1196));
  AND4_X1   g0996(.A1(new_n1004), .A2(new_n1195), .A3(new_n1040), .A4(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n507), .B2(new_n830), .C1(new_n463), .C2(new_n776), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1199));
  OAI21_X1  g0999(.A(new_n1193), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1199), .B2(new_n1198), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n747), .A2(G128), .B1(G150), .B2(new_n756), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n777), .A2(G125), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n771), .C2(new_n1111), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n782), .A2(G132), .B1(G137), .B2(new_n763), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT120), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT120), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT59), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n761), .B2(new_n752), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1201), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1191), .B1(new_n1213), .B2(new_n742), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1190), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1179), .B2(new_n988), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1189), .A2(new_n1217), .ZN(G375));
  AOI21_X1  g1018(.A(new_n952), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n724), .B1(new_n328), .B2(new_n817), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT123), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n349), .B1(new_n751), .B2(new_n791), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n767), .A2(new_n480), .B1(new_n507), .B2(new_n771), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G77), .C2(new_n760), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1039), .B1(new_n789), .B2(new_n792), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT124), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1226), .A2(new_n1227), .B1(new_n797), .B2(new_n776), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1227), .B2(new_n1226), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1225), .B(new_n1229), .C1(new_n463), .C2(new_n830), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1196), .B1(new_n771), .B2(new_n1034), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n244), .B1(new_n789), .B2(new_n828), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n786), .A2(G128), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1036), .B2(new_n829), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n796), .A2(new_n202), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n1109), .B2(new_n776), .C1(new_n830), .C2(new_n1111), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1222), .B1(new_n1238), .B2(new_n801), .C1(new_n885), .C2(new_n731), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1182), .B2(new_n1018), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1220), .A2(new_n1241), .ZN(G381));
  INV_X1    g1042(.A(new_n1154), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1150), .A2(new_n1139), .A3(new_n1152), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1140), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1189), .A2(new_n1245), .A3(new_n1217), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n989), .A2(new_n1015), .A3(new_n1089), .ZN(new_n1247));
  INV_X1    g1047(.A(G396), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1058), .A2(new_n1248), .A3(new_n1061), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(G384), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G381), .A2(new_n1246), .A3(new_n1247), .A4(new_n1250), .ZN(G407));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G343), .C2(new_n1246), .ZN(G409));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1249), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1247), .A2(KEYINPUT127), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1089), .B1(new_n989), .B2(new_n1015), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(KEYINPUT127), .A3(new_n1247), .A4(new_n1254), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1217), .C1(new_n1184), .C2(new_n1188), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n952), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1179), .A2(new_n1263), .A3(new_n1183), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1216), .B1(new_n1265), .B2(new_n988), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1245), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(KEYINPUT60), .B(new_n1148), .C1(new_n843), .C2(new_n1143), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n682), .B(new_n1149), .C1(new_n1270), .C2(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1273), .A2(new_n1241), .A3(G384), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1273), .B2(new_n1241), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n654), .A2(G213), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1269), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1262), .A2(new_n1268), .B1(G213), .B2(new_n654), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(KEYINPUT125), .A3(new_n1276), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT62), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1269), .A2(new_n1277), .ZN(new_n1284));
  INV_X1    g1084(.A(G2897), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1274), .A2(new_n1275), .B1(new_n1285), .B2(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1273), .A2(new_n1241), .ZN(new_n1287));
  INV_X1    g1087(.A(G384), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1273), .A2(new_n1241), .A3(G384), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1277), .A2(new_n1285), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(KEYINPUT62), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1261), .B1(new_n1283), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1299));
  AND4_X1   g1099(.A1(new_n1298), .A2(new_n1258), .A3(new_n1299), .A4(new_n1260), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1281), .A2(KEYINPUT126), .B1(new_n1292), .B2(new_n1286), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(KEYINPUT126), .B2(new_n1281), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1280), .A2(new_n1303), .A3(new_n1282), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1297), .A2(new_n1305), .ZN(G405));
  AND3_X1   g1106(.A1(new_n1258), .A2(new_n1260), .A3(new_n1276), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1276), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1246), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1245), .B1(new_n1189), .B2(new_n1217), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n1307), .A2(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1276), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1261), .A2(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1258), .A2(new_n1260), .A3(new_n1276), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1311), .A2(new_n1316), .ZN(G402));
endmodule


