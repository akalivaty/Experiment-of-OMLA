

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(G2105), .A2(n529), .ZN(n700) );
  BUF_X1 U556 ( .A(n697), .Z(n624) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n532), .Z(n697) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n533), .ZN(n899) );
  INV_X1 U559 ( .A(G2105), .ZN(n533) );
  XNOR2_X1 U560 ( .A(n522), .B(n772), .ZN(n521) );
  AND2_X1 U561 ( .A1(n771), .A2(G8), .ZN(n522) );
  NOR2_X2 U562 ( .A1(n758), .A2(G2084), .ZN(n775) );
  BUF_X4 U563 ( .A(n733), .Z(n758) );
  OR2_X1 U564 ( .A1(n988), .A2(n739), .ZN(n747) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n753) );
  XNOR2_X1 U566 ( .A(n725), .B(KEYINPUT31), .ZN(n774) );
  INV_X1 U567 ( .A(KEYINPUT108), .ZN(n791) );
  NAND2_X1 U568 ( .A1(n790), .A2(n789), .ZN(n792) );
  NOR2_X2 U569 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  BUF_X2 U570 ( .A(n620), .Z(n898) );
  AND2_X1 U571 ( .A1(n777), .A2(n717), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n712), .A2(n784), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n796), .A2(n783), .ZN(n790) );
  NAND2_X1 U574 ( .A1(n521), .A2(n527), .ZN(n796) );
  NOR2_X2 U575 ( .A1(n741), .A2(n989), .ZN(n740) );
  NOR2_X2 U576 ( .A1(n706), .A2(n705), .ZN(G160) );
  XNOR2_X1 U577 ( .A(n565), .B(KEYINPUT13), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n782), .A2(n781), .ZN(n526) );
  OR2_X1 U579 ( .A1(n779), .A2(n778), .ZN(n527) );
  INV_X1 U580 ( .A(KEYINPUT26), .ZN(n734) );
  INV_X1 U581 ( .A(G8), .ZN(n716) );
  NOR2_X1 U582 ( .A1(n997), .A2(n748), .ZN(n732) );
  INV_X1 U583 ( .A(KEYINPUT96), .ZN(n713) );
  INV_X1 U584 ( .A(KEYINPUT104), .ZN(n769) );
  XNOR2_X1 U585 ( .A(n709), .B(KEYINPUT64), .ZN(n715) );
  INV_X1 U586 ( .A(KEYINPUT109), .ZN(n800) );
  NOR2_X1 U587 ( .A1(G164), .A2(G1384), .ZN(n805) );
  NOR2_X2 U588 ( .A1(n644), .A2(n541), .ZN(n662) );
  NOR2_X1 U589 ( .A1(n529), .A2(n533), .ZN(n620) );
  BUF_X1 U590 ( .A(n700), .Z(n901) );
  NOR2_X1 U591 ( .A1(G651), .A2(n644), .ZN(n659) );
  XOR2_X1 U592 ( .A(KEYINPUT72), .B(n571), .Z(n1005) );
  INV_X1 U593 ( .A(G2104), .ZN(n529) );
  NAND2_X1 U594 ( .A1(n620), .A2(G114), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n528), .B(KEYINPUT90), .ZN(n531) );
  NAND2_X1 U596 ( .A1(G102), .A2(n901), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n537) );
  NAND2_X1 U598 ( .A1(G138), .A2(n697), .ZN(n535) );
  NAND2_X1 U599 ( .A1(G126), .A2(n899), .ZN(n534) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(G164) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT65), .B(n538), .Z(n561) );
  BUF_X1 U604 ( .A(n561), .Z(n658) );
  NAND2_X1 U605 ( .A1(G88), .A2(n658), .ZN(n540) );
  XOR2_X1 U606 ( .A(G543), .B(KEYINPUT0), .Z(n644) );
  INV_X1 U607 ( .A(G651), .ZN(n541) );
  NAND2_X1 U608 ( .A1(G75), .A2(n662), .ZN(n539) );
  NAND2_X1 U609 ( .A1(n540), .A2(n539), .ZN(n549) );
  NOR2_X1 U610 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U611 ( .A(KEYINPUT68), .B(n542), .Z(n543) );
  XNOR2_X1 U612 ( .A(KEYINPUT1), .B(n543), .ZN(n567) );
  BUF_X1 U613 ( .A(n567), .Z(n667) );
  NAND2_X1 U614 ( .A1(G62), .A2(n667), .ZN(n544) );
  XNOR2_X1 U615 ( .A(n544), .B(KEYINPUT84), .ZN(n546) );
  NAND2_X1 U616 ( .A1(G50), .A2(n659), .ZN(n545) );
  NAND2_X1 U617 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U618 ( .A(KEYINPUT85), .B(n547), .Z(n548) );
  NOR2_X1 U619 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U620 ( .A(KEYINPUT86), .B(n550), .Z(G303) );
  INV_X1 U621 ( .A(G303), .ZN(G166) );
  XOR2_X1 U622 ( .A(KEYINPUT111), .B(G2435), .Z(n552) );
  XNOR2_X1 U623 ( .A(G2430), .B(G2438), .ZN(n551) );
  XNOR2_X1 U624 ( .A(n552), .B(n551), .ZN(n559) );
  XOR2_X1 U625 ( .A(G2446), .B(G2454), .Z(n554) );
  XNOR2_X1 U626 ( .A(G2451), .B(G2443), .ZN(n553) );
  XNOR2_X1 U627 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U628 ( .A(n555), .B(G2427), .Z(n557) );
  XNOR2_X1 U629 ( .A(G1348), .B(G1341), .ZN(n556) );
  XNOR2_X1 U630 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U631 ( .A(n559), .B(n558), .ZN(n560) );
  AND2_X1 U632 ( .A1(n560), .A2(G14), .ZN(G401) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U634 ( .A(G860), .ZN(n613) );
  NAND2_X1 U635 ( .A1(n561), .A2(G81), .ZN(n562) );
  XNOR2_X1 U636 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U637 ( .A1(G68), .A2(n662), .ZN(n563) );
  NAND2_X1 U638 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G43), .A2(n659), .ZN(n566) );
  NAND2_X1 U640 ( .A1(n525), .A2(n566), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n567), .A2(G56), .ZN(n568) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n568), .Z(n569) );
  NOR2_X1 U643 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U644 ( .A1(n613), .A2(n1005), .ZN(G153) );
  INV_X1 U645 ( .A(G82), .ZN(G220) );
  INV_X1 U646 ( .A(G57), .ZN(G237) );
  INV_X1 U647 ( .A(G120), .ZN(G236) );
  NAND2_X1 U648 ( .A1(G52), .A2(n659), .ZN(n573) );
  NAND2_X1 U649 ( .A1(G64), .A2(n667), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G90), .A2(n658), .ZN(n575) );
  NAND2_X1 U652 ( .A1(G77), .A2(n662), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U654 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U655 ( .A1(n578), .A2(n577), .ZN(G171) );
  NAND2_X1 U656 ( .A1(n658), .A2(G89), .ZN(n579) );
  XNOR2_X1 U657 ( .A(KEYINPUT4), .B(n579), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n662), .A2(G76), .ZN(n580) );
  XOR2_X1 U659 ( .A(KEYINPUT73), .B(n580), .Z(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U661 ( .A(n583), .B(KEYINPUT5), .ZN(n590) );
  XNOR2_X1 U662 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n588) );
  NAND2_X1 U663 ( .A1(G63), .A2(n667), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n584), .B(KEYINPUT74), .ZN(n586) );
  NAND2_X1 U665 ( .A1(G51), .A2(n659), .ZN(n585) );
  NAND2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U667 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U669 ( .A(KEYINPUT7), .B(n591), .ZN(G168) );
  XOR2_X1 U670 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U671 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n592), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U673 ( .A(G223), .ZN(n855) );
  NAND2_X1 U674 ( .A1(n855), .A2(G567), .ZN(n593) );
  XOR2_X1 U675 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  INV_X1 U676 ( .A(G171), .ZN(G301) );
  NAND2_X1 U677 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G92), .A2(n658), .ZN(n595) );
  NAND2_X1 U679 ( .A1(G79), .A2(n662), .ZN(n594) );
  NAND2_X1 U680 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U681 ( .A1(G54), .A2(n659), .ZN(n597) );
  NAND2_X1 U682 ( .A1(G66), .A2(n667), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U685 ( .A(KEYINPUT15), .B(n600), .Z(n988) );
  INV_X1 U686 ( .A(n988), .ZN(n924) );
  INV_X1 U687 ( .A(G868), .ZN(n679) );
  NAND2_X1 U688 ( .A1(n924), .A2(n679), .ZN(n601) );
  NAND2_X1 U689 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U690 ( .A1(G53), .A2(n659), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n603), .B(KEYINPUT70), .ZN(n610) );
  NAND2_X1 U692 ( .A1(G91), .A2(n658), .ZN(n605) );
  NAND2_X1 U693 ( .A1(G65), .A2(n667), .ZN(n604) );
  NAND2_X1 U694 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U695 ( .A1(G78), .A2(n662), .ZN(n606) );
  XNOR2_X1 U696 ( .A(KEYINPUT69), .B(n606), .ZN(n607) );
  NOR2_X1 U697 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U698 ( .A1(n610), .A2(n609), .ZN(G299) );
  NOR2_X1 U699 ( .A1(G286), .A2(n679), .ZN(n612) );
  NOR2_X1 U700 ( .A1(G868), .A2(G299), .ZN(n611) );
  NOR2_X1 U701 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U702 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n614), .A2(n988), .ZN(n615) );
  XNOR2_X1 U704 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U705 ( .A1(n924), .A2(n679), .ZN(n616) );
  XOR2_X1 U706 ( .A(KEYINPUT76), .B(n616), .Z(n617) );
  NOR2_X1 U707 ( .A1(G559), .A2(n617), .ZN(n619) );
  NOR2_X1 U708 ( .A1(n1005), .A2(G868), .ZN(n618) );
  NOR2_X1 U709 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U710 ( .A1(G111), .A2(n898), .ZN(n622) );
  NAND2_X1 U711 ( .A1(G99), .A2(n901), .ZN(n621) );
  NAND2_X1 U712 ( .A1(n622), .A2(n621), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n899), .A2(G123), .ZN(n623) );
  XNOR2_X1 U714 ( .A(n623), .B(KEYINPUT18), .ZN(n626) );
  NAND2_X1 U715 ( .A1(G135), .A2(n624), .ZN(n625) );
  NAND2_X1 U716 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U717 ( .A(KEYINPUT77), .B(n627), .Z(n628) );
  NOR2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n937) );
  XOR2_X1 U719 ( .A(G2096), .B(n937), .Z(n630) );
  NOR2_X1 U720 ( .A1(G2100), .A2(n630), .ZN(n631) );
  XOR2_X1 U721 ( .A(KEYINPUT78), .B(n631), .Z(G156) );
  NAND2_X1 U722 ( .A1(G93), .A2(n658), .ZN(n633) );
  NAND2_X1 U723 ( .A1(G80), .A2(n662), .ZN(n632) );
  NAND2_X1 U724 ( .A1(n633), .A2(n632), .ZN(n639) );
  NAND2_X1 U725 ( .A1(G55), .A2(n659), .ZN(n634) );
  XNOR2_X1 U726 ( .A(n634), .B(KEYINPUT82), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n667), .A2(G67), .ZN(n635) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(n635), .Z(n636) );
  NAND2_X1 U729 ( .A1(n637), .A2(n636), .ZN(n638) );
  OR2_X1 U730 ( .A1(n639), .A2(n638), .ZN(n678) );
  NAND2_X1 U731 ( .A1(n988), .A2(G559), .ZN(n676) );
  XOR2_X1 U732 ( .A(n1005), .B(KEYINPUT79), .Z(n640) );
  XNOR2_X1 U733 ( .A(n676), .B(n640), .ZN(n641) );
  NOR2_X1 U734 ( .A1(G860), .A2(n641), .ZN(n642) );
  XNOR2_X1 U735 ( .A(n642), .B(KEYINPUT80), .ZN(n643) );
  XOR2_X1 U736 ( .A(n678), .B(n643), .Z(G145) );
  NAND2_X1 U737 ( .A1(G87), .A2(n644), .ZN(n646) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U739 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U740 ( .A1(n667), .A2(n647), .ZN(n649) );
  NAND2_X1 U741 ( .A1(n659), .A2(G49), .ZN(n648) );
  NAND2_X1 U742 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U743 ( .A1(n658), .A2(G85), .ZN(n650) );
  XNOR2_X1 U744 ( .A(n650), .B(KEYINPUT66), .ZN(n652) );
  NAND2_X1 U745 ( .A1(G72), .A2(n662), .ZN(n651) );
  NAND2_X1 U746 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U747 ( .A(KEYINPUT67), .B(n653), .ZN(n657) );
  NAND2_X1 U748 ( .A1(n667), .A2(G60), .ZN(n655) );
  NAND2_X1 U749 ( .A1(G47), .A2(n659), .ZN(n654) );
  AND2_X1 U750 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U751 ( .A1(n657), .A2(n656), .ZN(G290) );
  NAND2_X1 U752 ( .A1(G86), .A2(n658), .ZN(n661) );
  NAND2_X1 U753 ( .A1(G48), .A2(n659), .ZN(n660) );
  NAND2_X1 U754 ( .A1(n661), .A2(n660), .ZN(n666) );
  NAND2_X1 U755 ( .A1(G73), .A2(n662), .ZN(n663) );
  XNOR2_X1 U756 ( .A(n663), .B(KEYINPUT2), .ZN(n664) );
  XNOR2_X1 U757 ( .A(n664), .B(KEYINPUT83), .ZN(n665) );
  NOR2_X1 U758 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U759 ( .A1(G61), .A2(n667), .ZN(n668) );
  NAND2_X1 U760 ( .A1(n669), .A2(n668), .ZN(G305) );
  XOR2_X1 U761 ( .A(n678), .B(KEYINPUT19), .Z(n671) );
  INV_X1 U762 ( .A(G299), .ZN(n997) );
  XNOR2_X1 U763 ( .A(G288), .B(n997), .ZN(n670) );
  XNOR2_X1 U764 ( .A(n671), .B(n670), .ZN(n674) );
  XNOR2_X1 U765 ( .A(n1005), .B(G290), .ZN(n672) );
  XNOR2_X1 U766 ( .A(n672), .B(G166), .ZN(n673) );
  XNOR2_X1 U767 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U768 ( .A(n675), .B(G305), .ZN(n921) );
  XNOR2_X1 U769 ( .A(n676), .B(n921), .ZN(n677) );
  NAND2_X1 U770 ( .A1(n677), .A2(G868), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U773 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U774 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U775 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U776 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U777 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U778 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  XNOR2_X1 U779 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U780 ( .A1(G236), .A2(G237), .ZN(n686) );
  NAND2_X1 U781 ( .A1(G69), .A2(n686), .ZN(n687) );
  XNOR2_X1 U782 ( .A(KEYINPUT89), .B(n687), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n688), .A2(G108), .ZN(n860) );
  NAND2_X1 U784 ( .A1(n860), .A2(G567), .ZN(n695) );
  NOR2_X1 U785 ( .A1(G220), .A2(G219), .ZN(n690) );
  XNOR2_X1 U786 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n689) );
  XNOR2_X1 U787 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n691), .A2(G218), .ZN(n692) );
  XNOR2_X1 U789 ( .A(KEYINPUT88), .B(n692), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n693), .A2(G96), .ZN(n861) );
  NAND2_X1 U791 ( .A1(n861), .A2(G2106), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n862) );
  NAND2_X1 U793 ( .A1(G483), .A2(G661), .ZN(n696) );
  NOR2_X1 U794 ( .A1(n862), .A2(n696), .ZN(n859) );
  NAND2_X1 U795 ( .A1(n859), .A2(G36), .ZN(G176) );
  NAND2_X1 U796 ( .A1(G125), .A2(n899), .ZN(n699) );
  NAND2_X1 U797 ( .A1(G137), .A2(n697), .ZN(n698) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n706) );
  NAND2_X1 U799 ( .A1(G101), .A2(n700), .ZN(n702) );
  INV_X1 U800 ( .A(KEYINPUT23), .ZN(n701) );
  XNOR2_X1 U801 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n898), .A2(G113), .ZN(n703) );
  NAND2_X1 U803 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U804 ( .A1(G160), .A2(G40), .ZN(n804) );
  XNOR2_X1 U805 ( .A(n804), .B(KEYINPUT95), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n708), .A2(n805), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n715), .A2(G8), .ZN(n712) );
  NOR2_X1 U808 ( .A1(G1981), .A2(G305), .ZN(n710) );
  XOR2_X1 U809 ( .A(n710), .B(KEYINPUT24), .Z(n711) );
  NOR2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n803) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n712), .ZN(n714) );
  XNOR2_X1 U812 ( .A(n714), .B(n713), .ZN(n777) );
  INV_X1 U813 ( .A(n715), .ZN(n726) );
  INV_X1 U814 ( .A(n726), .ZN(n733) );
  NOR2_X1 U815 ( .A1(n775), .A2(n716), .ZN(n717) );
  XOR2_X1 U816 ( .A(KEYINPUT30), .B(n523), .Z(n718) );
  NOR2_X1 U817 ( .A1(G168), .A2(n718), .ZN(n719) );
  XNOR2_X1 U818 ( .A(n719), .B(KEYINPUT101), .ZN(n724) );
  INV_X1 U819 ( .A(n758), .ZN(n741) );
  NOR2_X1 U820 ( .A1(G1961), .A2(n741), .ZN(n721) );
  XOR2_X1 U821 ( .A(KEYINPUT25), .B(G2078), .Z(n966) );
  NOR2_X1 U822 ( .A1(n758), .A2(n966), .ZN(n720) );
  NOR2_X1 U823 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U824 ( .A(KEYINPUT97), .B(n722), .ZN(n755) );
  OR2_X1 U825 ( .A1(n755), .A2(G171), .ZN(n723) );
  NAND2_X1 U826 ( .A1(n724), .A2(n723), .ZN(n725) );
  AND2_X1 U827 ( .A1(n726), .A2(G2072), .ZN(n728) );
  XNOR2_X1 U828 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n727) );
  XNOR2_X1 U829 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U830 ( .A1(n758), .A2(G1956), .ZN(n729) );
  NAND2_X1 U831 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U832 ( .A(KEYINPUT99), .B(n731), .ZN(n748) );
  XOR2_X1 U833 ( .A(n732), .B(KEYINPUT28), .Z(n752) );
  INV_X1 U834 ( .A(G1996), .ZN(n961) );
  NOR2_X1 U835 ( .A1(n733), .A2(n961), .ZN(n735) );
  XNOR2_X1 U836 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U837 ( .A1(n758), .A2(G1341), .ZN(n736) );
  NAND2_X1 U838 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U839 ( .A1(n1005), .A2(n738), .ZN(n739) );
  NAND2_X1 U840 ( .A1(n988), .A2(n739), .ZN(n745) );
  INV_X1 U841 ( .A(G1348), .ZN(n989) );
  XOR2_X1 U842 ( .A(n740), .B(KEYINPUT100), .Z(n743) );
  NAND2_X1 U843 ( .A1(n741), .A2(G2067), .ZN(n742) );
  NAND2_X1 U844 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U845 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U846 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n997), .A2(n748), .ZN(n749) );
  NAND2_X1 U848 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n754) );
  XNOR2_X1 U850 ( .A(n754), .B(n753), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n755), .A2(G171), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n773) );
  NOR2_X1 U853 ( .A1(n758), .A2(G2090), .ZN(n759) );
  XNOR2_X1 U854 ( .A(n759), .B(KEYINPUT102), .ZN(n761) );
  NOR2_X1 U855 ( .A1(n712), .A2(G1971), .ZN(n760) );
  NOR2_X1 U856 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U857 ( .A(KEYINPUT103), .B(n762), .Z(n763) );
  NAND2_X1 U858 ( .A1(n763), .A2(G303), .ZN(n765) );
  AND2_X1 U859 ( .A1(n773), .A2(n765), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n774), .A2(n764), .ZN(n768) );
  INV_X1 U861 ( .A(n765), .ZN(n766) );
  OR2_X1 U862 ( .A1(n766), .A2(G286), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U864 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U865 ( .A(KEYINPUT105), .B(KEYINPUT32), .ZN(n772) );
  AND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n779) );
  NAND2_X1 U867 ( .A1(G8), .A2(n775), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U869 ( .A1(G303), .A2(G1971), .ZN(n780) );
  XOR2_X1 U870 ( .A(n780), .B(KEYINPUT106), .Z(n782) );
  INV_X1 U871 ( .A(KEYINPUT33), .ZN(n781) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n995) );
  NOR2_X1 U873 ( .A1(n526), .A2(n995), .ZN(n783) );
  NAND2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U875 ( .A(n992), .ZN(n784) );
  NOR2_X1 U876 ( .A1(KEYINPUT33), .A2(n524), .ZN(n788) );
  NAND2_X1 U877 ( .A1(KEYINPUT33), .A2(n995), .ZN(n785) );
  NOR2_X1 U878 ( .A1(n712), .A2(n785), .ZN(n786) );
  XOR2_X1 U879 ( .A(KEYINPUT107), .B(n786), .Z(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n792), .B(n791), .ZN(n793) );
  XOR2_X1 U882 ( .A(G1981), .B(G305), .Z(n985) );
  NAND2_X1 U883 ( .A1(n793), .A2(n985), .ZN(n799) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G8), .A2(n794), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n797), .A2(n712), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n801), .B(n800), .ZN(n802) );
  NOR2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n837) );
  NOR2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n849) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n847) );
  NAND2_X1 U893 ( .A1(G104), .A2(n901), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G140), .A2(n624), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n809) );
  XOR2_X1 U896 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n808) );
  XNOR2_X1 U897 ( .A(n809), .B(n808), .ZN(n814) );
  NAND2_X1 U898 ( .A1(G116), .A2(n898), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G128), .A2(n899), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n815), .ZN(n917) );
  NOR2_X1 U904 ( .A1(n847), .A2(n917), .ZN(n943) );
  NAND2_X1 U905 ( .A1(n849), .A2(n943), .ZN(n816) );
  XNOR2_X1 U906 ( .A(KEYINPUT92), .B(n816), .ZN(n845) );
  NAND2_X1 U907 ( .A1(G119), .A2(n899), .ZN(n823) );
  NAND2_X1 U908 ( .A1(G107), .A2(n898), .ZN(n818) );
  NAND2_X1 U909 ( .A1(G95), .A2(n901), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n821) );
  NAND2_X1 U911 ( .A1(G131), .A2(n624), .ZN(n819) );
  XNOR2_X1 U912 ( .A(KEYINPUT93), .B(n819), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U915 ( .A(n824), .B(KEYINPUT94), .ZN(n916) );
  AND2_X1 U916 ( .A1(G1991), .A2(n916), .ZN(n833) );
  NAND2_X1 U917 ( .A1(G117), .A2(n898), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G129), .A2(n899), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n901), .A2(G105), .ZN(n827) );
  XOR2_X1 U921 ( .A(KEYINPUT38), .B(n827), .Z(n828) );
  NOR2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n624), .A2(G141), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n895) );
  AND2_X1 U925 ( .A1(G1996), .A2(n895), .ZN(n832) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n945) );
  INV_X1 U927 ( .A(n849), .ZN(n834) );
  NOR2_X1 U928 ( .A1(n945), .A2(n834), .ZN(n842) );
  INV_X1 U929 ( .A(n842), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n845), .A2(n835), .ZN(n836) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n839) );
  XNOR2_X1 U932 ( .A(G1986), .B(G290), .ZN(n1001) );
  NAND2_X1 U933 ( .A1(n1001), .A2(n849), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n852) );
  NOR2_X1 U935 ( .A1(G1996), .A2(n895), .ZN(n948) );
  NOR2_X1 U936 ( .A1(G1986), .A2(G290), .ZN(n840) );
  NOR2_X1 U937 ( .A1(G1991), .A2(n916), .ZN(n938) );
  NOR2_X1 U938 ( .A1(n840), .A2(n938), .ZN(n841) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U940 ( .A1(n948), .A2(n843), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n844), .B(KEYINPUT39), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n848) );
  NAND2_X1 U943 ( .A1(n847), .A2(n917), .ZN(n955) );
  NAND2_X1 U944 ( .A1(n848), .A2(n955), .ZN(n850) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n852), .A2(n851), .ZN(n854) );
  XNOR2_X1 U947 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(G329) );
  NAND2_X1 U949 ( .A1(n855), .A2(G2106), .ZN(n856) );
  XNOR2_X1 U950 ( .A(n856), .B(KEYINPUT112), .ZN(G217) );
  AND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G661), .A2(n857), .ZN(G259) );
  NAND2_X1 U953 ( .A1(G3), .A2(G1), .ZN(n858) );
  NAND2_X1 U954 ( .A1(n859), .A2(n858), .ZN(G188) );
  INV_X1 U956 ( .A(G108), .ZN(G238) );
  INV_X1 U957 ( .A(G96), .ZN(G221) );
  NOR2_X1 U958 ( .A1(n861), .A2(n860), .ZN(G325) );
  INV_X1 U959 ( .A(G325), .ZN(G261) );
  INV_X1 U960 ( .A(n862), .ZN(G319) );
  XOR2_X1 U961 ( .A(G2100), .B(G2096), .Z(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT42), .B(G2678), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U964 ( .A(KEYINPUT43), .B(G2090), .Z(n866) );
  XNOR2_X1 U965 ( .A(G2067), .B(G2072), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U968 ( .A(G2078), .B(G2084), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(G227) );
  XOR2_X1 U970 ( .A(G1971), .B(G1961), .Z(n872) );
  XNOR2_X1 U971 ( .A(G1981), .B(G1966), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U973 ( .A(n873), .B(KEYINPUT41), .Z(n875) );
  XNOR2_X1 U974 ( .A(G1996), .B(G1991), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U976 ( .A(G2474), .B(G1956), .Z(n877) );
  XNOR2_X1 U977 ( .A(G1986), .B(G1976), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(G229) );
  NAND2_X1 U980 ( .A1(G124), .A2(n899), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n880), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n898), .A2(G112), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G100), .A2(n901), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G136), .A2(n624), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U987 ( .A1(n886), .A2(n885), .ZN(G162) );
  NAND2_X1 U988 ( .A1(G115), .A2(n898), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G127), .A2(n899), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G139), .A2(n624), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G103), .A2(n901), .ZN(n892) );
  XNOR2_X1 U995 ( .A(KEYINPUT115), .B(n892), .ZN(n893) );
  NOR2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n932) );
  XOR2_X1 U997 ( .A(G162), .B(n932), .Z(n897) );
  XOR2_X1 U998 ( .A(G164), .B(n895), .Z(n896) );
  XNOR2_X1 U999 ( .A(n897), .B(n896), .ZN(n912) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n898), .ZN(n909) );
  NAND2_X1 U1001 ( .A1(n899), .A2(G130), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(KEYINPUT113), .B(n900), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(G106), .A2(n901), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(G142), .A2(n624), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1006 ( .A(KEYINPUT45), .B(n904), .Z(n905) );
  XNOR2_X1 U1007 ( .A(KEYINPUT114), .B(n905), .ZN(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n910), .B(KEYINPUT48), .ZN(n911) );
  XOR2_X1 U1011 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1012 ( .A(G160), .B(KEYINPUT46), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n937), .B(n915), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n920), .ZN(G395) );
  XNOR2_X1 U1018 ( .A(n921), .B(KEYINPUT116), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(G171), .B(G286), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n926), .ZN(G397) );
  NOR2_X1 U1023 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(G401), .A2(n928), .ZN(n929) );
  AND2_X1 U1026 ( .A1(G319), .A2(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1031 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1043) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n981) );
  XOR2_X1 U1033 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n958) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n935) );
  INV_X1 U1035 ( .A(G2072), .ZN(n933) );
  XNOR2_X1 U1036 ( .A(n933), .B(n932), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1038 ( .A(KEYINPUT50), .B(n936), .Z(n954) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1040 ( .A(KEYINPUT117), .B(n939), .Z(n941) );
  XNOR2_X1 U1041 ( .A(G160), .B(G2084), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n951) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(n949), .B(KEYINPUT51), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(n952), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n958), .B(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n981), .A2(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n960), .A2(G29), .ZN(n1041) );
  XOR2_X1 U1056 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n974) );
  XNOR2_X1 U1057 ( .A(G32), .B(n961), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(G2072), .B(G33), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(G27), .B(n966), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n969), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n970), .B(KEYINPUT121), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n974), .B(n973), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G35), .B(G2090), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n979) );
  XOR2_X1 U1071 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1072 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n981), .B(n980), .ZN(n983) );
  INV_X1 U1075 ( .A(G29), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(G11), .A2(n984), .ZN(n1039) );
  XNOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .ZN(n1011) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n987), .B(KEYINPUT57), .ZN(n1009) );
  XNOR2_X1 U1082 ( .A(G301), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n989), .B(n988), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n1004) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G166), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT123), .B(n996), .Z(n999) );
  XNOR2_X1 U1089 ( .A(n997), .B(G1956), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT124), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1341), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1037) );
  INV_X1 U1098 ( .A(G16), .ZN(n1035) );
  XOR2_X1 U1099 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n1033) );
  XNOR2_X1 U1100 ( .A(KEYINPUT59), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT125), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G1348), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G1341), .B(G19), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G1981), .B(G6), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G20), .B(G1956), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(n1020), .B(KEYINPUT60), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(G1976), .B(G23), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(G1986), .B(G24), .Z(n1023) );
  NAND2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(G1966), .B(G21), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(G1961), .B(G5), .ZN(n1028) );
  NOR2_X1 U1119 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1121 ( .A(n1033), .B(n1032), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1126 ( .A(n1043), .B(n1042), .ZN(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

