//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G1gat), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT16), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT92), .B(G8gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n217), .B2(KEYINPUT93), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n216), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n224));
  OR3_X1    g023(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT89), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(G29gat), .A3(G36gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n224), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT91), .ZN(new_n238));
  XOR2_X1   g037(.A(G43gat), .B(G50gat), .Z(new_n239));
  INV_X1    g038(.A(KEYINPUT15), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n236), .A2(new_n238), .A3(new_n224), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n225), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n226), .A2(KEYINPUT90), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n225), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n234), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n218), .A2(new_n221), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G229gat), .A2(G233gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n247), .A2(KEYINPUT17), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n247), .A2(KEYINPUT17), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n222), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n253), .A3(new_n251), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n255), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n208), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n260), .A2(new_n251), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT18), .A3(new_n253), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(new_n263), .A3(new_n255), .A4(new_n207), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT36), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT34), .ZN(new_n272));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n204), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n276));
  NOR2_X1   g075(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n281), .B(KEYINPUT65), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n288), .A2(new_n278), .A3(KEYINPUT25), .A4(new_n280), .ZN(new_n289));
  OAI22_X1  g088(.A1(new_n287), .A2(KEYINPUT25), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n281), .B1(new_n279), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT68), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n300), .B(new_n281), .C1(new_n279), .C2(new_n297), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n301), .C1(KEYINPUT26), .C2(new_n275), .ZN(new_n302));
  INV_X1    g101(.A(new_n295), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n293), .A2(KEYINPUT66), .A3(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n296), .A2(new_n302), .A3(new_n284), .A4(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G127gat), .B(G134gat), .Z(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT1), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G113gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT69), .B(G113gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(new_n309), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n308), .A2(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n306), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n290), .A2(new_n305), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n290), .B2(new_n305), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n272), .B(new_n273), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n290), .A2(new_n305), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n307), .A2(new_n311), .B1(new_n316), .B2(new_n306), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n319), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n272), .B1(new_n327), .B2(new_n273), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n273), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n330), .A3(new_n319), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(KEYINPUT70), .A3(new_n332), .ZN(new_n336));
  XOR2_X1   g135(.A(G15gat), .B(G43gat), .Z(new_n337));
  XNOR2_X1  g136(.A(G71gat), .B(G99gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n331), .B2(KEYINPUT32), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n331), .B(KEYINPUT32), .C1(new_n332), .C2(new_n340), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n329), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT71), .A4(new_n329), .ZN(new_n348));
  AOI211_X1 g147(.A(new_n271), .B(new_n344), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n343), .ZN(new_n351));
  INV_X1    g150(.A(new_n329), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n349), .B1(new_n271), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT2), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G148gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G155gat), .ZN(new_n366));
  INV_X1    g165(.A(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n359), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n371), .A3(new_n359), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n364), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(new_n362), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n359), .B1(new_n368), .B2(KEYINPUT2), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n365), .A2(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT4), .B1(new_n379), .B2(new_n325), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n325), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n325), .B1(new_n379), .B2(new_n387), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n365), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n377), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n394), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n383), .B1(new_n392), .B2(new_n318), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n325), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n397), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT79), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n394), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n318), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n397), .B1(new_n409), .B2(new_n381), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(new_n396), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n399), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G197gat), .B(G204gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT73), .B(G218gat), .ZN(new_n420));
  INV_X1    g219(.A(G211gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n422), .B2(KEYINPUT22), .ZN(new_n423));
  XNOR2_X1  g222(.A(G211gat), .B(G218gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n290), .B2(new_n305), .ZN(new_n427));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n290), .B2(new_n305), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n425), .C1(new_n429), .C2(new_n427), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G8gat), .B(G36gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT30), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT74), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT74), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n432), .B2(new_n434), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(KEYINPUT30), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n435), .A2(new_n439), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(KEYINPUT30), .B2(new_n444), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n418), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n397), .B1(new_n385), .B2(new_n394), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n409), .A2(new_n381), .A3(new_n397), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT39), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n454), .B(new_n416), .C1(new_n450), .C2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n397), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n395), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n458), .B2(new_n417), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT84), .B(new_n453), .C1(new_n456), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT40), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n417), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n454), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(KEYINPUT83), .A3(new_n417), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(KEYINPUT40), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n466), .A2(new_n453), .B1(KEYINPUT84), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n449), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT86), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n449), .B(new_n471), .C1(new_n462), .C2(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n387), .B1(new_n425), .B2(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n392), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n425), .B1(new_n476), .B2(KEYINPUT29), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G228gat), .ZN(new_n479));
  INV_X1    g278(.A(G233gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n475), .A2(G228gat), .A3(G233gat), .A4(new_n477), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G50gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G22gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(KEYINPUT82), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n491), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n482), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496));
  INV_X1    g295(.A(new_n411), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n404), .B2(new_n407), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n496), .B(new_n416), .C1(new_n498), .C2(new_n399), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n400), .A2(new_n403), .A3(KEYINPUT79), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n406), .B1(new_n405), .B2(new_n394), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n411), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n399), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n417), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n412), .A2(KEYINPUT81), .A3(new_n417), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT6), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n499), .B1(new_n508), .B2(new_n418), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n432), .A2(new_n434), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n439), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT38), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n444), .A2(KEYINPUT38), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n513), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n495), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n358), .B1(new_n473), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n444), .A2(KEYINPUT30), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n439), .B2(new_n435), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n442), .B2(new_n445), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n499), .C1(new_n508), .C2(new_n418), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n495), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n495), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n350), .A2(new_n527), .A3(new_n353), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n499), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT81), .B1(new_n412), .B2(new_n417), .ZN(new_n532));
  NOR4_X1   g331(.A1(new_n498), .A2(new_n505), .A3(new_n399), .A4(new_n416), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n496), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n418), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n350), .A2(new_n527), .A3(KEYINPUT88), .A4(new_n353), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n530), .A2(new_n536), .A3(new_n523), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n492), .A2(new_n540), .A3(new_n494), .ZN(new_n541));
  AND4_X1   g340(.A1(new_n350), .A2(new_n355), .A3(new_n356), .A4(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(KEYINPUT87), .A3(new_n536), .A4(new_n523), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n350), .A2(new_n355), .A3(new_n541), .A4(new_n356), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n524), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n270), .B1(new_n526), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G183gat), .B(G211gat), .Z(new_n550));
  AND2_X1   g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(G57gat), .A2(G64gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n555), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT94), .Z(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n572));
  OR3_X1    g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n556), .A2(new_n562), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n250), .B1(KEYINPUT21), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n573), .B2(new_n574), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n550), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n574), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n576), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n583));
  INV_X1    g382(.A(new_n550), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(KEYINPUT8), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n597), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n600), .A2(new_n590), .A3(new_n601), .A4(new_n591), .ZN(new_n602));
  INV_X1    g401(.A(new_n594), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT96), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n257), .B2(new_n258), .ZN(new_n608));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n248), .B2(new_n606), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n587), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT97), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n615), .B(new_n587), .C1(new_n608), .C2(new_n612), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n608), .A2(new_n612), .A3(new_n587), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n614), .A2(new_n616), .A3(new_n617), .A4(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n625), .A3(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n586), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT99), .B(KEYINPUT10), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n602), .A2(new_n635), .A3(new_n603), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n603), .B1(new_n602), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n575), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n563), .B(new_n599), .C1(new_n604), .C2(new_n605), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n575), .A2(KEYINPUT10), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n606), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n632), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n632), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n648), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n549), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n536), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n211), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n654), .A2(new_n523), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT42), .B1(new_n657), .B2(KEYINPUT100), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  INV_X1    g462(.A(new_n657), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(G8gat), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n657), .A2(KEYINPUT101), .A3(new_n214), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n661), .B(new_n662), .C1(new_n665), .C2(new_n666), .ZN(G1325gat));
  INV_X1    g466(.A(new_n358), .ZN(new_n668));
  OAI21_X1  g467(.A(G15gat), .B1(new_n654), .B2(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n357), .A2(G15gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n654), .B2(new_n670), .ZN(G1326gat));
  NAND3_X1  g470(.A1(new_n549), .A2(new_n495), .A3(new_n653), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT102), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n580), .A2(new_n585), .ZN(new_n676));
  INV_X1    g475(.A(new_n652), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n630), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n536), .A2(G29gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n549), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n525), .A2(KEYINPUT103), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n524), .A2(new_n685), .A3(new_n495), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n520), .A2(new_n687), .B1(new_n539), .B2(new_n547), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n683), .B1(new_n688), .B2(new_n630), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n629), .A2(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n473), .A2(new_n519), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n692), .A2(new_n525), .A3(new_n668), .ZN(new_n693));
  AOI22_X1  g492(.A1(KEYINPUT35), .A2(new_n538), .B1(new_n543), .B2(new_n546), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n270), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n689), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n536), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1328gat));
  NAND2_X1  g500(.A1(new_n549), .A2(new_n679), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(G36gat), .A3(new_n523), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n697), .B2(new_n523), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n357), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n549), .A2(new_n708), .A3(new_n709), .A4(new_n679), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT105), .Z(new_n711));
  NAND4_X1  g510(.A1(new_n689), .A2(new_n358), .A3(new_n695), .A4(new_n696), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(G43gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n708), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n690), .B1(new_n526), .B2(new_n548), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n520), .A2(new_n687), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n548), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n629), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(new_n721), .B2(new_n683), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n722), .A2(KEYINPUT106), .A3(new_n358), .A4(new_n696), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n715), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI211_X1 g526(.A(KEYINPUT107), .B(new_n725), .C1(new_n717), .C2(new_n723), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n714), .B1(new_n727), .B2(new_n728), .ZN(G1330gat));
  NOR2_X1   g528(.A1(new_n702), .A2(new_n527), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n495), .A2(G50gat), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n730), .A2(G50gat), .B1(new_n697), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1331gat));
  NOR3_X1   g533(.A1(new_n631), .A2(new_n269), .A3(new_n677), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n536), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(G57gat), .Z(G1332gat));
  AOI211_X1 g537(.A(new_n523), .B(new_n736), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  NAND4_X1  g540(.A1(new_n720), .A2(G71gat), .A3(new_n358), .A4(new_n735), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n736), .A2(new_n357), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n743), .B(new_n744), .C1(G71gat), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n736), .A2(new_n527), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g548(.A1(new_n586), .A2(new_n269), .A3(new_n677), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n722), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n536), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n586), .A2(new_n269), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n720), .A2(new_n629), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(KEYINPUT110), .A3(new_n755), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n509), .A2(new_n596), .A3(new_n652), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n752), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  OAI21_X1  g562(.A(G92gat), .B1(new_n751), .B2(new_n523), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n523), .A2(G92gat), .A3(new_n677), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n763), .B(new_n764), .C1(new_n760), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n754), .A2(KEYINPUT111), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n755), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n767), .A2(new_n773), .ZN(G1337gat));
  NAND3_X1  g573(.A1(new_n722), .A2(new_n358), .A3(new_n750), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G99gat), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n357), .A2(G99gat), .A3(new_n677), .ZN(new_n777));
  OAI211_X1 g576(.A(KEYINPUT112), .B(new_n776), .C1(new_n760), .C2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779));
  INV_X1    g578(.A(new_n776), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n758), .B2(new_n759), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n751), .B2(new_n527), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n785));
  NOR3_X1   g584(.A1(new_n527), .A2(G106gat), .A3(new_n677), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n784), .B(new_n785), .C1(new_n760), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n770), .A3(new_n786), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n266), .B2(new_n253), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n260), .A2(new_n251), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n795), .A2(KEYINPUT117), .A3(G229gat), .A4(G233gat), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n252), .A2(new_n254), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n206), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(new_n268), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n801), .B(new_n632), .C1(new_n640), .C2(new_n642), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n648), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n644), .A2(new_n633), .ZN(new_n804));
  INV_X1    g603(.A(new_n642), .ZN(new_n805));
  INV_X1    g604(.A(new_n632), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n643), .A3(KEYINPUT114), .A4(KEYINPUT54), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n643), .A2(KEYINPUT54), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n640), .A2(new_n642), .A3(new_n632), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT116), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n813), .A2(KEYINPUT55), .A3(new_n808), .A4(new_n803), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT115), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n809), .A2(new_n818), .A3(KEYINPUT55), .A4(new_n813), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n649), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n629), .A2(new_n800), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n815), .A2(new_n269), .A3(new_n820), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n268), .A3(new_n652), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n629), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n676), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n586), .A2(new_n270), .A3(new_n630), .A4(new_n677), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n495), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n523), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n536), .A2(new_n357), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n270), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n826), .A2(new_n827), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n530), .A2(new_n537), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n536), .A2(new_n832), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n310), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n269), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n835), .A2(new_n841), .ZN(G1340gat));
  AOI21_X1  g641(.A(G120gat), .B1(new_n839), .B2(new_n652), .ZN(new_n843));
  INV_X1    g642(.A(new_n834), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n677), .A2(new_n308), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n834), .B2(new_n676), .ZN(new_n847));
  INV_X1    g646(.A(G127gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n839), .A2(new_n848), .A3(new_n586), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1342gat));
  OAI21_X1  g649(.A(G134gat), .B1(new_n834), .B2(new_n630), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n536), .B1(new_n826), .B2(new_n827), .ZN(new_n852));
  INV_X1    g651(.A(G134gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n630), .A2(new_n832), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n837), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT56), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n358), .A2(new_n527), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n836), .A2(new_n838), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n363), .A3(new_n269), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n668), .A2(new_n838), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n676), .A2(new_n269), .A3(new_n629), .A4(new_n652), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n817), .A2(new_n819), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n813), .A2(new_n808), .A3(new_n803), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n649), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n269), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n866), .B1(new_n865), .B2(new_n869), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT120), .B(new_n824), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n630), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n865), .A2(new_n869), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n269), .A3(new_n870), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT120), .B1(new_n877), .B2(new_n824), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n821), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n864), .B1(new_n879), .B2(new_n676), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n880), .A2(new_n881), .A3(new_n527), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n836), .B2(new_n495), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n269), .B(new_n863), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n861), .B1(new_n884), .B2(G141gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n824), .B1(new_n871), .B2(new_n872), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n630), .A3(new_n873), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n586), .B1(new_n892), .B2(new_n821), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT57), .B(new_n495), .C1(new_n893), .C2(new_n864), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n836), .A2(new_n495), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n881), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n270), .B(new_n862), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n860), .B1(new_n897), .B2(new_n363), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n888), .B1(new_n898), .B2(KEYINPUT58), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n886), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n887), .B1(new_n899), .B2(new_n900), .ZN(G1344gat));
  AND2_X1   g700(.A1(new_n852), .A2(new_n858), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n902), .A2(new_n361), .A3(new_n523), .A4(new_n652), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n881), .B(new_n495), .C1(new_n893), .C2(new_n864), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(KEYINPUT57), .ZN(new_n906));
  AND4_X1   g705(.A1(new_n652), .A2(new_n905), .A3(new_n906), .A4(new_n863), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n361), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n862), .B1(new_n894), .B2(new_n896), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n652), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(KEYINPUT122), .A3(new_n904), .A4(G148gat), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n677), .B(new_n862), .C1(new_n894), .C2(new_n896), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n904), .A2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n903), .B1(new_n911), .B2(new_n919), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n859), .A2(new_n366), .A3(new_n586), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n912), .A2(new_n586), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n366), .ZN(G1346gat));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n367), .A3(new_n854), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT124), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n912), .A2(new_n629), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n367), .B2(new_n926), .ZN(G1347gat));
  AOI21_X1  g726(.A(new_n509), .B1(new_n826), .B2(new_n827), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n837), .A2(new_n832), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n269), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n536), .A2(new_n832), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n357), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT125), .Z(new_n934));
  AND2_X1   g733(.A1(new_n831), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n270), .A2(new_n204), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  AOI21_X1  g736(.A(new_n274), .B1(new_n935), .B2(new_n652), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n930), .A2(new_n274), .A3(new_n652), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n938), .A2(new_n939), .ZN(G1349gat));
  OAI211_X1 g739(.A(new_n586), .B(new_n934), .C1(new_n829), .C2(new_n830), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G183gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n930), .A2(new_n291), .A3(new_n586), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n292), .A3(new_n629), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n831), .A2(new_n629), .A3(new_n934), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n947), .A2(new_n948), .A3(G190gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n947), .B2(G190gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  INV_X1    g750(.A(G197gat), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n905), .A2(new_n906), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n358), .A2(new_n932), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n269), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(KEYINPUT126), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(KEYINPUT126), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n858), .A2(new_n832), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n928), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n952), .A3(new_n269), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(G1352gat));
  INV_X1    g761(.A(new_n960), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n963), .A2(G204gat), .A3(new_n677), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n953), .A2(new_n652), .A3(new_n954), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G204gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n960), .A2(new_n421), .A3(new_n586), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n586), .A2(new_n905), .A3(new_n906), .A4(new_n954), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n421), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n905), .A2(new_n906), .A3(new_n586), .A4(new_n954), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n972), .A2(KEYINPUT63), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n960), .B2(new_n629), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n953), .A2(new_n954), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n630), .A2(new_n420), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1355gat));
endmodule


