//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n454), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT3), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n476), .A2(G137), .A3(new_n464), .A4(new_n466), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n467), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n479), .A2(G101), .A3(new_n464), .A4(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n474), .A2(new_n475), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G101), .A4(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(KEYINPUT70), .A3(new_n477), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n473), .B1(new_n486), .B2(new_n492), .ZN(G160));
  NAND2_X1  g068(.A1(new_n476), .A2(new_n466), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n464), .A2(G112), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n494), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n466), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT68), .B(G2104), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT3), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(new_n464), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n506), .B2(G136), .ZN(G162));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n503), .A2(new_n508), .A3(G126), .A4(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n476), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n476), .A2(G138), .A3(new_n464), .A4(new_n466), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n515));
  INV_X1    g090(.A(G138), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(G2105), .ZN(new_n517));
  AND4_X1   g092(.A1(new_n515), .A2(new_n517), .A3(new_n466), .A4(new_n468), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n521));
  INV_X1    g096(.A(G114), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G2105), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G164));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n531), .B1(new_n528), .B2(G543), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n532), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT6), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G88), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G50), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n535), .A2(new_n544), .ZN(G166));
  AND2_X1   g120(.A1(new_n532), .A2(new_n539), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n546), .A2(G89), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  INV_X1    g125(.A(G51), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n548), .B(new_n550), .C1(new_n551), .C2(new_n542), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n547), .A2(new_n552), .ZN(G168));
  AOI22_X1  g128(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n534), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(G90), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n540), .A2(new_n556), .B1(new_n542), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(G171));
  AOI22_X1  g134(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(new_n542), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n546), .A2(G81), .B1(new_n563), .B2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G188));
  AND3_X1   g147(.A1(new_n539), .A2(G53), .A3(G543), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT9), .Z(new_n574));
  NAND2_X1  g149(.A1(new_n546), .A2(G91), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n532), .A2(G65), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT76), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n546), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n563), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND4_X1  g162(.A1(new_n536), .A2(new_n538), .A3(G48), .A4(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT77), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n532), .A2(G86), .A3(new_n539), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n532), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n534), .C2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n534), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n540), .A2(new_n595), .B1(new_n542), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n594), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n546), .A2(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT78), .B(G66), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n532), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n530), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n563), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT79), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G168), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT80), .ZN(new_n614));
  XNOR2_X1  g189(.A(G299), .B(KEYINPUT81), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n609), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n609), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n488), .A2(new_n464), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(new_n469), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT83), .B(G2100), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT84), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n506), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n495), .A2(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n464), .A2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NOR2_X1   g213(.A1(new_n629), .A2(new_n630), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n632), .A2(new_n638), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT15), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2435), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2435), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n660), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n662), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n664), .B(new_n665), .C1(new_n661), .C2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(KEYINPUT18), .B1(new_n665), .B2(new_n658), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n665), .A2(KEYINPUT18), .A3(new_n658), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n676), .B2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(new_n506), .A2(G131), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n695));
  OR2_X1    g270(.A1(G95), .A2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT89), .Z(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G119), .B2(new_n495), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT90), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT35), .B(G1991), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n711), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n708), .A2(new_n715), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n722), .A2(KEYINPUT93), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G24), .ZN(new_n725));
  INV_X1    g300(.A(G290), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(new_n691), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n705), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT36), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  INV_X1    g306(.A(G34), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(KEYINPUT24), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G160), .B2(new_n731), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT98), .Z(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G2084), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G2090), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(G2090), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n716), .A2(KEYINPUT23), .A3(G20), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n746));
  INV_X1    g321(.A(G20), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G299), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n745), .B(new_n748), .C1(new_n749), .C2(new_n716), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1956), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n738), .A2(new_n743), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n731), .A2(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n731), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT101), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(G168), .A2(new_n716), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n716), .B2(G21), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n755), .A2(G2078), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n756), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n495), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  INV_X1    g339(.A(G105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(new_n625), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G141), .B2(new_n506), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT27), .B(G1996), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT99), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n637), .A2(new_n731), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT100), .Z(new_n773));
  NAND4_X1  g348(.A1(new_n752), .A2(new_n760), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n609), .A2(G16), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G4), .B2(G16), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n776), .A2(G4), .A3(G16), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT28), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n731), .A2(G26), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n495), .A2(G128), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n506), .A2(G140), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n464), .A2(G116), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n782), .B(new_n783), .C1(new_n789), .C2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n782), .B2(new_n783), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT96), .B(G2067), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n716), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n716), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n716), .A2(G19), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n565), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1341), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT30), .B(G28), .Z(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G29), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n768), .B2(new_n770), .ZN(new_n806));
  AND4_X1   g381(.A1(new_n797), .A2(new_n801), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n731), .A2(G33), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT25), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n506), .A2(G139), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT97), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n810), .B(new_n811), .C1(G2105), .C2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n731), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(G2072), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n737), .A2(G2084), .B1(G2078), .B2(new_n755), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n793), .A2(new_n807), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n774), .A2(new_n781), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(KEYINPUT103), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT103), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n774), .A2(new_n818), .A3(new_n821), .A4(new_n781), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n730), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(G311));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n730), .B(KEYINPUT104), .C1(new_n820), .C2(new_n822), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  AOI22_X1  g403(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n534), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n540), .A2(new_n831), .B1(new_n542), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT105), .B(G860), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n609), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n565), .B(new_n834), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT39), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n843), .B2(new_n836), .ZN(G145));
  XNOR2_X1  g419(.A(G160), .B(KEYINPUT106), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(G162), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n637), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n495), .A2(G130), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n464), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G142), .B2(new_n506), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n767), .B(new_n852), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n814), .B(new_n789), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n523), .B1(new_n509), .B2(new_n511), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT107), .ZN(new_n857));
  AOI211_X1 g432(.A(new_n857), .B(new_n518), .C1(new_n513), .C2(KEYINPUT4), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT107), .B1(new_n514), .B2(new_n519), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n627), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n855), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n701), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n854), .A2(new_n863), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g443(.A1(new_n835), .A2(new_n612), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n620), .B(new_n841), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n608), .B(G299), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(KEYINPUT41), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n602), .A2(new_n607), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n749), .A2(new_n608), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT108), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(KEYINPUT108), .A3(G299), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n874), .B1(KEYINPUT41), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n870), .B(new_n873), .C1(new_n871), .C2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(new_n870), .ZN(new_n885));
  XNOR2_X1  g460(.A(G166), .B(G288), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G290), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n885), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n869), .B1(new_n890), .B2(new_n612), .ZN(G295));
  OAI21_X1  g466(.A(new_n869), .B1(new_n890), .B2(new_n612), .ZN(G331));
  XNOR2_X1  g467(.A(G301), .B(G168), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n841), .B(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n873), .B(new_n894), .C1(new_n882), .C2(new_n871), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n884), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  INV_X1    g474(.A(new_n888), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g476(.A(KEYINPUT110), .B(new_n888), .C1(new_n895), .C2(new_n896), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n865), .B(new_n897), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n841), .A2(new_n893), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n841), .A2(new_n893), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT41), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n884), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n872), .A2(KEYINPUT111), .A3(KEYINPUT41), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n894), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n900), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n917), .B(new_n918), .C1(new_n901), .C2(new_n902), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n904), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n905), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n903), .A2(new_n904), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n904), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT45), .B1(new_n860), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n473), .ZN(new_n929));
  INV_X1    g504(.A(new_n492), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT70), .B1(new_n491), .B2(new_n477), .ZN(new_n931));
  OAI211_X1 g506(.A(G40), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G2067), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n789), .B(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n767), .B(G1996), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n701), .A2(new_n704), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n701), .A2(new_n704), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT113), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n691), .B2(new_n726), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n935), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n520), .A2(new_n857), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n514), .A2(KEYINPUT107), .A3(new_n519), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n952), .B2(new_n856), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n949), .B(new_n933), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n486), .A2(new_n492), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n956), .A2(new_n954), .A3(G40), .A4(new_n929), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n860), .A2(new_n927), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT116), .B(new_n957), .C1(new_n958), .C2(new_n932), .ZN(new_n959));
  INV_X1    g534(.A(G2090), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n856), .B2(new_n520), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n954), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n955), .A2(new_n959), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n525), .A2(new_n927), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n967), .A3(new_n933), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n719), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G8), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  NOR2_X1   g547(.A1(G166), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT55), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n974), .A2(KEYINPUT115), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(KEYINPUT115), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n975), .B(new_n976), .C1(KEYINPUT55), .C2(new_n973), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n710), .A2(G1976), .ZN(new_n980));
  OAI211_X1 g555(.A(G8), .B(new_n980), .C1(new_n958), .C2(new_n932), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT52), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n953), .A2(new_n933), .ZN(new_n983));
  NOR2_X1   g558(.A1(G305), .A2(G1981), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G305), .A2(G1981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(KEYINPUT49), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  AND2_X1   g563(.A1(G305), .A2(G1981), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n984), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n983), .A2(new_n987), .A3(G8), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n983), .A2(G8), .A3(new_n980), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n982), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n982), .A2(new_n991), .A3(new_n994), .A4(KEYINPUT117), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n969), .A2(KEYINPUT114), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n954), .B1(new_n525), .B2(new_n927), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(new_n932), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n860), .A2(new_n954), .A3(new_n927), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n960), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n968), .A2(new_n1005), .A3(new_n719), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(G8), .A3(new_n977), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n979), .A2(new_n999), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2084), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(new_n1010), .A3(new_n1003), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n966), .B(G1384), .C1(new_n856), .C2(new_n520), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n928), .A2(new_n1012), .A3(new_n932), .ZN(new_n1013));
  OAI211_X1 g588(.A(G168), .B(new_n1011), .C1(new_n1013), .C2(G1966), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(KEYINPUT122), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n933), .B1(new_n953), .B2(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n756), .B1(new_n1020), .B2(new_n1012), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1011), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(G8), .A3(G286), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT122), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1015), .A2(new_n1024), .A3(new_n1016), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT123), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1019), .A2(new_n1023), .A3(new_n1028), .A4(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n955), .A2(new_n962), .A3(new_n959), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT119), .B(G1956), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  AND4_X1   g609(.A1(new_n933), .A2(new_n964), .A3(new_n967), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G299), .B(KEYINPUT57), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1038), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(new_n1040), .A3(new_n1036), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT120), .B(G1996), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n964), .A2(new_n967), .A3(new_n933), .A4(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(new_n800), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n958), .B2(new_n932), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1049), .B2(new_n566), .ZN(new_n1050));
  AOI211_X1 g625(.A(KEYINPUT59), .B(new_n565), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1348), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n958), .A2(G2067), .A3(new_n932), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n875), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n860), .A2(new_n954), .A3(new_n927), .ZN(new_n1057));
  OAI211_X1 g632(.A(G160), .B(G40), .C1(new_n961), .C2(new_n954), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n780), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n953), .A2(new_n936), .A3(new_n933), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n608), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT60), .A4(new_n608), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1052), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1040), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1035), .B(new_n1038), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1042), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1056), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1041), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n968), .B2(G2078), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n796), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n928), .A2(new_n932), .ZN(new_n1076));
  INV_X1    g651(.A(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1074), .B(new_n1075), .C1(new_n1078), .C2(new_n1012), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1079), .B2(G301), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1077), .A4(new_n964), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(G301), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(G171), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1079), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1082), .A2(G171), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1072), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1069), .A2(new_n1071), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT62), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1030), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1027), .A2(KEYINPUT62), .A3(new_n1029), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1009), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n972), .B(G286), .C1(new_n1021), .C2(new_n1011), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n979), .A2(new_n999), .A3(new_n1008), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1007), .A2(G8), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n995), .B1(new_n1100), .B2(new_n978), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(KEYINPUT63), .A3(new_n1008), .A4(new_n1096), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1008), .A2(new_n995), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n991), .A2(new_n992), .A3(new_n710), .ZN(new_n1105));
  OAI211_X1 g680(.A(G8), .B(new_n983), .C1(new_n1105), .C2(new_n984), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1103), .A2(new_n1109), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n948), .B1(new_n1095), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n934), .B1(new_n937), .B2(new_n767), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n934), .A2(G1996), .ZN(new_n1115));
  NOR2_X1   g690(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT47), .ZN(new_n1119));
  INV_X1    g694(.A(new_n940), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n939), .A2(new_n1120), .B1(G2067), .B2(new_n789), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n935), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n945), .A2(new_n935), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT48), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n942), .B2(new_n934), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1119), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1112), .A2(new_n1127), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g703(.A1(new_n656), .A2(new_n462), .A3(new_n672), .ZN(new_n1130));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1131));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g706(.A1(new_n656), .A2(KEYINPUT126), .A3(new_n462), .A4(new_n672), .ZN(new_n1133));
  AOI21_X1  g707(.A(G229), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g708(.A1(new_n922), .A2(new_n867), .A3(new_n923), .A4(new_n1134), .ZN(G225));
  INV_X1    g709(.A(G225), .ZN(G308));
endmodule


