//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n217), .B1(new_n212), .B2(new_n211), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(KEYINPUT24), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT82), .ZN(new_n245));
  AND2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  OAI211_X1 g0047(.A(new_n207), .B(G87), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT81), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT81), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n250), .A2(new_n251), .A3(new_n207), .A4(G87), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT22), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(new_n252), .A3(KEYINPUT22), .ZN(new_n256));
  OR3_X1    g0056(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AND4_X1   g0061(.A1(new_n245), .A2(new_n255), .A3(new_n256), .A4(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n253), .B2(new_n254), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n245), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n244), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n255), .A2(new_n256), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT82), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n245), .A3(new_n256), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(KEYINPUT24), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n213), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n206), .A2(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G107), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G20), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT25), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n206), .A2(G33), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(new_n213), .A4(new_n270), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(G107), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n272), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT5), .A2(G41), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT5), .A2(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n206), .B(G45), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT66), .ZN(new_n287));
  AND2_X1   g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n213), .ZN(new_n289));
  AND2_X1   g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(KEYINPUT66), .A3(new_n291), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n286), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G294), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n294), .A2(KEYINPUT83), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(KEYINPUT83), .ZN(new_n296));
  OAI21_X1  g0096(.A(G33), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  OAI211_X1 g0098(.A(G250), .B(new_n298), .C1(new_n246), .C2(new_n247), .ZN(new_n299));
  OAI211_X1 g0099(.A(G257), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n288), .A2(new_n213), .ZN(new_n302));
  AOI22_X1  g0102(.A1(G264), .A2(new_n293), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n288), .A2(new_n287), .A3(new_n213), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT66), .B1(new_n290), .B2(new_n291), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n286), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(KEYINPUT77), .A3(G274), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT77), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n289), .A2(G274), .A3(new_n292), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n286), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G169), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n313), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n283), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n278), .A2(G116), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n281), .B2(G116), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G283), .ZN(new_n320));
  INV_X1    g0120(.A(G97), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n207), .C1(G33), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G116), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G20), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n271), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT80), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n326), .B2(new_n325), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(KEYINPUT80), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n319), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT21), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  OAI211_X1 g0133(.A(G264), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n334));
  OAI211_X1 g0134(.A(G257), .B(new_n298), .C1(new_n246), .C2(new_n247), .ZN(new_n335));
  INV_X1    g0135(.A(G303), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n250), .ZN(new_n337));
  AOI22_X1  g0137(.A1(G270), .A2(new_n293), .B1(new_n337), .B2(new_n302), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n332), .B(new_n333), .C1(new_n338), .C2(new_n312), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n312), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n315), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n331), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n338), .B2(new_n312), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n332), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n338), .A2(new_n312), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n331), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n303), .A2(new_n312), .A3(KEYINPUT84), .A4(new_n349), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT84), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n313), .B2(new_n347), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n313), .A2(G190), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n272), .A2(new_n282), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n278), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n321), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n280), .B2(new_n321), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT76), .ZN(new_n362));
  XNOR2_X1  g0162(.A(G97), .B(G107), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n364), .A2(new_n321), .A3(G107), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G20), .A2(G33), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(G20), .B1(G77), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT3), .ZN(new_n371));
  INV_X1    g0171(.A(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n207), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n379));
  NOR4_X1   g0179(.A1(new_n246), .A2(new_n247), .A3(new_n377), .A4(G20), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n370), .B1(new_n381), .B2(new_n275), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n362), .B1(new_n382), .B2(new_n271), .ZN(new_n383));
  AND4_X1   g0183(.A1(G257), .A2(new_n286), .A3(new_n289), .A4(new_n292), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n308), .B2(new_n311), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n298), .A2(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n250), .A2(G244), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G244), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n373), .B2(new_n374), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n387), .B(new_n320), .C1(new_n389), .C2(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n250), .A2(G250), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n298), .B1(new_n391), .B2(KEYINPUT4), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n302), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n385), .A2(new_n349), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(G200), .B1(new_n385), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n383), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n361), .B(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n366), .B1(new_n364), .B2(new_n363), .ZN(new_n399));
  INV_X1    g0199(.A(G77), .ZN(new_n400));
  INV_X1    g0200(.A(new_n369), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n399), .A2(new_n207), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n375), .A2(new_n377), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT72), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n405));
  INV_X1    g0205(.A(new_n380), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n407), .B2(G107), .ZN(new_n408));
  INV_X1    g0208(.A(new_n271), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n398), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n385), .A2(G179), .A3(new_n393), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n333), .B1(new_n385), .B2(new_n393), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(G238), .B(new_n298), .C1(new_n246), .C2(new_n247), .ZN(new_n414));
  OAI211_X1 g0214(.A(G244), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n372), .C2(new_n323), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n302), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n206), .A2(G45), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G250), .ZN(new_n419));
  INV_X1    g0219(.A(G274), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n306), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n417), .A2(G190), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n347), .B1(new_n417), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n250), .A2(new_n207), .A3(G68), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(G20), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(KEYINPUT19), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G87), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n321), .A3(new_n275), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(new_n430), .A3(new_n321), .A4(new_n275), .ZN(new_n434));
  NAND3_X1  g0234(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n432), .A2(new_n434), .B1(new_n207), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n271), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT15), .B(G87), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n359), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT79), .B1(new_n280), .B2(new_n430), .ZN(new_n440));
  OR3_X1    g0240(.A1(new_n280), .A2(KEYINPUT79), .A3(new_n430), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n437), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n417), .A2(G179), .A3(new_n422), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n416), .A2(new_n302), .B1(new_n306), .B2(new_n421), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n333), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n437), .B(new_n439), .C1(new_n438), .C2(new_n280), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n425), .A2(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n396), .A2(new_n413), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n317), .A2(new_n352), .A3(new_n358), .A4(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n369), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT8), .B(G58), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n207), .A2(G33), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n271), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n278), .A2(new_n202), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n271), .B1(new_n206), .B2(G20), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n202), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n289), .A2(new_n460), .A3(new_n292), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT67), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT67), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n289), .A2(new_n292), .A3(new_n463), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G226), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(G1698), .B1(new_n373), .B2(new_n374), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n246), .A2(new_n247), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n468), .A2(G222), .B1(new_n469), .B2(G77), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n298), .B1(new_n373), .B2(new_n374), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G223), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n302), .ZN(new_n474));
  INV_X1    g0274(.A(new_n310), .ZN(new_n475));
  INV_X1    g0275(.A(new_n460), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G179), .ZN(new_n480));
  OAI21_X1  g0280(.A(G169), .B1(new_n478), .B2(new_n467), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n459), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(G190), .ZN(new_n483));
  OAI21_X1  g0283(.A(G200), .B1(new_n467), .B2(new_n478), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n458), .B(KEYINPUT9), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT10), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n484), .B2(KEYINPUT68), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n488), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n482), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G20), .A2(G77), .ZN(new_n492));
  OAI221_X1 g0292(.A(new_n492), .B1(new_n451), .B2(new_n401), .C1(new_n452), .C2(new_n438), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n493), .A2(new_n271), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n359), .A2(new_n400), .ZN(new_n495));
  INV_X1    g0295(.A(new_n456), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n400), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n465), .A2(G244), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n471), .A2(G238), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n250), .A2(G232), .A3(new_n298), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n469), .A2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(new_n302), .B1(new_n475), .B2(new_n476), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n347), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n500), .A2(new_n505), .A3(new_n349), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(G169), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n500), .A2(new_n505), .A3(G179), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n498), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n465), .A2(G238), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT13), .ZN(new_n514));
  OAI211_X1 g0314(.A(G232), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n515));
  OAI211_X1 g0315(.A(G226), .B(new_n298), .C1(new_n246), .C2(new_n247), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n427), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n302), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n513), .A2(new_n514), .A3(new_n477), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n477), .A2(new_n518), .ZN(new_n520));
  INV_X1    g0320(.A(G238), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n462), .B2(new_n464), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT13), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n347), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G190), .B2(new_n524), .ZN(new_n526));
  INV_X1    g0326(.A(G68), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n369), .A2(G50), .B1(G20), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n400), .B2(new_n452), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT11), .B1(new_n529), .B2(new_n271), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(G68), .B2(new_n456), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(KEYINPUT11), .A3(new_n271), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n274), .A2(G20), .A3(new_n527), .ZN(new_n533));
  OR3_X1    g0333(.A1(new_n533), .A2(KEYINPUT69), .A3(KEYINPUT12), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT69), .B1(new_n533), .B2(KEYINPUT12), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(KEYINPUT12), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n509), .B(new_n512), .C1(new_n526), .C2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n491), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT75), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n306), .A2(G232), .A3(new_n460), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n477), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT74), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n372), .A2(new_n430), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n468), .B2(G223), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT73), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n471), .B2(G226), .ZN(new_n549));
  OAI211_X1 g0349(.A(G226), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n545), .B(new_n547), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n302), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n471), .A2(new_n548), .A3(G226), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n545), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n349), .B(new_n544), .C1(new_n553), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n477), .A2(new_n543), .ZN(new_n559));
  INV_X1    g0359(.A(new_n302), .ZN(new_n560));
  OAI211_X1 g0360(.A(G223), .B(new_n298), .C1(new_n246), .C2(new_n247), .ZN(new_n561));
  INV_X1    g0361(.A(new_n546), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n554), .B2(new_n555), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n545), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n547), .B1(new_n549), .B2(new_n551), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n559), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n558), .B1(new_n568), .B2(G200), .ZN(new_n569));
  INV_X1    g0369(.A(new_n451), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n359), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n496), .B2(new_n570), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT71), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT70), .ZN(new_n574));
  AND2_X1   g0374(.A1(G58), .A2(G68), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(G20), .C1(new_n575), .C2(new_n201), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n369), .A2(G159), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g0378(.A(G58), .B(G68), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n579), .B2(G20), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n573), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT7), .B1(new_n469), .B2(new_n207), .ZN(new_n582));
  OAI21_X1  g0382(.A(G68), .B1(new_n582), .B2(new_n380), .ZN(new_n583));
  OAI21_X1  g0383(.A(G20), .B1(new_n575), .B2(new_n201), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT70), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(KEYINPUT71), .A3(new_n576), .A4(new_n577), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT16), .A4(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n271), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT16), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n379), .A2(new_n380), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n527), .B1(new_n590), .B2(new_n405), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n581), .A2(new_n586), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n572), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n569), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT17), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n315), .B(new_n544), .C1(new_n553), .C2(new_n557), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n568), .B2(G169), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT18), .B1(new_n599), .B2(new_n594), .ZN(new_n600));
  INV_X1    g0400(.A(new_n572), .ZN(new_n601));
  INV_X1    g0401(.A(new_n592), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n407), .A2(G68), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT16), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n587), .A2(new_n271), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT18), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n544), .B1(new_n553), .B2(new_n557), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n333), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n606), .A2(new_n607), .A3(new_n598), .A4(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n569), .A2(new_n594), .A3(KEYINPUT17), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n597), .A2(new_n600), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n519), .A2(new_n523), .A3(G179), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n333), .B1(new_n519), .B2(new_n523), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT14), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI211_X1 g0417(.A(KEYINPUT14), .B(new_n333), .C1(new_n519), .C2(new_n523), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n538), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n541), .A2(new_n542), .A3(new_n613), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n491), .A2(new_n619), .A3(new_n540), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT75), .B1(new_n621), .B2(new_n612), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n449), .B1(new_n620), .B2(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n445), .A2(new_n446), .ZN(new_n625));
  INV_X1    g0425(.A(new_n413), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n447), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n425), .A2(new_n442), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n625), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n413), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n346), .B1(new_n283), .B2(new_n316), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n448), .A2(new_n358), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n625), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n624), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n600), .A2(new_n610), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n526), .A2(new_n539), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n512), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n619), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n569), .A2(KEYINPUT17), .A3(new_n594), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT17), .B1(new_n569), .B2(new_n594), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT85), .B1(new_n639), .B2(new_n619), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n489), .A2(new_n490), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n482), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n636), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(KEYINPUT87), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n273), .A2(KEYINPUT27), .A3(G20), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n273), .B2(G20), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G343), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n283), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n358), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n650), .B1(new_n283), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n317), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n317), .A2(new_n655), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n331), .A2(new_n655), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n346), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT86), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n352), .A2(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n346), .A2(KEYINPUT86), .A3(new_n665), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n346), .A2(new_n654), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n660), .B1(new_n659), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n210), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n432), .A2(new_n434), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n323), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n215), .B2(new_n680), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n385), .A2(new_n393), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n303), .A2(new_n444), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT88), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT88), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n303), .A2(new_n691), .A3(new_n444), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n341), .A2(new_n688), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n444), .B(KEYINPUT89), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n303), .B2(new_n312), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n687), .A4(new_n340), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n693), .B2(new_n694), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n655), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT31), .B(new_n655), .C1(new_n695), .C2(new_n699), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n702), .B(new_n703), .C1(new_n449), .C2(new_n655), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n633), .A2(new_n634), .ZN(new_n707));
  INV_X1    g0507(.A(new_n625), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n631), .A2(KEYINPUT91), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(new_n627), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n655), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n635), .A2(new_n654), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n706), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n686), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n670), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT92), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n671), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G13), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n680), .A2(G1), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n719), .B2(new_n720), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n213), .B1(G20), .B2(new_n333), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT96), .Z(new_n734));
  NOR2_X1   g0534(.A1(new_n678), .A2(new_n469), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G355), .B1(new_n323), .B2(new_n678), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n678), .A2(new_n250), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G45), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n216), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n239), .A2(G45), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n741), .B(new_n742), .C1(KEYINPUT93), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n743), .A2(KEYINPUT93), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n736), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n734), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n747), .B2(new_n746), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n315), .A2(new_n347), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n207), .A2(new_n349), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n347), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G50), .A2(new_n753), .B1(new_n756), .B2(G87), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G97), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n750), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n469), .B1(new_n764), .B2(G68), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n757), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n762), .A2(new_n758), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n315), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G77), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n751), .A2(new_n772), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n762), .A2(new_n754), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G58), .A2(new_n777), .B1(new_n779), .B2(G107), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n766), .A2(new_n771), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT98), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n778), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n752), .A2(new_n787), .B1(new_n755), .B2(new_n336), .ZN(new_n788));
  INV_X1    g0588(.A(new_n767), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n786), .B(new_n788), .C1(G329), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n776), .A2(new_n791), .B1(new_n773), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n250), .B(new_n793), .C1(new_n764), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n295), .A2(new_n296), .ZN(new_n796));
  INV_X1    g0596(.A(new_n760), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n790), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n783), .A2(new_n784), .A3(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n726), .B(new_n749), .C1(new_n732), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n668), .A2(new_n669), .A3(new_n731), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n722), .A2(new_n728), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n512), .A2(new_n654), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT100), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n498), .A2(new_n654), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n507), .A2(new_n508), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n498), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n804), .B(new_n805), .C1(new_n808), .C2(new_n512), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n511), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n333), .B1(new_n500), .B2(new_n505), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n499), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n509), .B2(new_n806), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n805), .B1(new_n814), .B2(new_n804), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n714), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n727), .B1(new_n817), .B2(new_n706), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n706), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n732), .A2(new_n729), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT99), .Z(new_n821));
  OAI21_X1  g0621(.A(new_n727), .B1(new_n821), .B2(G77), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n755), .A2(new_n275), .B1(new_n767), .B2(new_n792), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n250), .B(new_n823), .C1(G87), .C2(new_n779), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G294), .A2(new_n777), .B1(new_n774), .B2(G116), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G303), .A2(new_n753), .B1(new_n764), .B2(G283), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n824), .A2(new_n761), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n250), .B1(new_n755), .B2(new_n202), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n779), .A2(G68), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n767), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n828), .B(new_n831), .C1(G58), .C2(new_n760), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G137), .A2(new_n753), .B1(new_n774), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n776), .C1(new_n835), .C2(new_n763), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n827), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n822), .B1(new_n841), .B2(new_n732), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n816), .B2(new_n730), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n819), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  INV_X1    g0645(.A(G58), .ZN(new_n846));
  OAI21_X1  g0646(.A(G77), .B1(new_n846), .B2(new_n527), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n847), .A2(new_n215), .B1(G50), .B2(new_n527), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(G1), .A3(new_n723), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n214), .A2(G116), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT35), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n399), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n851), .B2(new_n399), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT36), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n624), .A2(new_n713), .A3(new_n716), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n624), .A2(new_n713), .A3(new_n859), .A4(new_n716), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n648), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT104), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n619), .A2(KEYINPUT101), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT101), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n864), .B(new_n538), .C1(new_n617), .C2(new_n618), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n655), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n599), .A2(new_n594), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT102), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n606), .A2(new_n871), .A3(new_n598), .A4(new_n609), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n606), .A2(new_n653), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n595), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n653), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n599), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n581), .A2(new_n583), .A3(new_n586), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n589), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n572), .B1(new_n588), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n877), .A2(new_n881), .B1(new_n594), .B2(new_n569), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n872), .A2(new_n875), .B1(new_n882), .B2(new_n869), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n876), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n612), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT39), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n873), .A2(new_n595), .A3(new_n874), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n606), .A2(new_n598), .A3(new_n609), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT37), .B1(new_n891), .B2(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n595), .A3(new_n874), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n890), .A2(new_n892), .B1(KEYINPUT37), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n874), .B1(new_n637), .B2(new_n643), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n868), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n653), .B1(new_n609), .B2(new_n598), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n595), .B1(new_n901), .B2(new_n880), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n890), .A2(new_n892), .B1(KEYINPUT37), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n884), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n637), .B2(new_n643), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n889), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n898), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n635), .A2(new_n816), .A3(new_n654), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n804), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n539), .A2(new_n654), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n526), .B2(new_n539), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n863), .A2(new_n911), .A3(new_n865), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n619), .A2(new_n654), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n907), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n637), .A2(new_n653), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n900), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n862), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n814), .A2(new_n804), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n809), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n912), .B2(new_n913), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n704), .B(new_n923), .C1(new_n886), .C2(new_n887), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n704), .A2(new_n914), .A3(new_n816), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n919), .B1(new_n896), .B2(new_n898), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n919), .A2(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n624), .A2(new_n704), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(G330), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n918), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n206), .B2(new_n724), .C1(new_n918), .C2(new_n931), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n856), .B1(new_n934), .B2(new_n935), .ZN(G367));
  NOR2_X1   g0736(.A1(new_n662), .A2(new_n674), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n396), .B(new_n413), .C1(new_n383), .C2(new_n654), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n626), .A2(new_n655), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT42), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n937), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n317), .B1(new_n942), .B2(new_n943), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n949), .A2(KEYINPUT107), .A3(new_n626), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT107), .B1(new_n949), .B2(new_n626), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n654), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n946), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n442), .A2(new_n654), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n625), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n447), .B2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n952), .A2(new_n948), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n961), .A2(new_n957), .A3(new_n956), .A4(new_n946), .ZN(new_n962));
  INV_X1    g0762(.A(new_n944), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n673), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n960), .B2(new_n962), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n679), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(new_n673), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT44), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n676), .B2(new_n944), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n676), .A2(new_n944), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n676), .A2(new_n970), .A3(new_n944), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n981), .A2(KEYINPUT108), .A3(new_n971), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n969), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n717), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n671), .A2(new_n662), .A3(new_n674), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n671), .B1(new_n662), .B2(new_n674), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n986), .A2(new_n987), .B1(KEYINPUT109), .B2(new_n937), .ZN(new_n988));
  INV_X1    g0788(.A(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n937), .A2(KEYINPUT109), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n990), .A3(new_n985), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n984), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n972), .A2(new_n973), .B1(new_n977), .B2(new_n978), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n981), .A2(KEYINPUT108), .A3(new_n971), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n673), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n983), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n968), .B1(new_n996), .B2(new_n717), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n725), .A2(G1), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n967), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n235), .A2(new_n738), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n734), .B1(new_n210), .B2(new_n438), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n727), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G97), .A2(new_n779), .B1(new_n774), .B2(G283), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n792), .B2(new_n752), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT46), .B1(new_n755), .B2(new_n323), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n323), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT110), .B(G317), .Z(new_n1008));
  OAI21_X1  g0808(.A(new_n469), .B1(new_n1008), .B2(new_n767), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n796), .A2(new_n763), .B1(new_n776), .B2(new_n336), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G107), .C2(new_n760), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n752), .A2(new_n834), .B1(new_n776), .B2(new_n835), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n763), .A2(new_n768), .B1(new_n773), .B2(new_n202), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G77), .A2(new_n779), .B1(new_n789), .B2(G137), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n760), .A2(G68), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n469), .B1(new_n756), .B2(G58), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1007), .A2(new_n1011), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT47), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n732), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1019), .B2(KEYINPUT47), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1002), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n956), .A2(new_n731), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n999), .A2(new_n1025), .ZN(G387));
  AOI22_X1  g0826(.A1(G322), .A2(new_n753), .B1(new_n774), .B2(G303), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n792), .B2(new_n763), .C1(new_n776), .C2(new_n1008), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT112), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1030), .A2(KEYINPUT48), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(KEYINPUT48), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n797), .A2(new_n785), .B1(new_n796), .B2(new_n755), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT49), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n469), .B1(new_n767), .B2(new_n787), .C1(new_n323), .C2(new_n778), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G50), .A2(new_n777), .B1(new_n789), .B2(G150), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n250), .C1(new_n321), .C2(new_n778), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n763), .A2(new_n451), .B1(new_n773), .B2(new_n527), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n752), .A2(new_n768), .B1(new_n755), .B2(new_n400), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n797), .A2(new_n438), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n732), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n683), .A2(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n683), .A2(KEYINPUT111), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n451), .A2(G50), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g0848(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n737), .C1(new_n739), .C2(new_n231), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n735), .A2(new_n682), .B1(new_n275), .B2(new_n678), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n726), .B1(new_n1053), .B2(new_n734), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1044), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n662), .B2(new_n731), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n991), .A2(new_n988), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n998), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n992), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n679), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1057), .A2(new_n717), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  NAND3_X1  g0862(.A1(new_n983), .A2(new_n995), .A3(new_n998), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n755), .A2(new_n527), .B1(new_n767), .B2(new_n834), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n469), .B(new_n1064), .C1(G87), .C2(new_n779), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT114), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n752), .A2(new_n835), .B1(new_n776), .B2(new_n768), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n760), .A2(G77), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n764), .B1(new_n774), .B2(new_n570), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n469), .B1(new_n778), .B2(new_n275), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G283), .A2(new_n756), .B1(new_n789), .B2(G322), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n294), .B2(new_n773), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT115), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n764), .A2(G303), .B1(new_n760), .B2(G116), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1072), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G317), .A2(new_n753), .B1(new_n777), .B2(G311), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  OAI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1021), .B1(new_n1071), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n734), .B1(new_n321), .B2(new_n210), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n738), .A2(new_n242), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n727), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT113), .Z(new_n1085));
  AOI211_X1 g0885(.A(new_n1081), .B(new_n1085), .C1(new_n963), .C2(new_n731), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n996), .A2(new_n679), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n983), .A2(new_n995), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1059), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G390));
  NAND2_X1  g0893(.A1(new_n896), .A2(new_n898), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n712), .A2(new_n816), .B1(new_n512), .B2(new_n654), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n914), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n868), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n804), .B2(new_n908), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n888), .B(new_n899), .C1(new_n1098), .C2(new_n867), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n706), .A2(new_n923), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n624), .A2(G330), .A3(new_n704), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n858), .A2(new_n648), .A3(new_n860), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n712), .A2(new_n816), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n804), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1096), .B1(new_n705), .B2(new_n922), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1100), .A3(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1100), .A2(new_n1109), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n909), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1104), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1103), .A2(new_n1113), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n679), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1103), .A2(new_n998), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n888), .A2(new_n729), .A3(new_n899), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n727), .B1(new_n821), .B2(new_n570), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n755), .A2(new_n835), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT116), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1122), .B1(new_n773), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G128), .A2(new_n753), .B1(new_n777), .B2(G132), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G137), .A2(new_n764), .B1(new_n789), .B2(G125), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n760), .A2(G159), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n469), .B1(new_n779), .B2(G50), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G116), .A2(new_n777), .B1(new_n789), .B2(G294), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n275), .B2(new_n763), .C1(new_n785), .C2(new_n752), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n250), .B1(new_n756), .B2(G87), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n774), .A2(G97), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1134), .A2(new_n829), .A3(new_n1069), .A4(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1126), .A2(new_n1131), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1120), .B1(new_n1137), .B2(new_n732), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1119), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1117), .A2(new_n1118), .A3(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(new_n1106), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1116), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n900), .A2(new_n916), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n915), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1147));
  NOR2_X1   g0947(.A1(new_n459), .A2(new_n876), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n491), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n491), .A2(new_n1149), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1147), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1152), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1147), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n928), .B2(G330), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n886), .A2(new_n887), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n919), .B1(new_n1159), .B2(new_n925), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1094), .A2(KEYINPUT40), .A3(new_n704), .A4(new_n923), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(G330), .A4(new_n1157), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1146), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1160), .A2(G330), .A3(new_n1161), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1157), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n917), .A3(new_n1162), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1143), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n680), .B1(new_n1142), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1106), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT119), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  AOI221_X4 g0974(.A(new_n1174), .B1(new_n1144), .B2(new_n1145), .C1(new_n1167), .C2(new_n1162), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1167), .A2(new_n1162), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT120), .B1(new_n1176), .B2(new_n1146), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1173), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1164), .A2(new_n1174), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(KEYINPUT120), .A3(new_n1146), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1171), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1170), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1166), .A2(new_n729), .ZN(new_n1186));
  INV_X1    g0986(.A(G137), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n763), .A2(new_n830), .B1(new_n773), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  INV_X1    g0989(.A(G128), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n752), .A2(new_n1189), .B1(new_n776), .B2(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1188), .B(new_n1191), .C1(G150), .C2(new_n760), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n755), .B2(new_n1125), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  INV_X1    g0995(.A(G41), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n372), .B(new_n1196), .C1(new_n778), .C2(new_n768), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT117), .B(G124), .Z(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n789), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1194), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n400), .A2(new_n755), .B1(new_n763), .B2(new_n321), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n752), .A2(new_n323), .B1(new_n778), .B2(new_n846), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n469), .A2(new_n1196), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G107), .B2(new_n777), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n773), .A2(new_n438), .B1(new_n767), .B2(new_n785), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1016), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G50), .B1(new_n372), .B2(new_n1196), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1208), .A2(new_n1209), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1200), .B(new_n1211), .C1(new_n1209), .C2(new_n1208), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n732), .B1(new_n1212), .B2(KEYINPUT118), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(KEYINPUT118), .B2(new_n1212), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n726), .B(new_n1214), .C1(new_n202), .C2(new_n820), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1185), .A2(new_n998), .B1(new_n1186), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1184), .A2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT121), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n968), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n1114), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1110), .B(new_n998), .C1(new_n1111), .C2(new_n909), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n727), .B1(new_n821), .B2(G68), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n752), .A2(new_n830), .B1(new_n776), .B2(new_n1187), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n469), .B(new_n1224), .C1(G58), .C2(new_n779), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n760), .A2(G50), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1124), .A2(new_n764), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n755), .A2(new_n768), .B1(new_n767), .B2(new_n1190), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G150), .B2(new_n774), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n469), .B1(new_n778), .B2(new_n400), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n323), .A2(new_n763), .B1(new_n776), .B2(new_n785), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1042), .A2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G97), .A2(new_n756), .B1(new_n789), .B2(G303), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G294), .A2(new_n753), .B1(new_n774), .B2(G107), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1223), .B1(new_n1238), .B2(new_n732), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n914), .B2(new_n730), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1222), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1221), .A2(new_n1242), .ZN(G381));
  NOR2_X1   g1043(.A1(G375), .A2(G378), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1092), .A2(new_n999), .A3(new_n1025), .ZN(new_n1246));
  OR3_X1    g1046(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G381), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(G407));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND2_X1  g1049(.A1(G387), .A2(G390), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(G393), .B(G396), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1250), .A2(new_n1246), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1250), .B2(new_n1246), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G378), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1180), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1142), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n968), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1164), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1168), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n998), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1186), .A2(new_n1215), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1256), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1184), .A2(G378), .A3(new_n1216), .ZN(new_n1267));
  INV_X1    g1067(.A(G343), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1266), .A2(new_n1267), .B1(G213), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT121), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT121), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1218), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT60), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n679), .B1(new_n1218), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1280), .B2(new_n1242), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n844), .B(new_n1241), .C1(new_n1276), .C2(new_n1279), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1269), .A2(new_n1270), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1268), .A2(G213), .A3(G2897), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1268), .A2(G213), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1287), .A2(KEYINPUT124), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1283), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1278), .B1(new_n1219), .B2(new_n1275), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n844), .B1(new_n1290), .B2(new_n1241), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1280), .A2(G384), .A3(new_n1242), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1288), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1286), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1284), .B(new_n1285), .C1(new_n1269), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1298), .A2(new_n1287), .A3(new_n1283), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(new_n1270), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1255), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1296), .B1(KEYINPUT123), .B2(new_n1269), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1269), .A2(KEYINPUT123), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1254), .A2(new_n1285), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1299), .B2(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1269), .A2(new_n1283), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1304), .A2(new_n1306), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1301), .A2(new_n1310), .ZN(G405));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1283), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1184), .A2(G378), .A3(new_n1216), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G378), .B1(new_n1184), .B2(new_n1216), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1312), .B(new_n1313), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1169), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n679), .B1(new_n1317), .B2(new_n1171), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n1259), .B2(new_n1143), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1185), .A2(new_n998), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1264), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1256), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1312), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1291), .A2(new_n1292), .A3(KEYINPUT125), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1322), .A2(new_n1267), .A3(new_n1323), .A4(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1316), .A2(new_n1254), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1316), .A2(new_n1325), .A3(new_n1254), .A4(KEYINPUT127), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1316), .A2(new_n1325), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT126), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1331), .A2(new_n1255), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1255), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(KEYINPUT126), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1330), .A2(new_n1333), .A3(new_n1335), .ZN(G402));
endmodule


