//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI211_X1 g003(.A(new_n204), .B(KEYINPUT89), .C1(G1gat), .C2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(G8gat), .Z(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT86), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT15), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT87), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(new_n212), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n216), .A2(new_n210), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT17), .B1(new_n221), .B2(KEYINPUT88), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n209), .A2(new_n213), .B1(new_n219), .B2(new_n215), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n206), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n206), .A2(new_n223), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n223), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n228), .B(KEYINPUT13), .Z(new_n234));
  AOI22_X1  g033(.A1(new_n230), .A2(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n227), .A2(new_n229), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n228), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G113gat), .B(G141gat), .Z(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G169gat), .B(G197gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT12), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OR3_X1    g044(.A1(new_n238), .A2(KEYINPUT90), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT90), .B1(new_n238), .B2(new_n245), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n246), .A2(new_n247), .B1(new_n238), .B2(new_n245), .ZN(new_n248));
  XOR2_X1   g047(.A(G1gat), .B(G29gat), .Z(new_n249));
  XNOR2_X1  g048(.A(G57gat), .B(G85gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n255), .A2(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(G134gat), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n254), .A2(KEYINPUT1), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(G113gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G120gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G155gat), .B(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT2), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(KEYINPUT73), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT2), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n278), .A3(new_n271), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  INV_X1    g079(.A(new_n272), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n275), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n268), .B1(new_n284), .B2(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n281), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n275), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(KEYINPUT75), .A3(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n258), .A2(new_n266), .A3(new_n275), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n282), .B2(new_n283), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT4), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(KEYINPUT76), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n305), .B(new_n297), .C1(new_n282), .C2(new_n283), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n296), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT5), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n284), .A2(new_n267), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(new_n310), .A3(new_n306), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n311), .B2(new_n301), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n253), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n305), .B1(new_n289), .B2(new_n297), .ZN(new_n315));
  INV_X1    g114(.A(new_n306), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT4), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n304), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n304), .B1(new_n303), .B2(new_n306), .ZN(new_n320));
  INV_X1    g119(.A(new_n318), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n320), .A2(KEYINPUT78), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n294), .B2(new_n295), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT79), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n317), .A2(new_n314), .A3(new_n318), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT78), .B1(new_n320), .B2(new_n321), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n285), .A2(KEYINPUT75), .A3(new_n291), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT75), .B1(new_n285), .B2(new_n291), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n324), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n313), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n253), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n330), .B2(new_n333), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n326), .A2(KEYINPUT79), .A3(new_n329), .A4(new_n328), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n308), .A2(new_n312), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT83), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n343), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n253), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT6), .B1(new_n342), .B2(new_n313), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT22), .ZN(new_n354));
  NAND2_X1  g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n352), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G211gat), .A2(G218gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(G211gat), .A2(G218gat), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT68), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  INV_X1    g160(.A(G218gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n353), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n366), .A2(new_n351), .B1(new_n357), .B2(KEYINPUT22), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT68), .B1(new_n357), .B2(new_n358), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n360), .A3(new_n355), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(KEYINPUT69), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT69), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n367), .A2(new_n372), .A3(new_n368), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(KEYINPUT70), .A3(new_n373), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G226gat), .ZN(new_n379));
  INV_X1    g178(.A(G233gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT23), .ZN(new_n383));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  AND4_X1   g185(.A1(KEYINPUT25), .A2(new_n383), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G183gat), .ZN(new_n388));
  INV_X1    g187(.A(G190gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT24), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(G183gat), .A3(G190gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n399));
  NOR2_X1   g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n390), .B2(new_n392), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n394), .B2(new_n395), .ZN(new_n406));
  NOR2_X1   g205(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n389), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT27), .B(G183gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(G190gat), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n382), .A2(KEYINPUT26), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n388), .B2(new_n389), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n384), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(new_n382), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n404), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n381), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n411), .ZN(new_n423));
  AND2_X1   g222(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT27), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n407), .ZN(new_n427));
  AOI21_X1  g226(.A(G190gat), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n428), .B2(KEYINPUT28), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n429), .A2(new_n418), .B1(new_n398), .B2(new_n403), .ZN(new_n430));
  INV_X1    g229(.A(new_n381), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n378), .B1(new_n422), .B2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n371), .A2(KEYINPUT70), .A3(new_n373), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT70), .B1(new_n371), .B2(new_n373), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n430), .B2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n381), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT71), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n436), .A2(new_n437), .A3(new_n438), .A4(KEYINPUT71), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n439), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT38), .B1(new_n450), .B2(KEYINPUT37), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(new_n442), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT72), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n446), .B1(new_n441), .B2(new_n442), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(KEYINPUT6), .B2(new_n344), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n345), .A2(new_n350), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT84), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n345), .A2(new_n350), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n449), .B1(new_n465), .B2(new_n453), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n466), .A2(KEYINPUT38), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n296), .A2(new_n329), .A3(new_n328), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n301), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT39), .C1(new_n301), .C2(new_n311), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n473), .A3(new_n301), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n474), .A2(new_n475), .A3(new_n339), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n474), .B2(new_n339), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT40), .B(new_n472), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n455), .A2(new_n482), .A3(new_n458), .ZN(new_n483));
  INV_X1    g282(.A(new_n447), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n456), .B2(KEYINPUT30), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n344), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G228gat), .A2(G233gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT80), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n291), .A2(new_n421), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n378), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n365), .B2(new_n370), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n284), .B1(KEYINPUT3), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n291), .A2(new_n421), .B1(new_n376), .B2(new_n377), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n284), .A2(new_n421), .A3(new_n373), .A4(new_n371), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n498));
  INV_X1    g297(.A(new_n488), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(G22gat), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n492), .A2(new_n498), .A3(new_n499), .A4(new_n497), .ZN(new_n503));
  INV_X1    g302(.A(new_n494), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n489), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G22gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT81), .ZN(new_n508));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT31), .B(G50gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  NAND4_X1  g310(.A1(new_n502), .A2(new_n507), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n508), .A3(new_n507), .ZN(new_n513));
  INV_X1    g312(.A(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n508), .B1(new_n502), .B2(new_n507), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n487), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n469), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n483), .A2(new_n485), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n347), .A2(new_n349), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n344), .A2(KEYINPUT6), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n420), .A2(new_n267), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n430), .A2(new_n268), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G227gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n380), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT66), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT34), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT32), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT33), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G15gat), .B(G43gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT65), .ZN(new_n541));
  INV_X1    g340(.A(G71gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G99gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n537), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n537), .B1(new_n539), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n535), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n539), .A2(new_n546), .ZN(new_n551));
  INV_X1    g350(.A(new_n537), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(new_n533), .A3(new_n534), .A4(new_n547), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(KEYINPUT36), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n550), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n535), .B(KEYINPUT67), .C1(new_n548), .C2(new_n549), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n525), .A2(new_n518), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n521), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n523), .A2(new_n524), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n517), .B1(new_n561), .B2(new_n560), .ZN(new_n567));
  INV_X1    g366(.A(new_n522), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n345), .A2(new_n524), .A3(new_n350), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n483), .A2(new_n572), .A3(new_n485), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n573), .A2(new_n517), .A3(new_n555), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n248), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  INV_X1    g380(.A(G92gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT94), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n222), .B2(new_n226), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n589), .B2(new_n223), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n389), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n588), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n587), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n221), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n225), .B1(new_n223), .B2(new_n224), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(G190gat), .B1(new_n600), .B2(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n362), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT93), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n595), .A2(new_n601), .A3(G218gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT95), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT93), .B1(new_n602), .B2(new_n362), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n611), .A3(new_n605), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n607), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n607), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n579), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n612), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n611), .B1(new_n610), .B2(new_n605), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n608), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n607), .A2(new_n609), .A3(new_n612), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n578), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G57gat), .B(G64gat), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G71gat), .B(G78gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n631), .B(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n206), .B1(new_n628), .B2(new_n627), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT92), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n637), .B(new_n640), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n589), .A2(new_n627), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n597), .A2(new_n626), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(G230gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n380), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(KEYINPUT96), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(KEYINPUT96), .A3(new_n647), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n649), .A2(new_n659), .A3(new_n654), .A4(new_n655), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n577), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n566), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n522), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n670), .A2(G8gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n673), .ZN(G1325gat));
  NOR3_X1   g474(.A1(new_n665), .A2(G15gat), .A3(new_n555), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n557), .A2(new_n562), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n666), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n676), .B1(G15gat), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT97), .Z(G1326gat));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n518), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n571), .A2(new_n574), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n572), .B1(new_n525), .B2(new_n567), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n570), .A2(new_n575), .A3(KEYINPUT101), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n467), .B1(new_n461), .B2(KEYINPUT84), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n519), .B1(new_n689), .B2(new_n464), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n687), .B(new_n688), .C1(new_n690), .C2(new_n563), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n615), .A2(new_n620), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n621), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n565), .B2(new_n576), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n641), .A2(new_n663), .ZN(new_n698));
  INV_X1    g497(.A(new_n248), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT100), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n693), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n667), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n217), .B1(new_n703), .B2(KEYINPUT102), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT102), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n692), .A2(new_n698), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT98), .Z(new_n707));
  NAND4_X1  g506(.A1(new_n707), .A2(new_n217), .A3(new_n667), .A4(new_n577), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT99), .B(KEYINPUT45), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n710), .ZN(G1328gat));
  NAND4_X1  g510(.A1(new_n707), .A2(new_n218), .A3(new_n522), .A4(new_n577), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT46), .Z(new_n713));
  AND2_X1   g512(.A1(new_n702), .A2(new_n522), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n218), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT103), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n713), .B(new_n717), .C1(new_n218), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n707), .A2(new_n720), .A3(new_n556), .A4(new_n577), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT104), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n702), .A2(new_n677), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1330gat));
  NAND2_X1  g525(.A1(new_n687), .A2(new_n688), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n563), .B1(new_n469), .B2(new_n520), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n692), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n694), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n565), .A2(new_n576), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n695), .ZN(new_n732));
  INV_X1    g531(.A(new_n701), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n730), .A2(new_n517), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G50gat), .ZN(new_n735));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n707), .A2(new_n736), .A3(new_n517), .A4(new_n577), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(KEYINPUT48), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  INV_X1    g538(.A(new_n737), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n735), .B2(KEYINPUT105), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n742), .A3(G50gat), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n739), .B(KEYINPUT48), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  NOR4_X1   g543(.A1(new_n693), .A2(new_n697), .A3(new_n518), .A4(new_n701), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT105), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n743), .A3(new_n737), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT106), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n738), .B1(new_n744), .B2(new_n749), .ZN(G1331gat));
  INV_X1    g549(.A(new_n691), .ZN(new_n751));
  INV_X1    g550(.A(new_n663), .ZN(new_n752));
  NOR4_X1   g551(.A1(new_n751), .A2(new_n699), .A3(new_n642), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n667), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g554(.A(new_n568), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT107), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n758), .B(new_n759), .Z(G1333gat));
  AOI21_X1  g559(.A(new_n542), .B1(new_n753), .B2(new_n677), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n555), .A2(G71gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n753), .A2(new_n517), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n693), .A2(new_n697), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n699), .A2(new_n641), .A3(new_n752), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(KEYINPUT108), .A3(new_n667), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n566), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(G85gat), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n729), .A2(new_n699), .A3(new_n641), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT51), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n667), .A2(new_n581), .A3(new_n663), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NAND4_X1  g578(.A1(new_n776), .A2(new_n582), .A3(new_n522), .A4(new_n663), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n769), .B2(new_n568), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n784), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n677), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G99gat), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n752), .A2(new_n555), .A3(G99gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n777), .B2(new_n789), .ZN(G1338gat));
  OAI21_X1  g589(.A(G106gat), .B1(new_n769), .B2(new_n518), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n752), .A2(new_n518), .A3(G106gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(KEYINPUT109), .A2(KEYINPUT53), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT109), .A2(KEYINPUT53), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT110), .ZN(new_n796));
  AND4_X1   g595(.A1(new_n791), .A2(new_n793), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n776), .A2(new_n792), .B1(KEYINPUT109), .B2(KEYINPUT53), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n791), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n799), .ZN(G1339gat));
  AND4_X1   g599(.A1(new_n248), .A2(new_n621), .A3(new_n641), .A4(new_n752), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n246), .A2(new_n247), .ZN(new_n802));
  INV_X1    g601(.A(new_n243), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n236), .A2(new_n228), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n233), .A2(new_n234), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n651), .A2(new_n647), .A3(new_n652), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n809));
  AOI21_X1  g608(.A(new_n659), .B1(new_n653), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n662), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(new_n808), .B2(new_n810), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n802), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n615), .A3(new_n620), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n815), .A2(new_n615), .A3(new_n818), .A4(new_n620), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n663), .A3(new_n806), .ZN(new_n820));
  INV_X1    g619(.A(new_n814), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n248), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n621), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n817), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n641), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n801), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n517), .A3(new_n555), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n667), .A3(new_n568), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n261), .A3(new_n248), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n825), .ZN(new_n830));
  INV_X1    g629(.A(new_n801), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n567), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n522), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n667), .A3(new_n834), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(new_n248), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n829), .B1(new_n261), .B2(new_n836), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n828), .B2(new_n752), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n663), .A2(new_n259), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT113), .Z(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n835), .B2(new_n840), .ZN(G1341gat));
  NOR3_X1   g640(.A1(new_n828), .A2(new_n255), .A3(new_n825), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT114), .B1(new_n835), .B2(new_n825), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n825), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G127gat), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(G1342gat));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n828), .B2(new_n621), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n621), .A2(G134gat), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n667), .A3(new_n834), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT56), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT116), .B1(new_n850), .B2(KEYINPUT56), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n847), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n851), .B(KEYINPUT115), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n857), .A2(new_n858), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT117), .A4(new_n848), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n677), .A2(new_n518), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n667), .A2(new_n832), .A3(new_n568), .A4(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(G141gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n699), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n677), .A2(new_n566), .A3(new_n522), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT118), .Z(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n826), .B2(new_n518), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n816), .A2(KEYINPUT112), .B1(new_n621), .B2(new_n822), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n641), .B1(new_n874), .B2(new_n819), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n517), .C1(new_n875), .C2(new_n801), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n248), .B(new_n871), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n873), .A2(new_n876), .ZN(new_n880));
  INV_X1    g679(.A(new_n871), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(KEYINPUT120), .A3(new_n248), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n865), .B(new_n869), .C1(new_n879), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n869), .B1(new_n877), .B2(new_n868), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT58), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n885), .B2(KEYINPUT58), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n663), .A3(new_n881), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(KEYINPUT59), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n890), .B2(new_n893), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n641), .B1(new_n823), .B2(new_n816), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n517), .B1(new_n897), .B2(new_n801), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n872), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n876), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n871), .A2(new_n752), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n892), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n894), .A2(new_n895), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n867), .A2(new_n892), .A3(new_n663), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n882), .B2(new_n825), .ZN(new_n906));
  INV_X1    g705(.A(G155gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n867), .A2(new_n907), .A3(new_n641), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1346gat));
  INV_X1    g708(.A(G162gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n867), .A2(new_n910), .A3(new_n692), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n882), .A2(new_n621), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  OAI21_X1  g712(.A(G162gat), .B1(new_n912), .B2(KEYINPUT122), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n826), .A2(new_n667), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n833), .A2(new_n568), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n699), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n667), .A2(new_n568), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n827), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G169gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n922), .A2(new_n923), .A3(new_n248), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n920), .A2(new_n924), .ZN(G1348gat));
  NAND4_X1  g724(.A1(new_n827), .A2(G176gat), .A3(new_n663), .A4(new_n921), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT123), .ZN(new_n927));
  AOI21_X1  g726(.A(G176gat), .B1(new_n919), .B2(new_n663), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(KEYINPUT123), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G1349gat));
  NAND3_X1  g729(.A1(new_n919), .A2(new_n410), .A3(new_n641), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n922), .A2(new_n825), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n424), .A2(new_n425), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n922), .B2(new_n621), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(KEYINPUT61), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n938), .A2(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n919), .A2(new_n389), .A3(new_n692), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(G1351gat));
  NAND3_X1  g741(.A1(new_n916), .A2(new_n522), .A3(new_n866), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(G197gat), .A3(new_n248), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT125), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n667), .A2(new_n677), .A3(new_n568), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n900), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n248), .ZN(new_n948));
  OAI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(KEYINPUT126), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(KEYINPUT126), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  NOR3_X1   g750(.A1(new_n943), .A2(G204gat), .A3(new_n752), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n947), .B2(new_n752), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1353gat));
  OR3_X1    g754(.A1(new_n943), .A2(G211gat), .A3(new_n825), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n947), .A2(new_n825), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(new_n361), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(KEYINPUT63), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n947), .B2(new_n621), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n692), .A2(new_n362), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n943), .B2(new_n963), .ZN(G1355gat));
endmodule


