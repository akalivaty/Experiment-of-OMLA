//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n462), .B2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n479), .B2(G2105), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT72), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n471), .B1(new_n466), .B2(KEYINPUT71), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n461), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n483), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(new_n461), .A2(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n476), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n484), .B2(new_n485), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n488), .B2(G126), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n504), .B1(new_n509), .B2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n505), .A2(new_n506), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT74), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n517), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n515), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT75), .B(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n507), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT76), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT76), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n510), .B2(new_n512), .ZN(new_n538));
  AND2_X1   g113(.A1(G77), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT77), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n513), .A2(G90), .A3(new_n514), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n507), .A2(G52), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n545), .B(G651), .C1(new_n538), .C2(new_n539), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT78), .A4(new_n546), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AOI22_X1  g127(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G651), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n513), .A2(new_n514), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT80), .B(G43), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(G81), .B1(new_n507), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  AND2_X1   g141(.A1(new_n513), .A2(G65), .ZN(new_n567));
  AND2_X1   g142(.A1(G78), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n557), .A2(G91), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n507), .A2(new_n572), .A3(G53), .ZN(new_n573));
  AND2_X1   g148(.A1(KEYINPUT6), .A2(G651), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  OAI211_X1 g150(.A(G53), .B(G543), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(new_n529), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT76), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n533), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT81), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n580), .B(new_n584), .C1(new_n581), .C2(new_n533), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  NAND2_X1  g163(.A1(new_n557), .A2(G87), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n507), .A2(G49), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  AOI22_X1  g167(.A1(new_n557), .A2(G86), .B1(G48), .B2(new_n507), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n510), .A2(new_n512), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n593), .A2(new_n598), .A3(KEYINPUT82), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT82), .B1(new_n593), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(G651), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n557), .A2(G85), .B1(G47), .B2(new_n507), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G171), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n557), .A2(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n595), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n615), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  AOI211_X1 g192(.A(KEYINPUT84), .B(new_n609), .C1(new_n608), .C2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(KEYINPUT84), .B2(new_n609), .ZN(G284));
  XNOR2_X1  g194(.A(G284), .B(KEYINPUT85), .ZN(G321));
  NOR2_X1   g195(.A1(G299), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n586), .ZN(G297));
  AOI21_X1  g197(.A(new_n621), .B1(G868), .B2(new_n586), .ZN(G280));
  INV_X1    g198(.A(new_n617), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n476), .A2(new_n467), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT13), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n486), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n488), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n461), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n634), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT88), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT87), .B(G2438), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n643), .B(new_n644), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(new_n647), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n651), .A3(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND4_X1  g235(.A1(new_n649), .A2(new_n651), .A3(KEYINPUT14), .A4(new_n655), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n657), .B2(new_n661), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT89), .ZN(G401));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT90), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n671), .A2(KEYINPUT91), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(KEYINPUT91), .ZN(new_n673));
  INV_X1    g248(.A(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n669), .B(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n672), .B(new_n673), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n667), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n667), .A2(new_n670), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT92), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n695), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT20), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n692), .A2(new_n693), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n689), .B(KEYINPUT19), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n694), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT93), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n698), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1991), .B(G1996), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n698), .A2(new_n701), .A3(new_n706), .A4(new_n708), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n712), .B1(new_n710), .B2(new_n713), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n688), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n718), .A2(new_n687), .A3(new_n714), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(G229));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G32), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT26), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G105), .B2(new_n467), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n486), .A2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n488), .A2(G129), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT99), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(G16), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n561), .B2(new_n738), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1341), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(G20), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT23), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n571), .A2(new_n578), .ZN(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT101), .B(G1956), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n736), .B(new_n741), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT31), .B(G11), .Z(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n722), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n639), .B2(new_n722), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n486), .A2(G139), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n755), .B(new_n756), .C1(new_n461), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n722), .A2(G33), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n753), .B1(new_n762), .B2(G2072), .ZN(new_n763));
  INV_X1    g338(.A(G2072), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n761), .A2(new_n764), .B1(new_n733), .B2(new_n734), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G27), .A2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G164), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n770), .C1(new_n747), .C2(new_n748), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT96), .Z(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n617), .B2(new_n745), .ZN(new_n774));
  INV_X1    g349(.A(G1348), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G34), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT24), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n722), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G160), .B2(new_n722), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2084), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n771), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G5), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G171), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n722), .A2(G35), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT100), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n490), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT29), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n745), .A2(G21), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G168), .B2(new_n745), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1966), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n722), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n488), .A2(G128), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT97), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n486), .B2(G140), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(G29), .ZN(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n793), .A2(new_n796), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n749), .A2(new_n783), .A3(new_n787), .A4(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G6), .B(G305), .S(G16), .Z(new_n812));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n814), .A2(new_n817), .A3(new_n815), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n738), .A2(G22), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n738), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n745), .A2(G23), .ZN(new_n825));
  INV_X1    g400(.A(G288), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n745), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT33), .B(G1976), .Z(new_n828));
  XOR2_X1   g403(.A(new_n827), .B(new_n828), .Z(new_n829));
  NAND4_X1  g404(.A1(new_n819), .A2(new_n820), .A3(new_n824), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G24), .B(G290), .S(new_n738), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1986), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n722), .A2(G25), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n486), .A2(G131), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n488), .A2(G119), .ZN(new_n837));
  OR2_X1    g412(.A1(G95), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n835), .B1(new_n840), .B2(new_n722), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G1991), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n834), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n830), .B2(KEYINPUT34), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT36), .B1(new_n832), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n831), .A4(new_n845), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n811), .B1(new_n847), .B2(new_n850), .ZN(G311));
  INV_X1    g426(.A(G311), .ZN(G150));
  NAND2_X1  g427(.A1(new_n624), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT102), .B(G55), .Z(new_n855));
  AOI22_X1  g430(.A1(new_n557), .A2(G93), .B1(new_n507), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n518), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n560), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n854), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(G145));
  NAND2_X1  g443(.A1(new_n486), .A2(G142), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n488), .A2(G130), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n461), .A2(KEYINPUT107), .A3(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT107), .B1(new_n461), .B2(G118), .ZN(new_n872));
  OR2_X1    g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n871), .A2(G2104), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n632), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n840), .A2(KEYINPUT108), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n876), .B1(new_n877), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n877), .A2(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n632), .ZN(new_n886));
  INV_X1    g461(.A(new_n875), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n502), .B(new_n731), .Z(new_n890));
  INV_X1    g465(.A(new_n806), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n502), .B(new_n731), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n806), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT106), .B1(new_n758), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(KEYINPUT106), .B2(new_n758), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(new_n897), .A3(new_n894), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n889), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G160), .B(new_n639), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G162), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n889), .A3(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n908), .B2(new_n901), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g487(.A(new_n859), .B(new_n627), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n744), .A2(new_n617), .ZN(new_n914));
  NAND3_X1  g489(.A1(G299), .A2(new_n612), .A3(new_n616), .ZN(new_n915));
  XOR2_X1   g490(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n915), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n913), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n913), .A2(new_n919), .ZN(new_n923));
  OR3_X1    g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT42), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n826), .B1(new_n605), .B2(new_n606), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n605), .A2(new_n826), .A3(new_n606), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT110), .B1(new_n930), .B2(new_n925), .ZN(new_n931));
  OAI21_X1  g506(.A(G166), .B1(new_n599), .B2(new_n600), .ZN(new_n932));
  NAND2_X1  g507(.A1(G305), .A2(G303), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n929), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n932), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(new_n927), .A3(new_n926), .A4(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT42), .B1(new_n922), .B2(new_n923), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n924), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n924), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n858), .A2(new_n608), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(G331));
  NAND3_X1  g520(.A1(new_n549), .A2(G168), .A3(new_n550), .ZN(new_n946));
  OAI211_X1 g521(.A(KEYINPUT111), .B(new_n946), .C1(G301), .C2(new_n586), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(KEYINPUT111), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n947), .A2(new_n859), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n859), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n919), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  INV_X1    g527(.A(new_n859), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n921), .A2(new_n918), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(new_n859), .A3(new_n948), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n957), .A3(new_n938), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n910), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n938), .B1(new_n951), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n914), .A2(new_n915), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n920), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n954), .A2(new_n964), .A3(new_n956), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n954), .B2(new_n956), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n937), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n910), .A4(new_n958), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n910), .A3(new_n958), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n974), .B2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n951), .A2(new_n957), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n937), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(new_n968), .A3(new_n910), .A4(new_n958), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n973), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n954), .A2(new_n964), .A3(new_n956), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n938), .B1(new_n980), .B2(new_n951), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n959), .B2(new_n981), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n973), .A2(new_n982), .A3(KEYINPUT44), .A4(new_n978), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n972), .B1(new_n979), .B2(new_n983), .ZN(G397));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n497), .B2(new_n501), .ZN(new_n987));
  OAI211_X1 g562(.A(G160), .B(G40), .C1(new_n987), .C2(KEYINPUT45), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n989), .B(G1384), .C1(new_n497), .C2(new_n501), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n823), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  INV_X1    g567(.A(new_n492), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n463), .B2(new_n464), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n994), .A2(KEYINPUT4), .B1(new_n476), .B2(new_n493), .ZN(new_n995));
  OAI211_X1 g570(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n996));
  INV_X1    g571(.A(new_n500), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n992), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n473), .A2(new_n474), .B1(G113), .B2(G2104), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n461), .B1(new_n1001), .B2(new_n477), .ZN(new_n1002));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n469), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n987), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n991), .B1(G2090), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1008), .B2(KEYINPUT117), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n792), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1012), .B2(new_n991), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n986), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n986), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(KEYINPUT114), .A3(new_n991), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(G8), .ZN(new_n1019));
  INV_X1    g594(.A(G1981), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n593), .A2(new_n598), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n593), .B2(new_n598), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT115), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1004), .B2(new_n987), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT115), .B(new_n1028), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1027), .B(new_n1032), .C1(new_n1031), .C2(G288), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1027), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G288), .A2(new_n1031), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT52), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n988), .B2(new_n990), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .A4(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1026), .B(G286), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1014), .A2(new_n1019), .A3(new_n1038), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT63), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(KEYINPUT118), .A3(new_n1045), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1037), .B(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1043), .A2(KEYINPUT63), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1016), .A2(new_n1018), .A3(G8), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n986), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(new_n1019), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1049), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1030), .A2(new_n1031), .A3(new_n826), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1034), .B1(new_n1057), .B2(new_n1021), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1019), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1040), .A2(G168), .A3(new_n1042), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(G168), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1066), .A3(G8), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n999), .A2(new_n989), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1004), .A3(new_n1071), .A4(new_n769), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT126), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1073), .A2(KEYINPUT53), .B1(new_n786), .B2(new_n1007), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(KEYINPUT126), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1068), .A2(new_n1069), .A3(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1074), .A2(G301), .A3(new_n1076), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT125), .B1(new_n1080), .B2(new_n1077), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT125), .B(KEYINPUT54), .C1(new_n1080), .C2(new_n1077), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1087));
  AOI21_X1  g662(.A(new_n572), .B1(new_n507), .B2(G53), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT120), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n573), .A2(new_n577), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(new_n569), .A3(new_n570), .A4(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(KEYINPUT121), .A3(new_n1094), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1097), .A2(new_n1098), .B1(new_n744), .B2(KEYINPUT57), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1070), .A2(new_n1004), .A3(new_n1071), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1011), .B2(G1956), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n479), .A2(G2105), .ZN(new_n1105));
  INV_X1    g680(.A(new_n469), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(G40), .A3(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1104), .A2(new_n990), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1108), .A2(new_n1100), .B1(new_n1007), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n571), .A2(KEYINPUT57), .A3(new_n578), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1093), .A2(KEYINPUT121), .A3(new_n1094), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT121), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1087), .B1(new_n1103), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1099), .A2(new_n1102), .A3(KEYINPUT122), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1007), .A2(new_n775), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1004), .A2(new_n808), .A3(new_n987), .ZN(new_n1124));
  AND4_X1   g699(.A1(KEYINPUT60), .A2(new_n1123), .A3(new_n617), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1996), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1070), .A2(new_n1004), .A3(new_n1071), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1107), .B2(new_n999), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1130), .A2(new_n561), .B1(new_n1131), .B2(KEYINPUT59), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n560), .B(new_n1133), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1125), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n617), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1137), .B2(new_n1136), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1116), .A2(new_n1122), .A3(new_n1135), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n624), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1118), .A2(new_n1121), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1086), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1079), .B1(new_n1085), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1014), .A2(new_n1019), .A3(new_n1038), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1056), .B(new_n1060), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1070), .A2(new_n1107), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1126), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(new_n731), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1148), .B(KEYINPUT113), .Z(new_n1151));
  XNOR2_X1  g726(.A(new_n806), .B(G2067), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n732), .A2(new_n1126), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1150), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n878), .B(new_n843), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(G290), .B(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1148), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1147), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1151), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1155), .A2(new_n842), .A3(new_n840), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n891), .A2(new_n808), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1152), .A2(new_n731), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT47), .Z(new_n1169));
  INV_X1    g744(.A(new_n1158), .ZN(new_n1170));
  NOR2_X1   g745(.A1(G290), .A2(G1986), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1148), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1165), .B(new_n1169), .C1(new_n1170), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1161), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n685), .B(G319), .C1(new_n663), .C2(new_n664), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n719), .B2(new_n717), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n1179), .A2(new_n911), .ZN(new_n1180));
  AOI211_X1 g754(.A(new_n1177), .B(new_n1180), .C1(new_n961), .C2(new_n969), .ZN(new_n1181));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1182));
  AOI21_X1  g756(.A(KEYINPUT127), .B1(new_n970), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1183), .ZN(G308));
  NAND2_X1  g758(.A1(new_n970), .A2(new_n1182), .ZN(G225));
endmodule


