//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT66), .A2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G143), .A3(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n189), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT66), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT66), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n193), .B1(new_n200), .B2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n189), .A2(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n195), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G104), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT80), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n207), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT3), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(KEYINPUT80), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n208), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n187), .B1(new_n205), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n220), .B1(new_n213), .B2(new_n215), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n214), .A2(KEYINPUT3), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n208), .B1(new_n210), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n219), .A3(KEYINPUT4), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n192), .A2(KEYINPUT0), .A3(G128), .A4(new_n194), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n195), .A3(KEYINPUT64), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(KEYINPUT0), .B2(G128), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n232), .A2(new_n234), .B1(KEYINPUT0), .B2(G128), .ZN(new_n235));
  AOI21_X1  g049(.A(G143), .B1(new_n190), .B2(new_n191), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G146), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n189), .A2(KEYINPUT65), .A3(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n235), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G101), .C1(new_n225), .C2(new_n227), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n229), .A2(new_n230), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(new_n246), .B2(G134), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G137), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT11), .B1(new_n249), .B2(G137), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n246), .A3(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n251), .B2(new_n256), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n225), .A2(new_n227), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n221), .B1(new_n260), .B2(new_n218), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n236), .A2(new_n241), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n195), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n197), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n264), .A3(KEYINPUT10), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n224), .A2(new_n245), .A3(new_n259), .A4(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(G227), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n224), .A2(new_n245), .A3(new_n265), .ZN(new_n274));
  INV_X1    g088(.A(new_n259), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n266), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT81), .B1(new_n261), .B2(new_n264), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n261), .A2(new_n204), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n198), .A2(new_n199), .A3(new_n238), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n282));
  OAI21_X1  g096(.A(G128), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n239), .B(new_n240), .C1(new_n200), .C2(G143), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n283), .A2(new_n284), .B1(new_n201), .B2(new_n196), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n223), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n280), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n275), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n278), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(G469), .B(new_n277), .C1(new_n293), .C2(new_n271), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n272), .B1(new_n291), .B2(new_n292), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n271), .B1(new_n276), .B2(new_n266), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n295), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n295), .A2(new_n296), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G221), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT9), .B(G234), .Z(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(new_n296), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G113), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G119), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT5), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G116), .B(G119), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(new_n315), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT2), .A2(G113), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n312), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n223), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n219), .A2(new_n319), .A3(new_n326), .A4(new_n222), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G122), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT8), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n283), .A2(new_n284), .ZN(new_n334));
  AOI21_X1  g148(.A(G125), .B1(new_n334), .B2(new_n197), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n242), .A2(G125), .A3(new_n230), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n268), .A2(G224), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT7), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n338), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n264), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n242), .A2(G125), .A3(new_n230), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT82), .B(new_n333), .C1(new_n339), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n324), .ZN(new_n346));
  NOR3_X1   g160(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n346), .A2(new_n347), .B1(new_n322), .B2(new_n312), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT70), .A3(new_n318), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT70), .B1(new_n325), .B2(new_n317), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n318), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n229), .A2(new_n349), .A3(new_n352), .A4(new_n244), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n331), .A3(new_n329), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n345), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n338), .B1(new_n335), .B2(new_n336), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n342), .A2(new_n343), .A3(new_n340), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT82), .B1(new_n358), .B2(new_n333), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n296), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n329), .ZN(new_n361));
  INV_X1    g175(.A(new_n331), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n354), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n342), .A2(new_n343), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n337), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(new_n367), .A3(new_n362), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n311), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n358), .A2(new_n333), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n354), .A3(new_n345), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n374), .A2(new_n296), .A3(new_n310), .A4(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n309), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G478), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT15), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n313), .A2(KEYINPUT14), .A3(G122), .ZN(new_n380));
  INV_X1    g194(.A(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n313), .A2(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(G107), .B(new_n380), .C1(new_n384), .C2(KEYINPUT14), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n383), .A3(new_n206), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n238), .A2(G128), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n195), .A2(G143), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n249), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n249), .B1(new_n387), .B2(new_n388), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n385), .B(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(G107), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n386), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT13), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n395), .B(G134), .C1(KEYINPUT13), .C2(new_n387), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n396), .A3(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n304), .A2(G217), .A3(new_n268), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n296), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n379), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n405), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(KEYINPUT88), .A3(new_n296), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n409), .B2(new_n379), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT86), .B(G475), .Z(new_n412));
  INV_X1    g226(.A(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n341), .A2(G140), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT16), .ZN(new_n416));
  OR3_X1    g230(.A1(new_n341), .A2(KEYINPUT16), .A3(G140), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(G146), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n189), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT76), .A4(G146), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(G237), .A2(G953), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G214), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n238), .ZN(new_n428));
  AND2_X1   g242(.A1(KEYINPUT83), .A2(G143), .ZN(new_n429));
  NOR2_X1   g243(.A1(KEYINPUT83), .A2(G143), .ZN(new_n430));
  OAI211_X1 g244(.A(G214), .B(new_n425), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G131), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n431), .A3(new_n252), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n252), .B1(new_n428), .B2(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n424), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(new_n252), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G125), .B(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n200), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT79), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT79), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n200), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n444), .A2(new_n189), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n440), .B(new_n443), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT85), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT84), .B(G104), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n439), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n439), .A2(new_n451), .ZN(new_n458));
  INV_X1    g272(.A(new_n455), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI211_X1 g274(.A(KEYINPUT87), .B(new_n455), .C1(new_n439), .C2(new_n451), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n412), .B1(new_n462), .B2(new_n296), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  INV_X1    g278(.A(new_n435), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(new_n437), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT19), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n444), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n200), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n418), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n450), .B1(new_n446), .B2(new_n448), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n441), .B(new_n252), .C1(new_n428), .C2(new_n431), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n432), .A2(new_n442), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n459), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n456), .ZN(new_n477));
  NOR2_X1   g291(.A1(G475), .A2(G902), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  AOI211_X1 g294(.A(KEYINPUT20), .B(new_n480), .C1(new_n476), .C2(new_n456), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n268), .A2(G952), .ZN(new_n483));
  NAND2_X1  g297(.A1(G234), .A2(G237), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(G902), .A3(G953), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT21), .B(G898), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR4_X1   g304(.A1(new_n411), .A2(new_n463), .A3(new_n482), .A4(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n307), .A2(new_n377), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n425), .A2(G210), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n493), .B(KEYINPUT27), .Z(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n246), .A2(G134), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n249), .A2(G137), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n252), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT68), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n264), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n230), .B(new_n242), .C1(new_n257), .C2(new_n258), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n352), .A2(new_n349), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT72), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n499), .A2(new_n500), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n502), .B1(new_n513), .B2(new_n252), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n501), .A2(KEYINPUT68), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n498), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT71), .B1(new_n285), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n264), .A2(new_n518), .A3(new_n498), .A4(new_n503), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n517), .A2(new_n519), .A3(new_n506), .A4(new_n505), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n506), .B1(new_n504), .B2(new_n505), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n497), .B1(new_n512), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n519), .A3(new_n505), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT30), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n504), .A2(new_n505), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n506), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n521), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT31), .B1(new_n533), .B2(new_n497), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n506), .B1(new_n527), .B2(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n536));
  NOR4_X1   g350(.A1(new_n535), .A2(new_n536), .A3(new_n521), .A4(new_n496), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n525), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(G472), .A2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT32), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n529), .B1(KEYINPUT30), .B2(new_n526), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n520), .B(new_n497), .C1(new_n542), .C2(new_n506), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n531), .A2(new_n532), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n545), .A2(KEYINPUT31), .A3(new_n520), .A4(new_n497), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n524), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n539), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n541), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n511), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n509), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n526), .A2(new_n532), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n508), .B1(new_n552), .B2(new_n520), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n496), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n512), .A2(new_n523), .A3(new_n497), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n496), .B1(new_n535), .B2(new_n521), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G472), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n540), .A2(new_n549), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G119), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT74), .B1(new_n564), .B2(G128), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT23), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT74), .B(new_n567), .C1(new_n564), .C2(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(G128), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT78), .B(G110), .ZN(new_n571));
  XNOR2_X1  g385(.A(G119), .B(G128), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT24), .B(G110), .Z(new_n573));
  OAI22_X1  g387(.A1(new_n570), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n446), .A2(new_n448), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n418), .ZN(new_n576));
  INV_X1    g390(.A(G110), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n570), .B2(KEYINPUT75), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n566), .A2(new_n579), .A3(new_n568), .A4(new_n569), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n578), .A2(new_n580), .B1(new_n572), .B2(new_n573), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT77), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G110), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n573), .A2(new_n572), .ZN(new_n586));
  AND4_X1   g400(.A1(KEYINPUT77), .A2(new_n585), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n576), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  INV_X1    g403(.A(G234), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n303), .A2(new_n590), .A3(G953), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n576), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n585), .A2(new_n582), .A3(new_n586), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n581), .A2(KEYINPUT77), .A3(new_n582), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n592), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G217), .B1(new_n590), .B2(G902), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT73), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n593), .A2(new_n601), .A3(new_n296), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT25), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n593), .A2(new_n601), .A3(KEYINPUT25), .A4(new_n296), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n607), .B1(new_n612), .B2(new_n604), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n492), .A2(new_n563), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT89), .B(G101), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G3));
  NAND2_X1  g430(.A1(KEYINPUT90), .A2(G472), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n538), .A2(new_n296), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n617), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n547), .B2(G902), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n490), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n377), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n399), .B2(KEYINPUT91), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n402), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n401), .B1(new_n392), .B2(new_n397), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n400), .A2(new_n402), .A3(new_n626), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n296), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G478), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n403), .A2(new_n378), .A3(new_n296), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n463), .A2(new_n482), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n624), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n613), .A2(new_n306), .A3(new_n302), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n622), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n412), .ZN(new_n644));
  INV_X1    g458(.A(new_n456), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n458), .A2(new_n459), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT87), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n458), .A2(new_n457), .A3(new_n459), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n644), .B1(new_n649), .B2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT94), .ZN(new_n651));
  AOI211_X1 g465(.A(KEYINPUT93), .B(new_n464), .C1(new_n477), .C2(new_n478), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n482), .B2(KEYINPUT93), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT94), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n463), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n651), .A2(new_n653), .A3(new_n655), .A4(new_n411), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n624), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n622), .A2(new_n657), .A3(new_n640), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT95), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n599), .A2(new_n662), .ZN(new_n663));
  AOI211_X1 g477(.A(KEYINPUT95), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n664));
  OAI22_X1  g478(.A1(new_n663), .A2(new_n664), .B1(KEYINPUT36), .B2(new_n592), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n588), .A2(KEYINPUT95), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n599), .A2(new_n662), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n592), .A2(KEYINPUT36), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n612), .A2(new_n604), .B1(new_n670), .B2(new_n605), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n661), .B1(new_n621), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n612), .A2(new_n604), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n605), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n618), .A2(new_n675), .A3(new_n620), .A4(KEYINPUT96), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n492), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n486), .B1(new_n488), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n656), .A2(new_n671), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(new_n563), .A3(new_n307), .A4(new_n377), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XOR2_X1   g498(.A(new_n681), .B(KEYINPUT39), .Z(new_n685));
  AND2_X1   g499(.A1(new_n307), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n688));
  OR3_X1    g502(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT40), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT40), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  INV_X1    g504(.A(G472), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n552), .A2(new_n520), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n692), .B2(new_n496), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n543), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(G472), .A2(G902), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT97), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n540), .A3(new_n549), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n370), .A2(new_n376), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT38), .Z(new_n701));
  OAI21_X1  g515(.A(new_n650), .B1(new_n479), .B2(new_n481), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n410), .A2(new_n309), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n699), .A2(new_n701), .A3(new_n675), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n689), .A2(new_n690), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR3_X1   g521(.A1(new_n671), .A2(new_n638), .A3(new_n681), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n563), .A2(new_n708), .A3(new_n307), .A4(new_n377), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(new_n291), .A2(new_n292), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n298), .B1(new_n711), .B2(new_n273), .ZN(new_n712));
  OAI21_X1  g526(.A(G469), .B1(new_n712), .B2(G902), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n306), .A3(new_n299), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT99), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(KEYINPUT99), .A3(new_n306), .A4(new_n299), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n563), .A2(new_n613), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n639), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  AND3_X1   g535(.A1(new_n540), .A2(new_n549), .A3(new_n562), .ZN(new_n722));
  INV_X1    g536(.A(new_n613), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n716), .A2(new_n717), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n657), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT100), .B(G116), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G18));
  AND3_X1   g542(.A1(new_n713), .A2(new_n306), .A3(new_n299), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n675), .A3(new_n377), .A4(new_n491), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT101), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n377), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n732), .A2(new_n671), .A3(new_n714), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n563), .A4(new_n491), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  AND4_X1   g551(.A1(new_n700), .A2(new_n702), .A3(new_n703), .A4(new_n623), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n716), .A3(new_n717), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n496), .B1(new_n554), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT102), .ZN(new_n742));
  OAI22_X1  g556(.A1(new_n741), .A2(new_n742), .B1(new_n534), .B2(new_n537), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n539), .ZN(new_n744));
  OAI21_X1  g558(.A(G472), .B1(new_n547), .B2(G902), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n613), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n381), .ZN(G24));
  NOR2_X1   g562(.A1(new_n638), .A2(new_n681), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n538), .A2(new_n296), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n750), .A2(G472), .B1(new_n743), .B2(new_n539), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n733), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NAND2_X1  g567(.A1(new_n302), .A2(KEYINPUT103), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n370), .A2(new_n308), .A3(new_n376), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n294), .A2(new_n299), .A3(new_n756), .A4(new_n301), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n306), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT104), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n305), .B1(new_n302), .B2(KEYINPUT103), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n755), .A4(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n724), .A3(new_n749), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n759), .A2(new_n762), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n549), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(KEYINPUT105), .B(new_n541), .C1(new_n547), .C2(new_n548), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n540), .A3(new_n562), .A4(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n638), .A2(new_n765), .A3(new_n681), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n613), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT106), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n771), .A2(new_n613), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n763), .A4(new_n772), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n766), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NOR2_X1   g593(.A1(new_n656), .A2(new_n681), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n763), .A2(new_n724), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT107), .B(G134), .Z(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(G36));
  NOR2_X1   g597(.A1(new_n636), .A2(new_n637), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n702), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT43), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n621), .A4(new_n675), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n755), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT109), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n787), .B2(new_n755), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n786), .A2(new_n621), .A3(new_n675), .ZN(new_n792));
  OAI22_X1  g606(.A1(new_n789), .A2(new_n791), .B1(KEYINPUT44), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n277), .B1(new_n293), .B2(new_n271), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n295), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n796), .B(KEYINPUT108), .C1(new_n795), .C2(new_n794), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n300), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n299), .B1(new_n801), .B2(KEYINPUT46), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n306), .A3(new_n685), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n793), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT110), .B(G137), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G39));
  NAND3_X1  g622(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n306), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n306), .B1(new_n802), .B2(new_n803), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n722), .A2(new_n723), .A3(new_n749), .A4(new_n755), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  AND2_X1   g630(.A1(new_n713), .A2(new_n299), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT49), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n613), .A2(new_n785), .A3(new_n306), .A4(new_n308), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n699), .A2(new_n818), .A3(new_n701), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  INV_X1    g635(.A(new_n702), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n411), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n638), .ZN(new_n824));
  INV_X1    g638(.A(new_n624), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n622), .A2(new_n824), .A3(new_n825), .A4(new_n640), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n677), .A2(new_n614), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n736), .A2(new_n726), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n725), .A2(new_n563), .A3(new_n613), .ZN(new_n829));
  INV_X1    g643(.A(new_n639), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n829), .A2(new_n830), .B1(new_n746), .B2(new_n739), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n828), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n735), .A2(new_n731), .B1(new_n718), .B2(new_n657), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n747), .B1(new_n718), .B2(new_n639), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT111), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n827), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n683), .A2(new_n752), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n760), .A2(new_n757), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n681), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n698), .A3(new_n671), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n838), .A2(KEYINPUT52), .A3(new_n709), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n683), .A3(new_n752), .A4(new_n709), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n744), .A2(new_n749), .A3(new_n745), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n759), .B2(new_n762), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n411), .A2(new_n681), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n655), .A2(new_n850), .A3(new_n651), .A4(new_n653), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n563), .A2(new_n307), .A3(new_n755), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n675), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n781), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n847), .A2(new_n854), .A3(new_n778), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n821), .B1(new_n837), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT112), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n821), .C1(new_n837), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n828), .A2(new_n831), .A3(new_n821), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n847), .A2(new_n862), .A3(new_n778), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n827), .A2(new_n853), .A3(new_n781), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(KEYINPUT113), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(KEYINPUT113), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n861), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n837), .A2(new_n855), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n856), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n786), .A2(new_n486), .ZN(new_n875));
  INV_X1    g689(.A(new_n746), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n714), .A2(new_n308), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n701), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT50), .Z(new_n879));
  INV_X1    g693(.A(new_n755), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n714), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n786), .A2(new_n486), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n675), .A3(new_n751), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n613), .A2(new_n699), .A3(new_n486), .A4(new_n881), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n822), .A3(new_n784), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n879), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n817), .A2(new_n305), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n809), .A2(new_n812), .A3(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n875), .A2(new_n876), .A3(new_n755), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n888), .B2(KEYINPUT114), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n638), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n875), .A2(new_n377), .A3(new_n729), .A4(new_n876), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n483), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT48), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n882), .A2(new_n775), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT117), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n892), .B2(new_n894), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n874), .A2(new_n895), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(G952), .A2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n820), .B1(new_n909), .B2(new_n910), .ZN(G75));
  NOR2_X1   g725(.A1(new_n268), .A2(G952), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT119), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n867), .B1(new_n857), .B2(new_n859), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n296), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(G210), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n364), .A2(new_n368), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(new_n366), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n917), .A2(new_n918), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(G210), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n915), .A2(new_n926), .A3(new_n296), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n923), .B1(new_n927), .B2(KEYINPUT56), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n914), .B1(new_n925), .B2(new_n928), .ZN(G51));
  XNOR2_X1  g743(.A(new_n300), .B(KEYINPUT57), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n861), .B1(new_n860), .B2(new_n868), .ZN(new_n931));
  AOI211_X1 g745(.A(KEYINPUT54), .B(new_n867), .C1(new_n857), .C2(new_n859), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n712), .B(KEYINPUT120), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n916), .A2(new_n799), .A3(new_n800), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n912), .B1(new_n935), .B2(new_n936), .ZN(G54));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n916), .A2(new_n477), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n477), .B1(new_n916), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n912), .ZN(G60));
  AND2_X1   g755(.A1(new_n630), .A2(new_n631), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT59), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n874), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n860), .A2(new_n868), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT54), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n869), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n945), .A2(new_n949), .A3(new_n914), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n947), .A2(new_n670), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n602), .B1(new_n915), .B2(new_n952), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n913), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n954), .A2(new_n955), .A3(new_n913), .A4(new_n957), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  INV_X1    g775(.A(G224), .ZN(new_n962));
  OAI21_X1  g776(.A(G953), .B1(new_n489), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n837), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(G953), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n919), .B1(G898), .B2(new_n268), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  XNOR2_X1  g781(.A(new_n542), .B(KEYINPUT122), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n468), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n775), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n840), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n804), .A2(new_n972), .A3(new_n306), .A4(new_n685), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n838), .A2(new_n709), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n781), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n973), .B(new_n975), .C1(new_n793), .C2(new_n805), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n778), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n813), .B2(new_n814), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n680), .A2(G953), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT125), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n985));
  INV_X1    g799(.A(new_n979), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n268), .B1(new_n986), .B2(new_n976), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n985), .B1(new_n987), .B2(new_n982), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n970), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n268), .B1(G227), .B2(G900), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n706), .A2(new_n974), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT123), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n880), .B1(new_n824), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n823), .A2(KEYINPUT123), .A3(new_n638), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n724), .A2(new_n996), .A3(new_n686), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n806), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n994), .A2(new_n815), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n970), .B1(new_n1001), .B2(new_n268), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n989), .A2(new_n991), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT126), .B1(new_n980), .B2(new_n983), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n987), .A2(new_n985), .A3(new_n982), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n969), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n990), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1004), .A2(new_n1008), .ZN(G72));
  XNOR2_X1  g823(.A(new_n695), .B(KEYINPUT63), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1010), .B1(new_n559), .B2(new_n543), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n872), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1001), .A2(new_n837), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1013), .A2(new_n1010), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n497), .B1(new_n535), .B2(new_n521), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n912), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n986), .A2(new_n976), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1010), .B1(new_n1018), .B2(new_n964), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n533), .A2(new_n496), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1023), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1016), .B1(new_n1022), .B2(new_n1024), .ZN(G57));
endmodule


