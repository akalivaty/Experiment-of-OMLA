

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U562 ( .A1(n703), .A2(n702), .ZN(n747) );
  NOR2_X1 U563 ( .A1(n765), .A2(n808), .ZN(n766) );
  NAND2_X1 U564 ( .A1(n940), .A2(n799), .ZN(n526) );
  XOR2_X1 U565 ( .A(KEYINPUT109), .B(n815), .Z(n527) );
  OR2_X1 U566 ( .A1(KEYINPUT33), .A2(n766), .ZN(n528) );
  OR2_X1 U567 ( .A1(n715), .A2(n707), .ZN(n714) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n741) );
  NAND2_X1 U569 ( .A1(G8), .A2(n747), .ZN(n808) );
  NOR2_X1 U570 ( .A1(n800), .A2(n526), .ZN(n801) );
  NOR2_X1 U571 ( .A1(G651), .A2(n657), .ZN(n659) );
  XNOR2_X1 U572 ( .A(KEYINPUT15), .B(n596), .ZN(n901) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U574 ( .A1(n651), .A2(G85), .ZN(n531) );
  XNOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n529), .B(KEYINPUT67), .ZN(n657) );
  XOR2_X1 U577 ( .A(G651), .B(KEYINPUT68), .Z(n532) );
  NOR2_X2 U578 ( .A1(n657), .A2(n532), .ZN(n646) );
  NAND2_X1 U579 ( .A1(G72), .A2(n646), .ZN(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n537) );
  NAND2_X1 U581 ( .A1(n659), .A2(G47), .ZN(n535) );
  NOR2_X1 U582 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n533), .Z(n663) );
  NAND2_X1 U584 ( .A1(G60), .A2(n663), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U586 ( .A1(n537), .A2(n536), .ZN(G290) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U588 ( .A1(G113), .A2(n883), .ZN(n539) );
  INV_X1 U589 ( .A(G2105), .ZN(n540) );
  NOR2_X1 U590 ( .A1(G2104), .A2(n540), .ZN(n884) );
  NAND2_X1 U591 ( .A1(G125), .A2(n884), .ZN(n538) );
  AND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n695) );
  AND2_X1 U593 ( .A1(G2104), .A2(n540), .ZN(n541) );
  XNOR2_X2 U594 ( .A(n541), .B(KEYINPUT64), .ZN(n880) );
  NAND2_X1 U595 ( .A1(n880), .A2(G101), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n542), .B(KEYINPUT23), .ZN(n543) );
  XNOR2_X1 U597 ( .A(KEYINPUT65), .B(n543), .ZN(n547) );
  NOR2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT17), .B(n544), .Z(n879) );
  NAND2_X1 U600 ( .A1(G137), .A2(n879), .ZN(n545) );
  XNOR2_X1 U601 ( .A(n545), .B(KEYINPUT66), .ZN(n546) );
  AND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n696) );
  AND2_X1 U603 ( .A1(n695), .A2(n696), .ZN(G160) );
  NAND2_X1 U604 ( .A1(n659), .A2(G52), .ZN(n548) );
  XNOR2_X1 U605 ( .A(KEYINPUT69), .B(n548), .ZN(n556) );
  NAND2_X1 U606 ( .A1(n651), .A2(G90), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G77), .A2(n646), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT9), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT70), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G64), .A2(n663), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  NAND2_X1 U616 ( .A1(n651), .A2(G89), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G76), .A2(n646), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(KEYINPUT79), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n659), .A2(G51), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G63), .A2(n663), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U627 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G138), .A2(n879), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G102), .A2(n880), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G114), .A2(n883), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G126), .A2(n884), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n573), .A2(n572), .ZN(G164) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n834) );
  NAND2_X1 U639 ( .A1(n834), .A2(G567), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  XOR2_X1 U641 ( .A(KEYINPUT74), .B(KEYINPUT12), .Z(n577) );
  NAND2_X1 U642 ( .A1(G81), .A2(n651), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G68), .A2(n646), .ZN(n578) );
  XNOR2_X1 U645 ( .A(KEYINPUT75), .B(n578), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U647 ( .A(KEYINPUT13), .B(KEYINPUT76), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G56), .A2(n663), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT14), .B(n583), .Z(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n659), .A2(G43), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n935) );
  INV_X1 U654 ( .A(G860), .ZN(n636) );
  OR2_X1 U655 ( .A1(n935), .A2(n636), .ZN(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U658 ( .A1(G54), .A2(n659), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n588), .B(KEYINPUT78), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n651), .A2(G92), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G66), .A2(n663), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G79), .A2(n646), .ZN(n591) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(n591), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U667 ( .A(n901), .ZN(n931) );
  INV_X1 U668 ( .A(G868), .ZN(n667) );
  NAND2_X1 U669 ( .A1(n931), .A2(n667), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U671 ( .A1(n659), .A2(G53), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G65), .A2(n663), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT73), .B(n601), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n646), .A2(G78), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT72), .B(n602), .Z(n605) );
  NAND2_X1 U677 ( .A1(G91), .A2(n651), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT71), .B(n603), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(G299) );
  NOR2_X1 U681 ( .A1(G286), .A2(n667), .ZN(n609) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n636), .A2(G559), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n610), .A2(n901), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n935), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n901), .A2(G868), .ZN(n612) );
  NOR2_X1 U689 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(G282) );
  XOR2_X1 U691 ( .A(G2100), .B(KEYINPUT82), .Z(n625) );
  XOR2_X1 U692 ( .A(G2096), .B(KEYINPUT81), .Z(n623) );
  NAND2_X1 U693 ( .A1(G135), .A2(n879), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G111), .A2(n883), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G123), .A2(n884), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n617), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n880), .A2(G99), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n982) );
  XNOR2_X1 U702 ( .A(n623), .B(n982), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G55), .A2(n659), .ZN(n626) );
  XOR2_X1 U705 ( .A(KEYINPUT86), .B(n626), .Z(n631) );
  NAND2_X1 U706 ( .A1(n651), .A2(G93), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G80), .A2(n646), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT85), .B(n629), .Z(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G67), .A2(n663), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n669) );
  XNOR2_X1 U713 ( .A(n669), .B(KEYINPUT84), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n935), .B(KEYINPUT83), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n901), .A2(G559), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n635), .B(n634), .ZN(n675) );
  NAND2_X1 U717 ( .A1(n675), .A2(n636), .ZN(n637) );
  XNOR2_X1 U718 ( .A(n638), .B(n637), .ZN(G145) );
  NAND2_X1 U719 ( .A1(G88), .A2(n651), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G50), .A2(n659), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G75), .A2(n646), .ZN(n641) );
  XNOR2_X1 U723 ( .A(KEYINPUT91), .B(n641), .ZN(n642) );
  NOR2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G62), .A2(n663), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U727 ( .A(G303), .ZN(G166) );
  NAND2_X1 U728 ( .A1(n646), .A2(G73), .ZN(n647) );
  XNOR2_X1 U729 ( .A(n647), .B(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G48), .A2(n659), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT90), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G61), .A2(n663), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G86), .A2(n651), .ZN(n652) );
  XNOR2_X1 U735 ( .A(KEYINPUT89), .B(n652), .ZN(n653) );
  NOR2_X1 U736 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(G305) );
  NAND2_X1 U738 ( .A1(G87), .A2(n657), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(KEYINPUT88), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n659), .A2(G49), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U743 ( .A1(G74), .A2(G651), .ZN(n664) );
  XOR2_X1 U744 ( .A(KEYINPUT87), .B(n664), .Z(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(G288) );
  NAND2_X1 U746 ( .A1(n667), .A2(n669), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n668), .B(KEYINPUT92), .ZN(n678) );
  XNOR2_X1 U748 ( .A(G299), .B(n669), .ZN(n674) );
  XNOR2_X1 U749 ( .A(G166), .B(G305), .ZN(n672) );
  XOR2_X1 U750 ( .A(KEYINPUT19), .B(G290), .Z(n670) );
  XNOR2_X1 U751 ( .A(G288), .B(n670), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n674), .B(n673), .ZN(n900) );
  XNOR2_X1 U754 ( .A(n900), .B(n675), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G868), .A2(n676), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U757 ( .A(KEYINPUT93), .B(n679), .Z(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(KEYINPUT94), .Z(n680) );
  XNOR2_X1 U760 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G2090), .ZN(n683) );
  XOR2_X1 U762 ( .A(KEYINPUT95), .B(n683), .Z(n684) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U766 ( .A1(G132), .A2(G82), .ZN(n686) );
  XNOR2_X1 U767 ( .A(n686), .B(KEYINPUT96), .ZN(n687) );
  XNOR2_X1 U768 ( .A(n687), .B(KEYINPUT22), .ZN(n688) );
  NOR2_X1 U769 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G96), .A2(n689), .ZN(n838) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n838), .ZN(n693) );
  NAND2_X1 U772 ( .A1(G108), .A2(G120), .ZN(n690) );
  NOR2_X1 U773 ( .A1(G237), .A2(n690), .ZN(n691) );
  NAND2_X1 U774 ( .A1(G69), .A2(n691), .ZN(n839) );
  NAND2_X1 U775 ( .A1(G567), .A2(n839), .ZN(n692) );
  NAND2_X1 U776 ( .A1(n693), .A2(n692), .ZN(n840) );
  NAND2_X1 U777 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U778 ( .A1(n840), .A2(n694), .ZN(n837) );
  NAND2_X1 U779 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U780 ( .A(G1986), .B(G290), .ZN(n925) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n703) );
  AND2_X1 U782 ( .A1(n695), .A2(G40), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U784 ( .A1(n703), .A2(n698), .ZN(n829) );
  NAND2_X1 U785 ( .A1(n925), .A2(n829), .ZN(n816) );
  XOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .Z(n952) );
  INV_X1 U787 ( .A(n698), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n952), .A2(n747), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT103), .ZN(n701) );
  XOR2_X1 U790 ( .A(KEYINPUT102), .B(G1961), .Z(n997) );
  NAND2_X1 U791 ( .A1(n997), .A2(n747), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n738) );
  NAND2_X1 U793 ( .A1(n738), .A2(G171), .ZN(n732) );
  XNOR2_X1 U794 ( .A(KEYINPUT107), .B(KEYINPUT29), .ZN(n730) );
  AND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n720) );
  AND2_X1 U796 ( .A1(n720), .A2(G1996), .ZN(n704) );
  XOR2_X1 U797 ( .A(n704), .B(KEYINPUT26), .Z(n706) );
  NAND2_X1 U798 ( .A1(n747), .A2(G1341), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n715) );
  OR2_X1 U800 ( .A1(n931), .A2(n935), .ZN(n707) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n747), .ZN(n708) );
  XNOR2_X1 U802 ( .A(KEYINPUT104), .B(n708), .ZN(n711) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n720), .ZN(n709) );
  XOR2_X1 U804 ( .A(KEYINPUT105), .B(n709), .Z(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U806 ( .A(KEYINPUT106), .B(n712), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n935), .A2(n715), .ZN(n716) );
  OR2_X1 U809 ( .A1(n901), .A2(n716), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n724) );
  INV_X1 U811 ( .A(G299), .ZN(n928) );
  NAND2_X1 U812 ( .A1(n720), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U813 ( .A(n719), .B(KEYINPUT27), .ZN(n722) );
  INV_X1 U814 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U815 ( .A1(n998), .A2(n720), .ZN(n721) );
  NOR2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U817 ( .A1(n928), .A2(n725), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U819 ( .A1(n928), .A2(n725), .ZN(n726) );
  XOR2_X1 U820 ( .A(n726), .B(KEYINPUT28), .Z(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n744) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n747), .ZN(n756) );
  NOR2_X1 U825 ( .A1(n808), .A2(G1966), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n733), .B(KEYINPUT101), .ZN(n758) );
  NAND2_X1 U827 ( .A1(G8), .A2(n758), .ZN(n734) );
  NOR2_X1 U828 ( .A1(n756), .A2(n734), .ZN(n736) );
  INV_X1 U829 ( .A(KEYINPUT30), .ZN(n735) );
  XNOR2_X1 U830 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U831 ( .A1(G168), .A2(n737), .ZN(n740) );
  NOR2_X1 U832 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U834 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n757) );
  AND2_X1 U836 ( .A1(G286), .A2(G8), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n757), .A2(n745), .ZN(n754) );
  INV_X1 U838 ( .A(G8), .ZN(n752) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n808), .ZN(n746) );
  XNOR2_X1 U840 ( .A(n746), .B(KEYINPUT108), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n747), .A2(G2090), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n750), .A2(G303), .ZN(n751) );
  OR2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U846 ( .A(n755), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X1 U847 ( .A1(G8), .A2(n756), .ZN(n760) );
  AND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n804) );
  NOR2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n767), .A2(n763), .ZN(n929) );
  NAND2_X1 U854 ( .A1(n804), .A2(n929), .ZN(n764) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n926) );
  NAND2_X1 U856 ( .A1(n764), .A2(n926), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n767), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n808), .A2(n768), .ZN(n800) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n940) );
  NAND2_X1 U860 ( .A1(G131), .A2(n879), .ZN(n770) );
  NAND2_X1 U861 ( .A1(G95), .A2(n880), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U863 ( .A(KEYINPUT98), .B(n771), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G107), .A2(n883), .ZN(n773) );
  NAND2_X1 U865 ( .A1(G119), .A2(n884), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n892) );
  AND2_X1 U868 ( .A1(n892), .A2(G1991), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n883), .A2(G117), .ZN(n776) );
  XOR2_X1 U870 ( .A(KEYINPUT99), .B(n776), .Z(n778) );
  NAND2_X1 U871 ( .A1(n884), .A2(G129), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U873 ( .A(KEYINPUT100), .B(n779), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n880), .A2(G105), .ZN(n780) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n780), .Z(n781) );
  NOR2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n879), .A2(G141), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n868) );
  AND2_X1 U879 ( .A1(G1996), .A2(n868), .ZN(n785) );
  NOR2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n974) );
  INV_X1 U881 ( .A(n829), .ZN(n787) );
  NOR2_X1 U882 ( .A1(n974), .A2(n787), .ZN(n820) );
  INV_X1 U883 ( .A(n820), .ZN(n798) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NAND2_X1 U885 ( .A1(G104), .A2(n880), .ZN(n788) );
  XOR2_X1 U886 ( .A(KEYINPUT97), .B(n788), .Z(n790) );
  NAND2_X1 U887 ( .A1(n879), .A2(G140), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n791), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G116), .A2(n883), .ZN(n793) );
  NAND2_X1 U891 ( .A1(G128), .A2(n884), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n794), .Z(n795) );
  NOR2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n797), .ZN(n896) );
  NOR2_X1 U896 ( .A1(n826), .A2(n896), .ZN(n988) );
  NAND2_X1 U897 ( .A1(n829), .A2(n988), .ZN(n824) );
  NAND2_X1 U898 ( .A1(n798), .A2(n824), .ZN(n812) );
  INV_X1 U899 ( .A(n812), .ZN(n799) );
  NAND2_X1 U900 ( .A1(n528), .A2(n801), .ZN(n814) );
  NOR2_X1 U901 ( .A1(G2090), .A2(G303), .ZN(n802) );
  NAND2_X1 U902 ( .A1(G8), .A2(n802), .ZN(n803) );
  NAND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n805) );
  AND2_X1 U904 ( .A1(n805), .A2(n808), .ZN(n810) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XOR2_X1 U906 ( .A(n806), .B(KEYINPUT24), .Z(n807) );
  NOR2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n527), .ZN(n832) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n868), .ZN(n977) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n892), .A2(G1991), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n817), .B(KEYINPUT110), .ZN(n983) );
  NOR2_X1 U916 ( .A1(n818), .A2(n983), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n977), .A2(n821), .ZN(n822) );
  XOR2_X1 U919 ( .A(KEYINPUT111), .B(n822), .Z(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n826), .A2(n896), .ZN(n972) );
  NAND2_X1 U923 ( .A1(n827), .A2(n972), .ZN(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT112), .B(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  XOR2_X1 U933 ( .A(G120), .B(KEYINPUT114), .Z(G236) );
  INV_X1 U935 ( .A(G132), .ZN(G219) );
  INV_X1 U936 ( .A(G108), .ZN(G238) );
  INV_X1 U937 ( .A(G82), .ZN(G220) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U940 ( .A(KEYINPUT115), .B(n840), .ZN(G319) );
  XNOR2_X1 U941 ( .A(G1956), .B(KEYINPUT118), .ZN(n850) );
  XOR2_X1 U942 ( .A(G1976), .B(G1981), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1971), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U945 ( .A(G1961), .B(G1966), .Z(n844) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U948 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U949 ( .A(G2474), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT117), .B(G2678), .Z(n852) );
  XNOR2_X1 U953 ( .A(KEYINPUT116), .B(KEYINPUT43), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2090), .Z(n854) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U958 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2100), .B(G2096), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U961 ( .A(G2078), .B(G2084), .Z(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U963 ( .A1(G124), .A2(n884), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n883), .A2(G112), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G136), .A2(n879), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G100), .A2(n880), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U970 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U971 ( .A(G160), .B(n868), .Z(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(n982), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G118), .A2(n883), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G130), .A2(n884), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G142), .A2(n879), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G106), .A2(n880), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U981 ( .A(n878), .B(n877), .Z(n891) );
  NAND2_X1 U982 ( .A1(G139), .A2(n879), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G103), .A2(n880), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G115), .A2(n883), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G127), .A2(n884), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n967) );
  XNOR2_X1 U990 ( .A(G164), .B(n967), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n898) );
  XOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n894) );
  XOR2_X1 U993 ( .A(n892), .B(G162), .Z(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U998 ( .A(n900), .B(G286), .Z(n903) );
  XNOR2_X1 U999 ( .A(n901), .B(G171), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n904), .B(n935), .Z(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G397) );
  XOR2_X1 U1003 ( .A(G2454), .B(G2435), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G2438), .B(G2427), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n914) );
  XOR2_X1 U1006 ( .A(KEYINPUT113), .B(G2446), .Z(n909) );
  XNOR2_X1 U1007 ( .A(G2443), .B(G2430), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1009 ( .A(n910), .B(G2451), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n915), .A2(G14), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G96), .ZN(G221) );
  INV_X1 U1022 ( .A(G69), .ZN(G235) );
  INV_X1 U1023 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1024 ( .A(KEYINPUT56), .B(G16), .ZN(n946) );
  XNOR2_X1 U1025 ( .A(G171), .B(G1961), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(G1971), .A2(G303), .ZN(n922) );
  NAND2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1028 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n939) );
  XNOR2_X1 U1030 ( .A(n928), .B(G1956), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n934) );
  XOR2_X1 U1032 ( .A(G1348), .B(n931), .Z(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT125), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1035 ( .A(G1341), .B(n935), .Z(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G168), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(n942), .B(KEYINPUT57), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n947), .B(KEYINPUT126), .ZN(n966) );
  XNOR2_X1 U1044 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(n948), .B(KEYINPUT54), .ZN(n964) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n961) );
  XOR2_X1 U1047 ( .A(G25), .B(G1991), .Z(n949) );
  NAND2_X1 U1048 ( .A1(n949), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(G27), .B(n952), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1059 ( .A(KEYINPUT124), .B(n962), .Z(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n1021) );
  NAND2_X1 U1061 ( .A1(n1021), .A2(KEYINPUT55), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n1030) );
  XOR2_X1 U1063 ( .A(G2072), .B(n967), .Z(n969) );
  XOR2_X1 U1064 ( .A(G164), .B(G2078), .Z(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT122), .B(n970), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n971), .B(KEYINPUT50), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n991) );
  XNOR2_X1 U1069 ( .A(G160), .B(G2084), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n981) );
  XOR2_X1 U1071 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1073 ( .A(KEYINPUT120), .B(n978), .Z(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT51), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT119), .B(n984), .Z(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT121), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1082 ( .A(n992), .B(KEYINPUT52), .Z(n993) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n993), .ZN(n995) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n996), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1087 ( .A(n997), .B(G5), .ZN(n1011) );
  XNOR2_X1 U1088 ( .A(G20), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G6), .B(G1981), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n1006) );
  XOR2_X1 U1097 ( .A(n1007), .B(n1006), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1020), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(KEYINPUT55), .A2(G29), .ZN(n1023) );
  INV_X1 U1111 ( .A(n1021), .ZN(n1022) );
  NAND2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(G11), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1031), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

