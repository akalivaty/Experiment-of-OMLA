

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781;

  XNOR2_X1 U374 ( .A(n573), .B(n377), .ZN(n397) );
  XNOR2_X1 U375 ( .A(n736), .B(KEYINPUT6), .ZN(n582) );
  XNOR2_X1 U376 ( .A(n352), .B(n351), .ZN(n581) );
  INV_X1 U377 ( .A(n380), .ZN(n351) );
  XNOR2_X1 U378 ( .A(n362), .B(G110), .ZN(n436) );
  BUF_X1 U379 ( .A(n689), .Z(n350) );
  XNOR2_X2 U380 ( .A(n402), .B(n580), .ZN(n592) );
  INV_X1 U381 ( .A(n352), .ZN(n382) );
  OR2_X2 U382 ( .A1(n411), .A2(n414), .ZN(n352) );
  INV_X1 U383 ( .A(G128), .ZN(n468) );
  XNOR2_X1 U384 ( .A(n557), .B(n464), .ZN(n624) );
  XNOR2_X1 U385 ( .A(KEYINPUT107), .B(n550), .ZN(n353) );
  XOR2_X1 U386 ( .A(n559), .B(KEYINPUT38), .Z(n354) );
  NAND2_X2 U387 ( .A1(n440), .A2(n439), .ZN(n559) );
  NAND2_X1 U388 ( .A1(n397), .A2(n582), .ZN(n579) );
  XNOR2_X2 U389 ( .A(n516), .B(n465), .ZN(n768) );
  XNOR2_X2 U390 ( .A(n539), .B(n467), .ZN(n516) );
  NAND2_X1 U391 ( .A1(n358), .A2(n356), .ZN(n652) );
  NAND2_X1 U392 ( .A1(n360), .A2(n359), .ZN(n358) );
  NAND2_X1 U393 ( .A1(n399), .A2(n357), .ZN(n356) );
  AND2_X1 U394 ( .A1(n373), .A2(n422), .ZN(n357) );
  AND2_X1 U395 ( .A1(n422), .A2(n644), .ZN(n359) );
  XNOR2_X1 U396 ( .A(n461), .B(KEYINPUT75), .ZN(n361) );
  OR2_X1 U397 ( .A1(n390), .A2(n387), .ZN(n557) );
  XNOR2_X1 U398 ( .A(n426), .B(n370), .ZN(n732) );
  AND2_X1 U399 ( .A1(n442), .A2(n441), .ZN(n440) );
  XNOR2_X1 U400 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U401 ( .A(n398), .B(n496), .ZN(n660) );
  XNOR2_X1 U402 ( .A(n355), .B(n398), .ZN(n689) );
  XNOR2_X1 U403 ( .A(n396), .B(n431), .ZN(n355) );
  XNOR2_X1 U404 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n534) );
  XNOR2_X2 U405 ( .A(n768), .B(n488), .ZN(n398) );
  XNOR2_X2 U406 ( .A(n762), .B(KEYINPUT71), .ZN(n396) );
  XNOR2_X2 U407 ( .A(n436), .B(n435), .ZN(n762) );
  INV_X1 U408 ( .A(n399), .ZN(n360) );
  AND2_X1 U409 ( .A1(n361), .A2(n354), .ZN(n616) );
  AND2_X1 U410 ( .A1(n361), .A2(n353), .ZN(n560) );
  XNOR2_X2 U411 ( .A(G101), .B(KEYINPUT88), .ZN(n362) );
  AND2_X2 U412 ( .A1(n363), .A2(n395), .ZN(n676) );
  NAND2_X1 U413 ( .A1(n365), .A2(n363), .ZN(n434) );
  NAND2_X1 U414 ( .A1(n651), .A2(n650), .ZN(n363) );
  BUF_X1 U415 ( .A(n571), .Z(n364) );
  INV_X1 U416 ( .A(KEYINPUT46), .ZN(n400) );
  INV_X1 U417 ( .A(KEYINPUT30), .ZN(n462) );
  NAND2_X1 U418 ( .A1(G902), .A2(G469), .ZN(n415) );
  XNOR2_X1 U419 ( .A(n534), .B(n466), .ZN(n465) );
  XNOR2_X1 U420 ( .A(KEYINPUT70), .B(G137), .ZN(n466) );
  XNOR2_X1 U421 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n536) );
  AND2_X1 U422 ( .A1(n456), .A2(n646), .ZN(n422) );
  NOR2_X1 U423 ( .A1(n430), .A2(n551), .ZN(n429) );
  NOR2_X1 U424 ( .A1(n455), .A2(n453), .ZN(n452) );
  NOR2_X1 U425 ( .A1(n598), .A2(n463), .ZN(n455) );
  NAND2_X1 U426 ( .A1(n430), .A2(KEYINPUT76), .ZN(n454) );
  NAND2_X1 U427 ( .A1(G902), .A2(G472), .ZN(n391) );
  INV_X1 U428 ( .A(KEYINPUT96), .ZN(n554) );
  INV_X1 U429 ( .A(KEYINPUT1), .ZN(n380) );
  INV_X1 U430 ( .A(G113), .ZN(n493) );
  XNOR2_X1 U431 ( .A(KEYINPUT3), .B(G119), .ZN(n494) );
  INV_X1 U432 ( .A(KEYINPUT64), .ZN(n433) );
  XNOR2_X1 U433 ( .A(n526), .B(n525), .ZN(n432) );
  XOR2_X1 U434 ( .A(KEYINPUT93), .B(KEYINPUT77), .Z(n525) );
  INV_X1 U435 ( .A(G146), .ZN(n488) );
  INV_X1 U436 ( .A(KEYINPUT39), .ZN(n444) );
  INV_X1 U437 ( .A(n707), .ZN(n617) );
  NAND2_X1 U438 ( .A1(n427), .A2(n479), .ZN(n426) );
  BUF_X1 U439 ( .A(n557), .Z(n736) );
  XNOR2_X1 U440 ( .A(G107), .B(G104), .ZN(n435) );
  XNOR2_X1 U441 ( .A(n639), .B(n408), .ZN(n407) );
  NOR2_X1 U442 ( .A1(n640), .A2(n369), .ZN(n409) );
  INV_X1 U443 ( .A(KEYINPUT80), .ZN(n408) );
  NAND2_X1 U444 ( .A1(n413), .A2(n479), .ZN(n412) );
  INV_X1 U445 ( .A(G469), .ZN(n413) );
  NAND2_X1 U446 ( .A1(n457), .A2(KEYINPUT48), .ZN(n456) );
  NAND2_X1 U447 ( .A1(n366), .A2(n649), .ZN(n441) );
  NAND2_X1 U448 ( .A1(n389), .A2(n479), .ZN(n388) );
  INV_X1 U449 ( .A(G472), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n423), .B(G146), .ZN(n535) );
  INV_X1 U451 ( .A(G125), .ZN(n423) );
  XNOR2_X1 U452 ( .A(G140), .B(G119), .ZN(n446) );
  XNOR2_X1 U453 ( .A(G137), .B(G128), .ZN(n447) );
  XNOR2_X1 U454 ( .A(KEYINPUT94), .B(KEYINPUT23), .ZN(n449) );
  INV_X1 U455 ( .A(G134), .ZN(n467) );
  INV_X1 U456 ( .A(n544), .ZN(n649) );
  XNOR2_X1 U457 ( .A(G143), .B(G113), .ZN(n497) );
  XOR2_X1 U458 ( .A(G122), .B(G104), .Z(n498) );
  INV_X1 U459 ( .A(n677), .ZN(n427) );
  XOR2_X1 U460 ( .A(G101), .B(G116), .Z(n490) );
  XNOR2_X1 U461 ( .A(n535), .B(KEYINPUT10), .ZN(n506) );
  XNOR2_X1 U462 ( .A(n448), .B(n445), .ZN(n474) );
  XNOR2_X1 U463 ( .A(n450), .B(n449), .ZN(n448) );
  XNOR2_X1 U464 ( .A(n447), .B(n446), .ZN(n445) );
  XNOR2_X1 U465 ( .A(G110), .B(KEYINPUT24), .ZN(n450) );
  XNOR2_X1 U466 ( .A(n419), .B(n543), .ZN(n669) );
  XNOR2_X1 U467 ( .A(n428), .B(KEYINPUT28), .ZN(n625) );
  INV_X1 U468 ( .A(n579), .ZN(n417) );
  INV_X1 U469 ( .A(KEYINPUT105), .ZN(n464) );
  XNOR2_X1 U470 ( .A(n432), .B(n524), .ZN(n431) );
  AND2_X1 U471 ( .A1(n548), .A2(n458), .ZN(n645) );
  INV_X1 U472 ( .A(n710), .ZN(n443) );
  XNOR2_X1 U473 ( .A(n620), .B(n378), .ZN(n421) );
  INV_X1 U474 ( .A(KEYINPUT31), .ZN(n459) );
  INV_X1 U475 ( .A(n741), .ZN(n437) );
  INV_X1 U476 ( .A(KEYINPUT84), .ZN(n574) );
  INV_X1 U477 ( .A(n556), .ZN(n430) );
  AND2_X1 U478 ( .A1(n395), .A2(G475), .ZN(n365) );
  XOR2_X1 U479 ( .A(n547), .B(n546), .Z(n366) );
  XOR2_X1 U480 ( .A(n578), .B(KEYINPUT104), .Z(n367) );
  AND2_X1 U481 ( .A1(n577), .A2(n429), .ZN(n368) );
  NOR2_X1 U482 ( .A1(KEYINPUT47), .A2(n643), .ZN(n369) );
  XOR2_X1 U483 ( .A(n481), .B(KEYINPUT25), .Z(n370) );
  AND2_X1 U484 ( .A1(n556), .A2(n463), .ZN(n371) );
  AND2_X1 U485 ( .A1(n598), .A2(n597), .ZN(n372) );
  OR2_X1 U486 ( .A1(n457), .A2(KEYINPUT48), .ZN(n373) );
  AND2_X1 U487 ( .A1(n588), .A2(n587), .ZN(n374) );
  OR2_X1 U488 ( .A1(n366), .A2(n649), .ZN(n375) );
  XOR2_X1 U489 ( .A(n569), .B(KEYINPUT0), .Z(n376) );
  XOR2_X1 U490 ( .A(n572), .B(KEYINPUT22), .Z(n377) );
  XOR2_X1 U491 ( .A(n619), .B(KEYINPUT112), .Z(n378) );
  XNOR2_X1 U492 ( .A(KEYINPUT59), .B(n684), .ZN(n379) );
  INV_X1 U493 ( .A(G122), .ZN(n515) );
  NAND2_X1 U494 ( .A1(n394), .A2(n415), .ZN(n414) );
  NAND2_X1 U495 ( .A1(n660), .A2(G472), .ZN(n392) );
  NAND2_X1 U496 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U497 ( .A(n555), .B(n554), .ZN(n598) );
  INV_X1 U498 ( .A(n458), .ZN(n381) );
  INV_X1 U499 ( .A(n382), .ZN(n383) );
  NAND2_X1 U500 ( .A1(n624), .A2(n368), .ZN(n428) );
  NAND2_X1 U501 ( .A1(n409), .A2(n407), .ZN(n457) );
  BUF_X1 U502 ( .A(n438), .Z(n384) );
  NAND2_X1 U503 ( .A1(n381), .A2(n720), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n559), .A2(n720), .ZN(n629) );
  BUF_X1 U505 ( .A(n421), .Z(n386) );
  NAND2_X1 U506 ( .A1(n689), .A2(G469), .ZN(n394) );
  XNOR2_X1 U507 ( .A(n396), .B(n763), .ZN(n419) );
  NOR2_X1 U508 ( .A1(n660), .A2(n388), .ZN(n387) );
  XNOR2_X1 U509 ( .A(n558), .B(n462), .ZN(n393) );
  NAND2_X1 U510 ( .A1(n393), .A2(n454), .ZN(n453) );
  INV_X1 U511 ( .A(n395), .ZN(n717) );
  NAND2_X1 U512 ( .A1(n657), .A2(n656), .ZN(n395) );
  AND2_X1 U513 ( .A1(n397), .A2(n374), .ZN(n699) );
  XNOR2_X1 U514 ( .A(n416), .B(n400), .ZN(n399) );
  XNOR2_X1 U515 ( .A(n401), .B(KEYINPUT72), .ZN(n590) );
  NAND2_X1 U516 ( .A1(n403), .A2(n592), .ZN(n401) );
  NAND2_X1 U517 ( .A1(n417), .A2(n367), .ZN(n402) );
  NOR2_X2 U518 ( .A1(n607), .A2(n699), .ZN(n403) );
  XNOR2_X2 U519 ( .A(n586), .B(KEYINPUT35), .ZN(n607) );
  INV_X1 U520 ( .A(n384), .ZN(n719) );
  XNOR2_X2 U521 ( .A(n404), .B(KEYINPUT33), .ZN(n438) );
  NAND2_X1 U522 ( .A1(n406), .A2(n405), .ZN(n404) );
  INV_X1 U523 ( .A(n582), .ZN(n405) );
  XNOR2_X1 U524 ( .A(n596), .B(KEYINPUT106), .ZN(n406) );
  INV_X1 U525 ( .A(n652), .ZN(n715) );
  XNOR2_X1 U526 ( .A(n652), .B(KEYINPUT74), .ZN(n647) );
  NAND2_X1 U527 ( .A1(n410), .A2(KEYINPUT44), .ZN(n609) );
  INV_X1 U528 ( .A(n608), .ZN(n410) );
  XNOR2_X1 U529 ( .A(n608), .B(n515), .ZN(n780) );
  NOR2_X1 U530 ( .A1(n689), .A2(n412), .ZN(n411) );
  AND2_X2 U531 ( .A1(n581), .A2(n729), .ZN(n596) );
  NAND2_X1 U532 ( .A1(n421), .A2(n420), .ZN(n416) );
  XNOR2_X1 U533 ( .A(n418), .B(KEYINPUT85), .ZN(n611) );
  NAND2_X1 U534 ( .A1(n609), .A2(n610), .ZN(n418) );
  INV_X1 U535 ( .A(n781), .ZN(n420) );
  XNOR2_X1 U536 ( .A(n386), .B(G131), .ZN(G33) );
  XNOR2_X1 U537 ( .A(n424), .B(n686), .ZN(G60) );
  NAND2_X1 U538 ( .A1(n425), .A2(n685), .ZN(n424) );
  XNOR2_X1 U539 ( .A(n434), .B(n379), .ZN(n425) );
  XNOR2_X2 U540 ( .A(n433), .B(G953), .ZN(n771) );
  NAND2_X1 U541 ( .A1(n571), .A2(n437), .ZN(n460) );
  NAND2_X1 U542 ( .A1(n364), .A2(n372), .ZN(n695) );
  NAND2_X1 U543 ( .A1(n438), .A2(n364), .ZN(n584) );
  XNOR2_X2 U544 ( .A(n570), .B(n376), .ZN(n571) );
  OR2_X1 U545 ( .A1(n669), .A2(n375), .ZN(n439) );
  NAND2_X1 U546 ( .A1(n669), .A2(n366), .ZN(n442) );
  XNOR2_X2 U547 ( .A(n629), .B(KEYINPUT19), .ZN(n633) );
  AND2_X1 U548 ( .A1(n618), .A2(n443), .ZN(n714) );
  XNOR2_X1 U549 ( .A(n616), .B(n444), .ZN(n618) );
  NAND2_X1 U550 ( .A1(n452), .A2(n451), .ZN(n461) );
  NAND2_X1 U551 ( .A1(n598), .A2(n371), .ZN(n451) );
  INV_X1 U552 ( .A(n559), .ZN(n458) );
  XNOR2_X2 U553 ( .A(n460), .B(n459), .ZN(n709) );
  INV_X1 U554 ( .A(KEYINPUT76), .ZN(n463) );
  XNOR2_X2 U555 ( .A(n468), .B(G143), .ZN(n539) );
  NAND2_X1 U556 ( .A1(n729), .A2(n383), .ZN(n555) );
  OR2_X1 U557 ( .A1(G902), .A2(n680), .ZN(n469) );
  INV_X1 U558 ( .A(G902), .ZN(n479) );
  AND2_X1 U559 ( .A1(n621), .A2(n733), .ZN(n470) );
  INV_X1 U560 ( .A(KEYINPUT48), .ZN(n644) );
  INV_X1 U561 ( .A(KEYINPUT68), .ZN(n552) );
  XNOR2_X1 U562 ( .A(n614), .B(n613), .ZN(n655) );
  INV_X1 U563 ( .A(KEYINPUT82), .ZN(n653) );
  BUF_X1 U564 ( .A(n581), .Z(n730) );
  XOR2_X1 U565 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n472) );
  XNOR2_X1 U566 ( .A(G902), .B(KEYINPUT15), .ZN(n544) );
  NAND2_X1 U567 ( .A1(G234), .A2(n544), .ZN(n471) );
  XNOR2_X1 U568 ( .A(n472), .B(n471), .ZN(n480) );
  AND2_X1 U569 ( .A1(n480), .A2(G221), .ZN(n473) );
  XNOR2_X1 U570 ( .A(n473), .B(KEYINPUT21), .ZN(n733) );
  INV_X1 U571 ( .A(n733), .ZN(n551) );
  INV_X1 U572 ( .A(n506), .ZN(n475) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n478) );
  NAND2_X1 U574 ( .A1(n771), .A2(G234), .ZN(n476) );
  XOR2_X1 U575 ( .A(KEYINPUT8), .B(n476), .Z(n511) );
  NAND2_X1 U576 ( .A1(G221), .A2(n511), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n677) );
  NAND2_X1 U578 ( .A1(G217), .A2(n480), .ZN(n481) );
  INV_X1 U579 ( .A(n732), .ZN(n577) );
  NAND2_X1 U580 ( .A1(G234), .A2(G237), .ZN(n482) );
  XNOR2_X1 U581 ( .A(n482), .B(KEYINPUT14), .ZN(n485) );
  NAND2_X1 U582 ( .A1(G952), .A2(n485), .ZN(n483) );
  XNOR2_X1 U583 ( .A(KEYINPUT90), .B(n483), .ZN(n748) );
  NOR2_X1 U584 ( .A1(n748), .A2(G953), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n484), .B(KEYINPUT91), .ZN(n566) );
  NAND2_X1 U586 ( .A1(G902), .A2(n485), .ZN(n562) );
  NOR2_X1 U587 ( .A1(G900), .A2(n562), .ZN(n486) );
  INV_X1 U588 ( .A(n771), .ZN(n664) );
  NAND2_X1 U589 ( .A1(n486), .A2(n664), .ZN(n487) );
  NAND2_X1 U590 ( .A1(n566), .A2(n487), .ZN(n556) );
  XNOR2_X1 U591 ( .A(KEYINPUT5), .B(G131), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n492) );
  NOR2_X1 U593 ( .A1(G953), .A2(G237), .ZN(n503) );
  NAND2_X1 U594 ( .A1(n503), .A2(G210), .ZN(n491) );
  XNOR2_X1 U595 ( .A(n492), .B(n491), .ZN(n495) );
  XNOR2_X1 U596 ( .A(n494), .B(n493), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n495), .B(n532), .ZN(n496) );
  XNOR2_X1 U598 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n509) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n502) );
  XOR2_X1 U600 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n500) );
  XNOR2_X1 U601 ( .A(KEYINPUT97), .B(KEYINPUT12), .ZN(n499) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U603 ( .A(n502), .B(n501), .Z(n505) );
  NAND2_X1 U604 ( .A1(G214), .A2(n503), .ZN(n504) );
  XNOR2_X1 U605 ( .A(n505), .B(n504), .ZN(n507) );
  XOR2_X1 U606 ( .A(G131), .B(G140), .Z(n526) );
  XOR2_X1 U607 ( .A(n506), .B(n526), .Z(n770) );
  XNOR2_X1 U608 ( .A(n507), .B(n770), .ZN(n684) );
  NOR2_X1 U609 ( .A1(G902), .A2(n684), .ZN(n508) );
  XNOR2_X1 U610 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U611 ( .A(G475), .ZN(n683) );
  XNOR2_X1 U612 ( .A(n510), .B(n683), .ZN(n599) );
  NAND2_X1 U613 ( .A1(n511), .A2(G217), .ZN(n520) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n513) );
  XNOR2_X1 U615 ( .A(G107), .B(KEYINPUT7), .ZN(n512) );
  XNOR2_X1 U616 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U617 ( .A(n514), .B(KEYINPUT101), .Z(n518) );
  XNOR2_X1 U618 ( .A(n515), .B(G116), .ZN(n531) );
  XNOR2_X1 U619 ( .A(n516), .B(n531), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U621 ( .A(n520), .B(n519), .ZN(n680) );
  XNOR2_X1 U622 ( .A(G478), .B(n469), .ZN(n600) );
  INV_X1 U623 ( .A(n600), .ZN(n521) );
  NAND2_X1 U624 ( .A1(n599), .A2(n521), .ZN(n707) );
  NOR2_X1 U625 ( .A1(n582), .A2(n707), .ZN(n522) );
  NAND2_X1 U626 ( .A1(n368), .A2(n522), .ZN(n523) );
  XNOR2_X1 U627 ( .A(KEYINPUT108), .B(n523), .ZN(n630) );
  NAND2_X1 U628 ( .A1(n771), .A2(G227), .ZN(n524) );
  INV_X1 U629 ( .A(n730), .ZN(n587) );
  INV_X1 U630 ( .A(G237), .ZN(n527) );
  NAND2_X1 U631 ( .A1(n479), .A2(n527), .ZN(n545) );
  NAND2_X1 U632 ( .A1(n545), .A2(G214), .ZN(n720) );
  NAND2_X1 U633 ( .A1(n587), .A2(n720), .ZN(n528) );
  NOR2_X1 U634 ( .A1(n630), .A2(n528), .ZN(n530) );
  XNOR2_X1 U635 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n529) );
  XNOR2_X1 U636 ( .A(n530), .B(n529), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n531), .B(KEYINPUT16), .ZN(n533) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n763) );
  XNOR2_X1 U639 ( .A(n535), .B(n534), .ZN(n538) );
  XNOR2_X1 U640 ( .A(n536), .B(KEYINPUT18), .ZN(n537) );
  XNOR2_X1 U641 ( .A(n538), .B(n537), .ZN(n542) );
  NAND2_X1 U642 ( .A1(n771), .A2(G224), .ZN(n540) );
  XNOR2_X1 U643 ( .A(n539), .B(n540), .ZN(n541) );
  XNOR2_X1 U644 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U645 ( .A1(n545), .A2(G210), .ZN(n547) );
  XNOR2_X1 U646 ( .A(KEYINPUT79), .B(KEYINPUT89), .ZN(n546) );
  XOR2_X1 U647 ( .A(G140), .B(KEYINPUT119), .Z(n549) );
  XOR2_X1 U648 ( .A(n645), .B(n549), .Z(G42) );
  NAND2_X1 U649 ( .A1(n599), .A2(n600), .ZN(n550) );
  NAND2_X1 U650 ( .A1(n732), .A2(n733), .ZN(n553) );
  XNOR2_X2 U651 ( .A(n553), .B(n552), .ZN(n729) );
  NAND2_X1 U652 ( .A1(n624), .A2(n720), .ZN(n558) );
  NAND2_X1 U653 ( .A1(n560), .A2(n381), .ZN(n638) );
  XNOR2_X1 U654 ( .A(G143), .B(KEYINPUT118), .ZN(n561) );
  XNOR2_X1 U655 ( .A(n638), .B(n561), .ZN(G45) );
  INV_X1 U656 ( .A(n562), .ZN(n564) );
  INV_X1 U657 ( .A(G898), .ZN(n563) );
  AND2_X1 U658 ( .A1(n563), .A2(G953), .ZN(n764) );
  NAND2_X1 U659 ( .A1(n564), .A2(n764), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U661 ( .A(n567), .B(KEYINPUT92), .ZN(n568) );
  NAND2_X1 U662 ( .A1(n633), .A2(n568), .ZN(n570) );
  INV_X1 U663 ( .A(KEYINPUT67), .ZN(n569) );
  NOR2_X1 U664 ( .A1(n599), .A2(n600), .ZN(n621) );
  NAND2_X1 U665 ( .A1(n571), .A2(n470), .ZN(n573) );
  INV_X1 U666 ( .A(KEYINPUT73), .ZN(n572) );
  XNOR2_X1 U667 ( .A(n579), .B(n574), .ZN(n576) );
  NOR2_X1 U668 ( .A1(n730), .A2(n577), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n576), .A2(n575), .ZN(n605) );
  XNOR2_X1 U670 ( .A(n605), .B(G101), .ZN(G3) );
  NAND2_X1 U671 ( .A1(n730), .A2(n577), .ZN(n578) );
  XNOR2_X1 U672 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n592), .B(G119), .ZN(G21) );
  INV_X1 U674 ( .A(KEYINPUT34), .ZN(n583) );
  XNOR2_X1 U675 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n585), .A2(n353), .ZN(n586) );
  NOR2_X1 U677 ( .A1(n624), .A2(n732), .ZN(n588) );
  INV_X1 U678 ( .A(KEYINPUT44), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n590), .A2(n589), .ZN(n595) );
  NAND2_X1 U680 ( .A1(KEYINPUT72), .A2(KEYINPUT44), .ZN(n591) );
  NOR2_X1 U681 ( .A1(n699), .A2(n591), .ZN(n593) );
  NAND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n596), .A2(n736), .ZN(n741) );
  INV_X1 U685 ( .A(n736), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n709), .A2(n695), .ZN(n602) );
  INV_X1 U687 ( .A(n599), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n601), .A2(n600), .ZN(n710) );
  NAND2_X1 U689 ( .A1(n707), .A2(n710), .ZN(n641) );
  NAND2_X1 U690 ( .A1(n602), .A2(n641), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n603), .B(KEYINPUT102), .ZN(n604) );
  NAND2_X1 U692 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U693 ( .A(n606), .B(KEYINPUT103), .ZN(n610) );
  INV_X1 U694 ( .A(n607), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n614) );
  XOR2_X1 U696 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n613) );
  NAND2_X1 U697 ( .A1(n655), .A2(n649), .ZN(n615) );
  XNOR2_X1 U698 ( .A(n615), .B(KEYINPUT81), .ZN(n648) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U700 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n619) );
  INV_X1 U701 ( .A(n621), .ZN(n722) );
  NAND2_X1 U702 ( .A1(n354), .A2(n720), .ZN(n723) );
  NOR2_X1 U703 ( .A1(n722), .A2(n723), .ZN(n622) );
  XOR2_X1 U704 ( .A(KEYINPUT41), .B(n622), .Z(n623) );
  XNOR2_X1 U705 ( .A(KEYINPUT113), .B(n623), .ZN(n749) );
  INV_X1 U706 ( .A(n383), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT110), .B(n627), .Z(n635) );
  NOR2_X1 U709 ( .A1(n749), .A2(n635), .ZN(n628) );
  XNOR2_X1 U710 ( .A(n628), .B(KEYINPUT42), .ZN(n781) );
  NOR2_X1 U711 ( .A1(n630), .A2(n385), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT36), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n632), .A2(n730), .ZN(n713) );
  INV_X1 U714 ( .A(n633), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n642) );
  INV_X1 U716 ( .A(n642), .ZN(n705) );
  NAND2_X1 U717 ( .A1(n705), .A2(KEYINPUT47), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n713), .A2(n636), .ZN(n640) );
  INV_X1 U719 ( .A(n641), .ZN(n724) );
  NAND2_X1 U720 ( .A1(n724), .A2(KEYINPUT47), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n714), .A2(n645), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n649), .A2(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n652), .A2(KEYINPUT2), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n657) );
  BUF_X1 U728 ( .A(n655), .Z(n656) );
  NAND2_X1 U729 ( .A1(n676), .A2(G472), .ZN(n662) );
  XNOR2_X1 U730 ( .A(KEYINPUT87), .B(KEYINPUT114), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n658), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n662), .B(n661), .ZN(n665) );
  INV_X1 U733 ( .A(G952), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n685) );
  NAND2_X1 U735 ( .A1(n665), .A2(n685), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n676), .A2(G210), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n667), .B(KEYINPUT55), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n672), .A2(n685), .ZN(n675) );
  XNOR2_X1 U743 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n673), .B(KEYINPUT83), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(G51) );
  BUF_X2 U746 ( .A(n676), .Z(n687) );
  NAND2_X1 U747 ( .A1(n687), .A2(G217), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(n679) );
  INV_X1 U749 ( .A(n685), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n679), .A2(n692), .ZN(G66) );
  NAND2_X1 U751 ( .A1(n687), .A2(G478), .ZN(n681) );
  XNOR2_X1 U752 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U753 ( .A1(n682), .A2(n692), .ZN(G63) );
  XNOR2_X1 U754 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n687), .A2(G469), .ZN(n691) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XNOR2_X1 U757 ( .A(n350), .B(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n691), .B(n690), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(G54) );
  NOR2_X1 U760 ( .A1(n707), .A2(n695), .ZN(n694) );
  XOR2_X1 U761 ( .A(G104), .B(n694), .Z(G6) );
  NOR2_X1 U762 ( .A1(n710), .A2(n695), .ZN(n697) );
  XNOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U765 ( .A(G107), .B(n698), .ZN(G9) );
  XNOR2_X1 U766 ( .A(n699), .B(G110), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT115), .ZN(G12) );
  NOR2_X1 U768 ( .A1(n705), .A2(n710), .ZN(n704) );
  XOR2_X1 U769 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n702) );
  XNOR2_X1 U770 ( .A(G128), .B(KEYINPUT117), .ZN(n701) );
  XNOR2_X1 U771 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U772 ( .A(n704), .B(n703), .ZN(G30) );
  NOR2_X1 U773 ( .A1(n705), .A2(n707), .ZN(n706) );
  XOR2_X1 U774 ( .A(G146), .B(n706), .Z(G48) );
  NOR2_X1 U775 ( .A1(n707), .A2(n709), .ZN(n708) );
  XOR2_X1 U776 ( .A(G113), .B(n708), .Z(G15) );
  NOR2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U778 ( .A(G116), .B(n711), .Z(G18) );
  XOR2_X1 U779 ( .A(G125), .B(KEYINPUT37), .Z(n712) );
  XNOR2_X1 U780 ( .A(n713), .B(n712), .ZN(G27) );
  XOR2_X1 U781 ( .A(G134), .B(n714), .Z(G36) );
  INV_X1 U782 ( .A(n656), .ZN(n756) );
  NOR2_X1 U783 ( .A1(n756), .A2(n715), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n716), .A2(KEYINPUT2), .ZN(n718) );
  NOR2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n754) );
  NOR2_X1 U786 ( .A1(n354), .A2(n720), .ZN(n721) );
  NOR2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n726) );
  NOR2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U789 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U790 ( .A(KEYINPUT121), .B(n727), .Z(n728) );
  NOR2_X1 U791 ( .A1(n719), .A2(n728), .ZN(n745) );
  NOR2_X1 U792 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U793 ( .A(KEYINPUT50), .B(n731), .Z(n739) );
  NOR2_X1 U794 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U795 ( .A(KEYINPUT49), .B(n734), .Z(n735) );
  NOR2_X1 U796 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U797 ( .A(KEYINPUT120), .B(n737), .ZN(n738) );
  NAND2_X1 U798 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U799 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U800 ( .A(KEYINPUT51), .B(n742), .ZN(n743) );
  NOR2_X1 U801 ( .A1(n749), .A2(n743), .ZN(n744) );
  NOR2_X1 U802 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U803 ( .A(n746), .B(KEYINPUT52), .ZN(n747) );
  NOR2_X1 U804 ( .A1(n748), .A2(n747), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n749), .A2(n719), .ZN(n750) );
  NOR2_X1 U806 ( .A1(n751), .A2(n750), .ZN(n752) );
  INV_X1 U807 ( .A(G953), .ZN(n774) );
  NAND2_X1 U808 ( .A1(n752), .A2(n774), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U810 ( .A(n755), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U811 ( .A1(n756), .A2(G953), .ZN(n761) );
  NAND2_X1 U812 ( .A1(G953), .A2(G224), .ZN(n757) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n757), .ZN(n758) );
  NAND2_X1 U814 ( .A1(n758), .A2(G898), .ZN(n759) );
  XOR2_X1 U815 ( .A(KEYINPUT124), .B(n759), .Z(n760) );
  NOR2_X1 U816 ( .A1(n761), .A2(n760), .ZN(n767) );
  XNOR2_X1 U817 ( .A(n762), .B(n763), .ZN(n765) );
  NOR2_X1 U818 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U819 ( .A(n767), .B(n766), .Z(G69) );
  XOR2_X1 U820 ( .A(n768), .B(KEYINPUT125), .Z(n769) );
  XOR2_X1 U821 ( .A(n770), .B(n769), .Z(n775) );
  XNOR2_X1 U822 ( .A(n715), .B(n775), .ZN(n772) );
  NAND2_X1 U823 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U824 ( .A(n773), .B(KEYINPUT126), .ZN(n779) );
  XNOR2_X1 U825 ( .A(G227), .B(n775), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U827 ( .A1(G953), .A2(n777), .ZN(n778) );
  NAND2_X1 U828 ( .A1(n779), .A2(n778), .ZN(G72) );
  XNOR2_X1 U829 ( .A(n780), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U830 ( .A(G137), .B(n781), .Z(G39) );
endmodule

