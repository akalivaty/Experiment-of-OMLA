//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1245, new_n1246,
    new_n1247;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n464), .B2(G2105), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT66), .A4(new_n471), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(new_n471), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n482), .A2(KEYINPUT67), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT67), .B1(new_n482), .B2(new_n483), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n480), .A2(new_n484), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n471), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n481), .A2(G126), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT68), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n497), .A3(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n490), .A2(new_n491), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n492), .A2(new_n493), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT69), .A3(G62), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n515), .A2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT70), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(new_n528), .A3(new_n520), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n527), .A2(new_n529), .A3(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n533));
  INV_X1    g108(.A(G63), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n508), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n505), .B(new_n507), .C1(new_n525), .C2(new_n526), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT71), .B(G89), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n536), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n532), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n508), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(new_n538), .B2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n530), .A2(G52), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  AOI22_X1  g131(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n518), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n530), .A2(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n538), .A2(G81), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n508), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n527), .A2(new_n529), .A3(G53), .A4(G543), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g154(.A(KEYINPUT74), .B(new_n573), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  NAND2_X1  g158(.A1(new_n515), .A2(new_n523), .ZN(G303));
  NAND2_X1  g159(.A1(new_n530), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n538), .A2(G87), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n518), .ZN(new_n590));
  NAND2_X1  g165(.A1(G48), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n508), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n590), .B1(new_n521), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT75), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n530), .A2(G47), .B1(G85), .B2(new_n538), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT76), .B1(new_n537), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n521), .A2(new_n512), .A3(new_n603), .A4(G92), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT10), .B1(new_n602), .B2(new_n604), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n527), .A2(new_n529), .A3(G543), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n607), .A2(new_n608), .B1(new_n609), .B2(new_n518), .ZN(new_n610));
  NOR3_X1   g185(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G171), .B2(new_n613), .ZN(G321));
  XNOR2_X1  g190(.A(G321), .B(KEYINPUT77), .ZN(G284));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n581), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n561), .A2(new_n613), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n611), .A2(new_n620), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n622), .B1(new_n625), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n479), .A2(G135), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT80), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2100), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2438), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2438), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n650), .A3(new_n648), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n656), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n643), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n642), .A3(new_n661), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n666), .A3(G14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2084), .B(G2090), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT82), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT83), .Z(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT17), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT84), .Z(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n671), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(new_n670), .C1(new_n673), .C2(new_n675), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT85), .Z(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT86), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n691), .A2(new_n694), .A3(new_n696), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n699), .B(new_n700), .C1(new_n698), .C2(new_n697), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1981), .B(G1986), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(new_n703), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n706), .B1(new_n704), .B2(new_n707), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n689), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n704), .A2(new_n707), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(new_n705), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(new_n708), .A3(new_n688), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  NOR2_X1   g291(.A1(G5), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G171), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT96), .B(G1961), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G28), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(G28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n724), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(G168), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G16), .B2(G21), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT89), .B(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n562), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G1341), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n734), .A2(G19), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n730), .B1(new_n732), .B2(new_n733), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT27), .B(G1996), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G32), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n479), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n481), .A2(G129), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n746), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n742), .B(new_n745), .C1(new_n754), .C2(new_n721), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n751), .B(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n744), .B1(new_n759), .B2(G29), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n760), .A2(KEYINPUT94), .A3(new_n742), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n729), .B(new_n740), .C1(new_n757), .C2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n763));
  INV_X1    g338(.A(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n488), .B2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(new_n767), .B2(new_n763), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT99), .B(G2090), .Z(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n765), .C1(new_n767), .C2(new_n763), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n771), .A2(new_n774), .A3(new_n772), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G34), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(KEYINPUT24), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(KEYINPUT24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n721), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G160), .B2(new_n721), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n760), .A2(new_n742), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n762), .A2(new_n778), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n635), .A2(new_n721), .ZN(new_n788));
  INV_X1    g363(.A(new_n734), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n789), .A2(KEYINPUT23), .A3(G20), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n791));
  INV_X1    g366(.A(G20), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n734), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G16), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n790), .B(new_n793), .C1(new_n581), .C2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1956), .Z(new_n796));
  NAND3_X1  g371(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT25), .Z(new_n798));
  AND2_X1   g373(.A1(new_n461), .A2(new_n463), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n799), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n800));
  INV_X1    g375(.A(G139), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n798), .B1(new_n800), .B2(new_n471), .C1(new_n478), .C2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G33), .B(new_n802), .S(G29), .Z(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G2072), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n721), .A2(G27), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G164), .B2(new_n721), .ZN(new_n806));
  INV_X1    g381(.A(G2078), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n732), .A2(new_n733), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n796), .A2(new_n804), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n787), .A2(new_n788), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n789), .A2(G22), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n789), .ZN(new_n814));
  INV_X1    g389(.A(G1971), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n794), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n794), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT33), .B(G1976), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT90), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n794), .A2(G6), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n594), .B2(new_n794), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT32), .B(G1981), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n816), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT34), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n829), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G290), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n734), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G24), .B2(new_n734), .ZN(new_n838));
  INV_X1    g413(.A(G1986), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n721), .A2(G25), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n481), .A2(G119), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT87), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n479), .A2(G131), .ZN(new_n846));
  OR2_X1    g421(.A1(G95), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT88), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT88), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n842), .B1(new_n853), .B2(G29), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT35), .B(G1991), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n840), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n838), .A2(new_n839), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n812), .B1(new_n835), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g437(.A(KEYINPUT36), .B(new_n860), .C1(new_n832), .C2(new_n834), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n720), .B(new_n811), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT28), .ZN(new_n865));
  INV_X1    g440(.A(G26), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(G29), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(G29), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n479), .A2(G140), .B1(G128), .B2(new_n481), .ZN(new_n869));
  OR2_X1    g444(.A1(G104), .A2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT92), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n868), .B1(new_n873), .B2(G29), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n867), .B1(new_n874), .B2(new_n865), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G2067), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n794), .A2(G4), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n611), .B2(new_n794), .ZN(new_n878));
  INV_X1    g453(.A(G1348), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n864), .A2(new_n876), .A3(new_n881), .ZN(G311));
  INV_X1    g457(.A(new_n787), .ZN(new_n883));
  INV_X1    g458(.A(new_n788), .ZN(new_n884));
  INV_X1    g459(.A(new_n810), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n835), .A2(new_n861), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT36), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n835), .A2(new_n812), .A3(new_n861), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n876), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n880), .A4(new_n720), .ZN(G150));
  AND2_X1   g467(.A1(new_n530), .A2(G55), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n894));
  INV_X1    g469(.A(G93), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n894), .A2(new_n518), .B1(new_n895), .B2(new_n537), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G860), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT37), .Z(new_n900));
  NAND2_X1  g475(.A1(new_n611), .A2(G559), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n897), .A2(KEYINPUT101), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n893), .B2(new_n896), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n562), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n898), .A2(new_n904), .A3(new_n561), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n902), .B(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n900), .B1(new_n911), .B2(G860), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT102), .ZN(G145));
  XNOR2_X1  g488(.A(new_n873), .B(G164), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n802), .B1(new_n752), .B2(new_n753), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n751), .A2(new_n802), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n873), .B(new_n501), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n916), .C1(new_n759), .C2(new_n802), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n481), .A2(G130), .ZN(new_n922));
  NOR2_X1   g497(.A1(G106), .A2(G2105), .ZN(new_n923));
  OAI21_X1  g498(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n924));
  INV_X1    g499(.A(G142), .ZN(new_n925));
  OAI221_X1 g500(.A(new_n922), .B1(new_n923), .B2(new_n924), .C1(new_n478), .C2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(new_n638), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n638), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n853), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n853), .A2(new_n929), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(KEYINPUT103), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n853), .A2(new_n929), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n936), .B2(new_n930), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n921), .A2(new_n933), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n635), .A2(G160), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n635), .A2(G160), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n488), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(G162), .A3(new_n939), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n921), .A2(new_n933), .A3(new_n937), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n933), .A2(new_n937), .ZN(new_n948));
  INV_X1    g523(.A(new_n921), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n934), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n946), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n942), .A2(new_n944), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n931), .A2(new_n932), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n947), .B(new_n952), .C1(new_n953), .C2(new_n921), .ZN(new_n954));
  INV_X1    g529(.A(G37), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT105), .B1(new_n951), .B2(new_n956), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(KEYINPUT40), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT40), .ZN(new_n962));
  INV_X1    g537(.A(new_n956), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n947), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n938), .A3(new_n945), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n958), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n951), .A2(new_n956), .A3(KEYINPUT105), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(G395));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND2_X1  g546(.A1(G166), .A2(G288), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n818), .A2(G303), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n594), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n973), .A3(G305), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n975), .A2(new_n836), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n836), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G290), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n975), .A2(new_n836), .A3(new_n976), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(KEYINPUT108), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n985));
  OR3_X1    g560(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT42), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n579), .A2(new_n580), .A3(new_n611), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n611), .B1(new_n579), .B2(new_n580), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT107), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n581), .A2(new_n612), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT41), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n579), .A2(new_n580), .A3(new_n611), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT41), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n908), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n625), .B(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n625), .B(new_n908), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n996), .B(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n987), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n985), .B(new_n986), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G868), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n897), .A2(G868), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n970), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n613), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1015), .A2(KEYINPUT109), .A3(new_n1012), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(G295));
  NAND2_X1  g592(.A1(new_n1011), .A2(new_n1013), .ZN(G331));
  AND2_X1   g593(.A1(new_n540), .A2(new_n543), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(KEYINPUT110), .A3(new_n531), .A4(new_n536), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n532), .B2(new_n544), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G301), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT110), .B(G168), .C1(new_n553), .C2(new_n554), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n908), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1023), .A2(new_n907), .A3(new_n906), .A4(new_n1024), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n994), .B2(new_n998), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1028), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n996), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1028), .B(new_n1033), .C1(new_n994), .C2(new_n998), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1030), .A2(new_n984), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(new_n955), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1037));
  INV_X1    g612(.A(new_n984), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT43), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n996), .A2(new_n997), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n990), .A2(KEYINPUT41), .A3(new_n993), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1028), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AND4_X1   g620(.A1(KEYINPUT43), .A2(new_n1035), .A3(new_n1045), .A4(new_n955), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT44), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n1049), .A2(new_n1035), .A3(new_n1045), .A4(new_n955), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(G397));
  INV_X1    g628(.A(G1384), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n501), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT112), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n873), .B(G2067), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n751), .A2(G1996), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(new_n1061), .C1(new_n759), .C2(G1996), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n853), .B(new_n855), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(G290), .B(G1986), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1059), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n501), .A2(new_n1054), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT45), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1054), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1057), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n733), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1056), .B1(new_n1067), .B2(KEYINPUT50), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n501), .A2(new_n1074), .A3(new_n1054), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n784), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(KEYINPUT123), .A3(new_n1076), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(G168), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1080), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT123), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G286), .A2(G8), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(G8), .C1(new_n1077), .C2(G286), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1083), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1961), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT124), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1054), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n1096));
  NOR4_X1   g671(.A1(new_n1095), .A2(new_n1055), .A3(new_n1056), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1069), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1067), .A2(KEYINPUT113), .A3(new_n1068), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n807), .A3(new_n1057), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1094), .A2(new_n1103), .A3(KEYINPUT125), .A4(G301), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1093), .B(new_n1097), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(G301), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1094), .A2(G301), .A3(new_n1103), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1092), .B(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G8), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G166), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT55), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1075), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1073), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1074), .B1(new_n501), .B2(new_n1054), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT116), .B1(new_n1117), .B2(new_n1056), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1114), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G2090), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1099), .A2(new_n1057), .A3(new_n1100), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1119), .A2(new_n1120), .B1(new_n1121), .B2(new_n815), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1113), .B1(new_n1122), .B2(new_n1110), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n815), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1073), .A2(new_n1120), .A3(new_n1075), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(G8), .A3(new_n1112), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n818), .A2(G1976), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(G8), .C1(new_n1067), .C2(new_n1056), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT52), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1067), .A2(new_n1056), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1110), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n1133));
  OAI21_X1  g708(.A(G1981), .B1(new_n590), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT49), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT49), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1136), .B(G1981), .C1(new_n590), .C2(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G305), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n594), .A3(new_n1137), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1132), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1976), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT52), .B1(G288), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1132), .A2(new_n1128), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1130), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1123), .A2(new_n1127), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1106), .A2(G301), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT54), .B(new_n1149), .C1(new_n1150), .C2(G301), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1091), .A2(new_n1109), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT56), .B(G2072), .Z(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1119), .A2(G1956), .B1(new_n1121), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n573), .A2(KEYINPUT117), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(new_n577), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1159), .ZN(new_n1161));
  OAI221_X1 g736(.A(new_n1161), .B1(new_n1121), .B2(new_n1154), .C1(new_n1119), .C2(G1956), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT61), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1131), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(G2067), .ZN(new_n1165));
  AOI21_X1  g740(.A(G1348), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT60), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n611), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1168), .A2(new_n611), .A3(new_n1170), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1163), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(G1996), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1099), .A2(new_n1174), .A3(new_n1057), .A4(new_n1100), .ZN(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT58), .B(G1341), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n1164), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1175), .A2(KEYINPUT120), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT120), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n561), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT122), .Z(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1185));
  OR3_X1    g760(.A1(new_n1180), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1155), .A2(KEYINPUT119), .A3(new_n1159), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT119), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1188));
  OAI211_X1 g763(.A(KEYINPUT61), .B(new_n1162), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1184), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1173), .A2(new_n1186), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1187), .A2(new_n1188), .B1(new_n612), .B2(new_n1167), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1162), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1152), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1141), .A2(new_n1142), .A3(new_n818), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1195), .B1(G1981), .B2(G305), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1132), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1145), .B(KEYINPUT115), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1197), .B1(new_n1198), .B2(new_n1127), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1077), .A2(G8), .A3(G168), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1200), .B1(new_n1147), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1126), .A2(G8), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1201), .B1(new_n1203), .B2(new_n1113), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT115), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1145), .B(new_n1205), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1204), .A2(new_n1206), .A3(KEYINPUT63), .A4(new_n1127), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1199), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1106), .A2(G301), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1089), .B1(new_n1081), .B2(G8), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1090), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1209), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1083), .A2(new_n1088), .A3(new_n1214), .A4(new_n1090), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1148), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1208), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1066), .B1(new_n1194), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n1059), .A2(new_n1174), .ZN(new_n1220));
  OR2_X1    g795(.A1(new_n1220), .A2(KEYINPUT46), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1060), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1059), .B1(new_n1222), .B2(new_n751), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1220), .A2(KEYINPUT46), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1221), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  XOR2_X1   g800(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1226));
  XNOR2_X1  g801(.A(new_n1225), .B(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n853), .A2(new_n855), .ZN(new_n1228));
  XOR2_X1   g803(.A(new_n1228), .B(KEYINPUT126), .Z(new_n1229));
  OAI22_X1  g804(.A1(new_n1229), .A2(new_n1062), .B1(G2067), .B2(new_n873), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1064), .A2(new_n1059), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1059), .A2(new_n839), .A3(new_n836), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT48), .ZN(new_n1233));
  AOI22_X1  g808(.A1(new_n1230), .A2(new_n1059), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  AND2_X1   g809(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1219), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g811(.A1(new_n715), .A2(new_n667), .A3(G319), .ZN(new_n1238));
  OAI21_X1  g812(.A(new_n1238), .B1(new_n951), .B2(new_n956), .ZN(new_n1239));
  INV_X1    g813(.A(new_n1039), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n1035), .A2(new_n955), .ZN(new_n1241));
  OAI21_X1  g815(.A(KEYINPUT43), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g816(.A(new_n1051), .ZN(new_n1243));
  AOI211_X1 g817(.A(G227), .B(new_n1239), .C1(new_n1242), .C2(new_n1243), .ZN(G308));
  NAND2_X1  g818(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  INV_X1    g819(.A(G227), .ZN(new_n1246));
  INV_X1    g820(.A(new_n957), .ZN(new_n1247));
  NAND4_X1  g821(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1238), .ZN(G225));
endmodule


