//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  AOI21_X1  g000(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT96), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G64gat), .Z(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT96), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G71gat), .B(G78gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n211), .B(new_n212), .Z(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G211gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n218), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT92), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n225), .A2(G183gat), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(G183gat), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(G231gat), .A2(G233gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n227), .B2(new_n228), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n217), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n231), .A2(new_n232), .A3(new_n217), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n214), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n213), .A3(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT97), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT41), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G43gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G50gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT15), .B1(new_n246), .B2(KEYINPUT88), .ZN(new_n247));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G29gat), .ZN(new_n250));
  INV_X1    g049(.A(G36gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT14), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT14), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G29gat), .B2(G36gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(G29gat), .A2(G36gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT89), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n249), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n256), .A2(KEYINPUT15), .A3(new_n248), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT17), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n267), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270));
  INV_X1    g069(.A(G85gat), .ZN(new_n271));
  INV_X1    g070(.A(G92gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(KEYINPUT8), .A2(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT7), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n271), .B2(new_n272), .ZN(new_n275));
  NAND3_X1  g074(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G99gat), .B(G106gat), .Z(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(KEYINPUT99), .A3(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(KEYINPUT99), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT100), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n244), .B1(new_n269), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G190gat), .B(G218gat), .Z(new_n286));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n283), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT101), .ZN(new_n290));
  XOR2_X1   g089(.A(G134gat), .B(G162gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT98), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n242), .A2(new_n243), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n288), .B2(new_n289), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(KEYINPUT101), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n240), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G230gat), .A2(G233gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT10), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n208), .B1(new_n282), .B2(new_n281), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n279), .A2(new_n280), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n208), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n283), .A2(KEYINPUT10), .A3(new_n208), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT102), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT102), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(new_n308), .B2(new_n309), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n303), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G204gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n305), .A2(new_n307), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n314), .B(new_n320), .C1(new_n303), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n310), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n303), .B(KEYINPUT103), .Z(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n303), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n302), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT87), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G183gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT64), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT65), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT24), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n343), .A2(new_n344), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n341), .A2(new_n345), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n340), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g152(.A(G169gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(new_n316), .ZN(new_n355));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT23), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n340), .A2(new_n349), .A3(new_n362), .A4(new_n351), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n353), .A2(KEYINPUT25), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n345), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n351), .B(new_n365), .C1(G183gat), .C2(G190gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n361), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n355), .A2(KEYINPUT26), .A3(new_n356), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n356), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n336), .A2(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT28), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT28), .B1(new_n376), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n372), .B(new_n373), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT68), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n373), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT28), .ZN(new_n384));
  AND2_X1   g183(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT66), .B(G190gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT28), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT68), .A3(new_n372), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n334), .B1(new_n370), .B2(new_n393), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n383), .B(new_n371), .C1(new_n389), .C2(new_n390), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n333), .B(new_n395), .C1(new_n364), .C2(new_n369), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT73), .B(G218gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n216), .ZN(new_n399));
  OR2_X1    g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(G211gat), .A2(G218gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(KEYINPUT74), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n399), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n394), .A2(new_n396), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n333), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(KEYINPUT29), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n363), .A2(new_n361), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n368), .B1(new_n352), .B2(KEYINPUT67), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n411), .A2(new_n412), .B1(new_n368), .B2(new_n367), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n413), .B2(new_n395), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n370), .A2(new_n393), .A3(new_n409), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n406), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT37), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(G8gat), .B(G36gat), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G64gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G92gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n370), .A2(new_n393), .A3(new_n409), .ZN(new_n423));
  INV_X1    g222(.A(new_n410), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n370), .B2(new_n380), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n407), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n370), .A2(new_n380), .A3(new_n409), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n369), .A2(new_n364), .B1(new_n382), .B2(new_n392), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n406), .C1(new_n429), .C2(new_n334), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT86), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n408), .A2(new_n416), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n427), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n422), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT38), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n331), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n406), .B1(new_n423), .B2(new_n425), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n428), .B(new_n407), .C1(new_n429), .C2(new_n334), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT37), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n420), .B(KEYINPUT76), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n432), .B2(new_n435), .ZN(new_n445));
  AND2_X1   g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G141gat), .B(G148gat), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT2), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(G155gat), .B2(G162gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G141gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G148gat), .ZN(new_n454));
  INV_X1    g253(.A(G148gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G141gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G155gat), .B(G162gat), .ZN(new_n458));
  INV_X1    g257(.A(G155gat), .ZN(new_n459));
  INV_X1    g258(.A(G162gat), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT2), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g263(.A(G134gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G127gat), .ZN(new_n466));
  INV_X1    g265(.A(G127gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G134gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G113gat), .B(G120gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(KEYINPUT1), .ZN(new_n471));
  INV_X1    g270(.A(G120gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G113gat), .ZN(new_n473));
  INV_X1    g272(.A(G113gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G120gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G127gat), .B(G134gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT1), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n481));
  NAND3_X1  g280(.A1(new_n452), .A2(new_n462), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485));
  INV_X1    g284(.A(new_n463), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n471), .A2(new_n479), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n452), .A2(new_n471), .A3(new_n462), .A4(new_n479), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n483), .B(new_n484), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n484), .ZN(new_n492));
  AND4_X1   g291(.A1(new_n462), .A2(new_n452), .A3(new_n471), .A4(new_n479), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n462), .A2(new_n452), .B1(new_n471), .B2(new_n479), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT78), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT78), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n491), .A2(new_n497), .A3(KEYINPUT5), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(new_n485), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT79), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n501), .A2(KEYINPUT79), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n492), .A2(KEYINPUT5), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n483), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT0), .B(G57gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(G85gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G1gat), .B(G29gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n499), .A2(KEYINPUT85), .A3(new_n505), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT85), .B1(new_n499), .B2(new_n505), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n513), .A2(new_n514), .A3(new_n510), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n510), .A3(new_n505), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT80), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n499), .A2(KEYINPUT80), .A3(new_n505), .A4(new_n510), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n512), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n445), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n426), .A2(new_n430), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n420), .B1(new_n524), .B2(KEYINPUT37), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n434), .B1(new_n433), .B2(new_n427), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n431), .A2(KEYINPUT86), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n433), .A2(new_n420), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n438), .A2(new_n523), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n420), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n524), .B2(new_n443), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n524), .A2(new_n421), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n493), .A2(new_n494), .A3(new_n492), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT84), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n502), .A2(new_n503), .A3(new_n483), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n539), .B2(new_n492), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT39), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT39), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n543), .A3(new_n492), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n510), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n515), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n542), .A2(KEYINPUT40), .A3(new_n510), .A4(new_n544), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n536), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G22gat), .B(G50gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G78gat), .B(G106gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT31), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n482), .A2(new_n332), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n406), .A2(KEYINPUT81), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT81), .B1(new_n406), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G228gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n399), .A2(new_n403), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n400), .A2(new_n401), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n332), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n481), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n560), .B1(new_n565), .B2(new_n463), .ZN(new_n566));
  INV_X1    g365(.A(new_n402), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT29), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(KEYINPUT82), .B(new_n463), .C1(new_n570), .C2(KEYINPUT3), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT29), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n572), .B(new_n463), .C1(new_n404), .C2(new_n405), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT82), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n464), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(new_n406), .B2(new_n555), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n406), .A2(new_n576), .A3(new_n555), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n571), .B(new_n575), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI221_X4 g378(.A(new_n554), .B1(new_n558), .B2(new_n566), .C1(new_n579), .C2(new_n560), .ZN(new_n580));
  INV_X1    g379(.A(new_n554), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n571), .A2(new_n575), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n578), .A2(new_n577), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n560), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n558), .A2(new_n566), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n552), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n573), .A2(new_n574), .A3(new_n464), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n574), .B1(new_n573), .B2(new_n464), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n577), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n406), .A2(new_n576), .A3(new_n555), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n559), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n585), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n554), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n584), .A2(new_n581), .A3(new_n585), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n551), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n550), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n531), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT30), .B1(new_n433), .B2(new_n442), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n530), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n506), .A2(new_n511), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n518), .A2(new_n604), .A3(new_n519), .A4(new_n520), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n512), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n606), .A3(new_n532), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n587), .A2(new_n598), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n370), .A2(new_n393), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n480), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n429), .A2(new_n487), .ZN(new_n612));
  INV_X1    g411(.A(G227gat), .ZN(new_n613));
  INV_X1    g412(.A(G233gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT34), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT69), .B(G71gat), .ZN(new_n619));
  INV_X1    g418(.A(G99gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G15gat), .B(G43gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n616), .B1(new_n611), .B2(new_n612), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(KEYINPUT33), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT32), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n612), .ZN(new_n629));
  AOI221_X4 g428(.A(new_n626), .B1(KEYINPUT33), .B2(new_n623), .C1(new_n629), .C2(new_n615), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n618), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT71), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n610), .A2(new_n480), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n429), .A2(new_n487), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n615), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT32), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n638), .A3(new_n623), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT34), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n617), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n627), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n631), .A2(new_n632), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n642), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(KEYINPUT71), .A3(new_n618), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT70), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n631), .A2(new_n650), .A3(new_n643), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(KEYINPUT70), .A3(new_n618), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT36), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n601), .A2(new_n609), .A3(new_n649), .A4(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n536), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT35), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n522), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n647), .A2(new_n655), .A3(new_n599), .A4(new_n657), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n608), .B(new_n607), .C1(new_n651), .C2(new_n652), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT11), .B(G169gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G197gat), .ZN(new_n663));
  XOR2_X1   g462(.A(G113gat), .B(G141gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT90), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n224), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n224), .A2(new_n667), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n267), .B1(new_n262), .B2(new_n264), .ZN(new_n670));
  AOI211_X1 g469(.A(KEYINPUT17), .B(new_n263), .C1(new_n259), .C2(new_n261), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n225), .A2(new_n265), .ZN(new_n673));
  NAND2_X1  g472(.A1(G229gat), .A2(G233gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT91), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT18), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n225), .B(new_n265), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n675), .B(KEYINPUT13), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT93), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n672), .A2(KEYINPUT93), .A3(new_n673), .A4(new_n676), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n678), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n666), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n684), .A2(KEYINPUT94), .A3(new_n678), .A4(new_n685), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n666), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT94), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n687), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n661), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT95), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT95), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n661), .A2(new_n697), .A3(new_n694), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n330), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n606), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT104), .B(G1gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1324gat));
  NAND2_X1  g502(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n704));
  OR2_X1    g503(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n699), .A2(new_n536), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n697), .B1(new_n661), .B2(new_n694), .ZN(new_n709));
  AOI211_X1 g508(.A(KEYINPUT95), .B(new_n693), .C1(new_n654), .C2(new_n660), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n536), .B(new_n329), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G8gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n711), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(KEYINPUT42), .A3(new_n704), .A4(new_n705), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n708), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT105), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n708), .A2(new_n717), .A3(new_n714), .A4(new_n712), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1325gat));
  AOI21_X1  g518(.A(G15gat), .B1(new_n699), .B2(new_n647), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n649), .A2(new_n653), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(G15gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n720), .B1(new_n699), .B2(new_n726), .ZN(G1326gat));
  NAND2_X1  g526(.A1(new_n699), .A2(new_n608), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT107), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n728), .B(new_n730), .ZN(G1327gat));
  INV_X1    g530(.A(new_n328), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n240), .A2(new_n300), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n696), .B2(new_n698), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n250), .A3(new_n700), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT45), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(KEYINPUT45), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n240), .A2(new_n694), .A3(new_n732), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n299), .A2(KEYINPUT44), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT108), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT108), .B1(new_n607), .B2(new_n608), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n601), .A2(new_n742), .A3(new_n649), .A4(new_n653), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n660), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT109), .B1(new_n743), .B2(new_n660), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n739), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n661), .A2(new_n300), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n738), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n749), .A2(new_n700), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n736), .A2(new_n737), .B1(new_n250), .B2(new_n750), .ZN(G1328gat));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n536), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n749), .A2(KEYINPUT110), .A3(new_n536), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(G36gat), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n251), .A3(new_n536), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(G1329gat));
  INV_X1    g559(.A(new_n647), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(G43gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n734), .A2(new_n762), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n721), .B(new_n738), .C1(new_n746), .C2(new_n748), .ZN(new_n764));
  OAI211_X1 g563(.A(KEYINPUT47), .B(new_n763), .C1(new_n764), .C2(new_n245), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n245), .B1(new_n749), .B2(new_n725), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n734), .B2(new_n762), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n769));
  INV_X1    g568(.A(G50gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n749), .B2(new_n608), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n608), .A2(new_n770), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n734), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n749), .A2(new_n777), .A3(new_n608), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G50gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n749), .B2(new_n608), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n781), .B2(new_n769), .ZN(G1331gat));
  OR2_X1    g581(.A1(new_n744), .A2(new_n745), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n302), .A2(new_n732), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n693), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n700), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g587(.A1(new_n785), .A2(new_n655), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  OR3_X1    g592(.A1(new_n785), .A2(G71gat), .A3(new_n761), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795));
  OAI21_X1  g594(.A(G71gat), .B1(new_n785), .B2(new_n724), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(G1334gat));
  NAND2_X1  g598(.A1(new_n786), .A2(new_n608), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g600(.A1(new_n746), .A2(new_n748), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n240), .A2(new_n693), .A3(new_n328), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT113), .Z(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n271), .A3(new_n606), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n743), .A2(new_n660), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n694), .A2(new_n239), .A3(new_n299), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n328), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n700), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n806), .B1(new_n815), .B2(new_n271), .ZN(G1336gat));
  AND2_X1   g615(.A1(new_n802), .A2(new_n804), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n272), .B1(new_n817), .B2(new_n536), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n813), .A2(new_n272), .A3(new_n328), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n655), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G92gat), .B1(new_n805), .B2(new_n655), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n822), .B(new_n823), .C1(new_n655), .C2(new_n819), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(G1337gat));
  NAND3_X1  g624(.A1(new_n814), .A2(new_n620), .A3(new_n647), .ZN(new_n826));
  OAI21_X1  g625(.A(G99gat), .B1(new_n805), .B2(new_n724), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1338gat));
  NAND4_X1  g627(.A1(new_n802), .A2(G106gat), .A3(new_n608), .A4(new_n804), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n810), .A2(new_n608), .A3(new_n328), .A4(new_n812), .ZN(new_n830));
  INV_X1    g629(.A(G106gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n832), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(KEYINPUT115), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n833), .A2(new_n834), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(G1339gat));
  NAND2_X1  g638(.A1(new_n672), .A2(new_n673), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n675), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n842), .B(new_n843), .C1(new_n680), .C2(new_n681), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n665), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n692), .A2(new_n682), .A3(new_n688), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n323), .A2(new_n324), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n314), .A2(KEYINPUT54), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n320), .B1(new_n325), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n851), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n849), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n851), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n854), .A2(new_n857), .A3(new_n322), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n300), .B1(new_n847), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n299), .B1(new_n693), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n847), .A2(new_n732), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n860), .B(new_n240), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n301), .A2(new_n693), .A3(new_n732), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n608), .B1(new_n651), .B2(new_n652), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n536), .A2(new_n606), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n474), .A3(new_n694), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n761), .A2(new_n608), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n868), .ZN(new_n873));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n693), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(G1340gat));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n472), .A3(new_n328), .ZN(new_n876));
  OAI21_X1  g675(.A(G120gat), .B1(new_n873), .B2(new_n732), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1341gat));
  AOI21_X1  g677(.A(G127gat), .B1(new_n869), .B2(new_n239), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n873), .A2(new_n467), .A3(new_n240), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(G1342gat));
  NAND3_X1  g680(.A1(new_n869), .A2(new_n465), .A3(new_n300), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n873), .B2(new_n299), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT58), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n721), .A2(new_n868), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n599), .B1(new_n863), .B2(new_n864), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  AOI211_X1 g691(.A(new_n892), .B(new_n599), .C1(new_n863), .C2(new_n864), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n694), .B(new_n889), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n887), .A2(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n694), .A2(new_n453), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT118), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n724), .A2(new_n890), .A3(new_n868), .A4(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AND4_X1   g699(.A1(new_n888), .A2(new_n895), .A3(new_n896), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n894), .B2(G141gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n888), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(G1344gat));
  OR2_X1    g703(.A1(new_n891), .A2(new_n893), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n889), .B(KEYINPUT120), .Z(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n328), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n890), .A2(new_n724), .A3(new_n868), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n455), .A3(new_n328), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n328), .B(new_n889), .C1(new_n891), .C2(new_n893), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(G148gat), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n908), .B(new_n910), .C1(KEYINPUT59), .C2(new_n912), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n239), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT121), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n905), .A2(new_n889), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n240), .A2(new_n459), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n915), .A2(new_n459), .B1(new_n916), .B2(new_n917), .ZN(G1346gat));
  AOI21_X1  g717(.A(G162gat), .B1(new_n909), .B2(new_n300), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n299), .A2(new_n460), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n916), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n655), .A2(new_n700), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n867), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n354), .A3(new_n694), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n872), .A2(new_n922), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n693), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n316), .A3(new_n328), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  OAI21_X1  g728(.A(G176gat), .B1(new_n925), .B2(new_n732), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  NAND4_X1  g732(.A1(new_n865), .A2(new_n871), .A3(new_n239), .A4(new_n922), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(G183gat), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n923), .A2(new_n377), .A3(new_n239), .ZN(new_n939));
  AND2_X1   g738(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n923), .A2(new_n376), .A3(new_n300), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n872), .A2(new_n300), .A3(new_n922), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(G190gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n945), .B2(G190gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  AND2_X1   g748(.A1(new_n724), .A2(new_n922), .ZN(new_n950));
  XOR2_X1   g749(.A(KEYINPUT125), .B(G197gat), .Z(new_n951));
  NAND4_X1  g750(.A1(new_n950), .A2(new_n694), .A3(new_n890), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT126), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n905), .A2(new_n694), .A3(new_n950), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n955), .B2(new_n951), .ZN(G1352gat));
  NAND3_X1  g755(.A1(new_n905), .A2(new_n328), .A3(new_n950), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n950), .A2(new_n318), .A3(new_n328), .A4(new_n890), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n959), .B2(KEYINPUT62), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n958), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(G1353gat));
  AND2_X1   g763(.A1(new_n950), .A2(new_n890), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n216), .A3(new_n239), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n950), .B(new_n239), .C1(new_n891), .C2(new_n893), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n965), .B2(new_n300), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n905), .A2(new_n950), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n299), .A2(new_n398), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1355gat));
endmodule


