//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n199), .A2(G128), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n200), .B(new_n202), .C1(new_n203), .C2(KEYINPUT23), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(G119), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  AOI22_X1  g021(.A1(new_n204), .A2(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n198), .A2(new_n208), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n204), .A2(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n210), .B(new_n197), .C1(G146), .C2(new_n193), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G137), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XOR2_X1   g029(.A(new_n213), .B(new_n215), .Z(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n209), .A2(new_n211), .A3(new_n216), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G902), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(new_n222), .B(KEYINPUT25), .Z(new_n223));
  XOR2_X1   g037(.A(KEYINPUT74), .B(G217), .Z(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G234), .B2(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(G902), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n199), .B2(G116), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT70), .A3(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n199), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n234), .B2(new_n235), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n232), .A2(KEYINPUT70), .A3(G119), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT70), .B1(new_n232), .B2(G119), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n235), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n240), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n232), .A2(G119), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n231), .B2(new_n233), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n240), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT71), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(new_n255), .B2(G134), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(G137), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(G134), .B2(new_n255), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n258), .A2(KEYINPUT11), .A3(G137), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n263), .B(new_n264), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n262), .A2(new_n268), .A3(KEYINPUT67), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n270), .A3(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n195), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  AOI21_X1  g090(.A(G128), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(KEYINPUT1), .A3(G146), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n273), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G143), .B(G146), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT69), .B(new_n278), .C1(new_n281), .C2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n272), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G131), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n268), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n274), .A2(new_n276), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  OR2_X1    g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n281), .A2(KEYINPUT0), .A3(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(KEYINPUT65), .A3(G131), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n290), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n254), .A2(new_n286), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G237), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G237), .ZN(new_n304));
  AOI21_X1  g118(.A(G953), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n308), .A3(G210), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n307), .B2(new_n309), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n300), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n272), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n271), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n285), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n290), .A2(new_n298), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n296), .B(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT30), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n286), .A2(new_n299), .A3(KEYINPUT30), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n249), .A2(new_n252), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n314), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT31), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n314), .B(new_n328), .C1(new_n322), .C2(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n300), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n278), .B1(new_n281), .B2(G128), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n333), .A2(new_n273), .B1(new_n281), .B2(new_n283), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n272), .A2(new_n315), .B1(new_n282), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n335), .A2(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n336));
  INV_X1    g150(.A(new_n324), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n300), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n332), .B1(new_n338), .B2(KEYINPUT28), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n327), .B(new_n329), .C1(new_n339), .C2(new_n313), .ZN(new_n340));
  NOR2_X1   g154(.A1(G472), .A2(G902), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT32), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n318), .B2(new_n321), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n254), .A2(new_n286), .A3(new_n299), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT28), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n331), .ZN(new_n351));
  INV_X1    g165(.A(new_n253), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n249), .A2(new_n252), .A3(KEYINPUT71), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n286), .A2(new_n299), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT73), .B(KEYINPUT28), .C1(new_n348), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n331), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n353), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n290), .A2(new_n297), .A3(new_n298), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n282), .A2(new_n334), .B1(new_n269), .B2(new_n271), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n330), .B1(new_n361), .B2(new_n300), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n355), .B(KEYINPUT29), .C1(new_n357), .C2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n351), .A2(new_n363), .A3(new_n313), .ZN(new_n364));
  INV_X1    g178(.A(new_n313), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n300), .B(new_n365), .C1(new_n322), .C2(new_n325), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n367), .B2(new_n350), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G472), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n229), .B1(new_n346), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n303), .A2(G237), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n376));
  OAI211_X1 g190(.A(G214), .B(new_n214), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n275), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n263), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n198), .B1(new_n380), .B2(KEYINPUT17), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n377), .A2(new_n275), .ZN(new_n382));
  AOI21_X1  g196(.A(G143), .B1(new_n305), .B2(G214), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT17), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n263), .A3(new_n379), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT18), .A2(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n378), .A2(new_n379), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n193), .B(G146), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT18), .B(G131), .C1(new_n382), .C2(new_n383), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND4_X1   g211(.A1(KEYINPUT86), .A2(new_n388), .A3(new_n391), .A4(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n381), .A2(new_n387), .B1(new_n395), .B2(new_n396), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT86), .B1(new_n399), .B2(new_n391), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n384), .A2(new_n386), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n193), .B(KEYINPUT19), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n402), .B(new_n197), .C1(G146), .C2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n391), .B1(new_n404), .B2(new_n397), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n373), .B(new_n374), .C1(new_n401), .C2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(new_n391), .A3(new_n397), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n399), .A2(KEYINPUT86), .A3(new_n391), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n374), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n399), .A2(new_n391), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n221), .B1(new_n401), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G475), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n201), .A2(G143), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n275), .A2(G128), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT13), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT13), .B1(new_n275), .B2(G128), .ZN(new_n423));
  OAI21_X1  g237(.A(G134), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT88), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n420), .A2(new_n419), .A3(new_n258), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n427));
  INV_X1    g241(.A(G122), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(G116), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n232), .A2(KEYINPUT87), .A3(G122), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n232), .B2(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G107), .ZN(new_n433));
  INV_X1    g247(.A(G107), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n431), .B(new_n434), .C1(new_n232), .C2(G122), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n426), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT89), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(G116), .B2(new_n428), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n434), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n258), .B1(new_n420), .B2(new_n419), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n435), .B1(new_n426), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n437), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT9), .B(G234), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n224), .A2(G953), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n437), .B(new_n447), .C1(new_n442), .C2(new_n444), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n451), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(G234), .A2(G237), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(G952), .A3(new_n214), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n457), .B(KEYINPUT90), .Z(new_n458));
  AND3_X1   g272(.A1(new_n456), .A2(G902), .A3(G953), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n418), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n446), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT77), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n285), .A2(KEYINPUT10), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n434), .A3(G104), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n390), .A2(G107), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n390), .A2(G107), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT75), .B1(new_n472), .B2(new_n468), .ZN(new_n473));
  INV_X1    g287(.A(G101), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n434), .A2(G104), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT75), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n471), .A2(new_n473), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n470), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n466), .B1(new_n467), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(KEYINPUT77), .A3(KEYINPUT10), .A4(new_n285), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n476), .B1(new_n475), .B2(KEYINPUT3), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n469), .A2(new_n470), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n474), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n296), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n471), .A2(new_n477), .A3(new_n473), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G101), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT10), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n283), .A2(new_n274), .A3(new_n276), .A4(KEYINPUT76), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n278), .C1(G128), .C2(new_n281), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT76), .B1(new_n281), .B2(new_n283), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n478), .B(new_n480), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n491), .A2(new_n494), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n290), .A2(new_n298), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n290), .A2(new_n503), .A3(new_n298), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n485), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G140), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n214), .A2(G227), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT12), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT79), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n501), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n499), .B1(new_n483), .B2(new_n285), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n319), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n319), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n492), .A2(new_n490), .A3(G101), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n478), .A2(KEYINPUT4), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n297), .B(new_n522), .C1(new_n523), .C2(new_n489), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n499), .A2(new_n495), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n482), .B2(new_n484), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT80), .B1(new_n527), .B2(new_n501), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n485), .A2(new_n500), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT80), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n319), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n507), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n510), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n521), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n221), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n533), .B1(new_n520), .B2(new_n506), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n528), .A2(new_n531), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n511), .ZN(new_n539));
  OAI21_X1  g353(.A(G469), .B1(new_n539), .B2(G902), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n465), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G214), .B1(G237), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G210), .B1(G237), .B2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n494), .A2(new_n324), .A3(new_n522), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n547));
  OAI21_X1  g361(.A(G113), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n241), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n483), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n546), .A2(new_n553), .A3(new_n551), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(KEYINPUT6), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n297), .A2(new_n191), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT81), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n285), .B2(G125), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n334), .A2(KEYINPUT81), .A3(new_n191), .A4(new_n282), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G224), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n562), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT6), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n552), .A2(new_n567), .A3(new_n554), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n557), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT84), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n550), .A2(new_n481), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n553), .B(KEYINPUT8), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n548), .B(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT82), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n251), .A2(new_n577), .A3(KEYINPUT5), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n481), .B1(new_n579), .B2(new_n252), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n570), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n572), .B1(new_n550), .B2(new_n481), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT83), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n548), .B(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n577), .B1(new_n251), .B2(KEYINPUT5), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n241), .B1(new_n586), .B2(new_n578), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT84), .B(new_n582), .C1(new_n587), .C2(new_n481), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n564), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n562), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(new_n588), .A3(new_n591), .A4(new_n556), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n560), .A2(new_n561), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n558), .B1(new_n593), .B2(KEYINPUT85), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT85), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n560), .A2(new_n595), .A3(new_n561), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n590), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n221), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n545), .B1(new_n569), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(KEYINPUT85), .ZN(new_n600));
  INV_X1    g414(.A(new_n558), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(new_n596), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n589), .B2(new_n564), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n591), .A2(new_n556), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n581), .A2(new_n588), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n557), .A2(new_n566), .A3(new_n568), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(new_n221), .A3(new_n544), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n543), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n463), .A2(new_n541), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n372), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n474), .ZN(G3));
  NAND2_X1  g426(.A1(new_n327), .A2(new_n329), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n313), .B1(new_n349), .B2(new_n331), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n221), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G472), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n342), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n229), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n541), .ZN(new_n619));
  INV_X1    g433(.A(new_n462), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n449), .A2(new_n450), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT91), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n445), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n448), .A2(KEYINPUT92), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n450), .A2(KEYINPUT92), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n445), .A2(new_n624), .A3(new_n626), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n623), .B1(new_n631), .B2(KEYINPUT33), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n452), .A2(G902), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI22_X1  g448(.A1(new_n632), .A2(new_n634), .B1(new_n451), .B2(G478), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n418), .A2(new_n635), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n621), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n619), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND3_X1  g454(.A1(new_n414), .A2(new_n455), .A3(new_n417), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n621), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n618), .A3(new_n541), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n217), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n212), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n227), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n226), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n617), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(new_n463), .A3(new_n541), .A4(new_n609), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  AND3_X1   g468(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n344), .B1(new_n340), .B2(new_n341), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n370), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n541), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n649), .A2(new_n609), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n459), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n458), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n414), .A2(new_n417), .A3(new_n455), .A4(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XOR2_X1   g481(.A(new_n662), .B(KEYINPUT39), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n541), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT40), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n322), .A2(new_n325), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n365), .B1(new_n671), .B2(new_n300), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n361), .A2(new_n300), .A3(new_n365), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n221), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT93), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n346), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n650), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n599), .A2(new_n608), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT38), .Z(new_n680));
  AOI22_X1  g494(.A1(new_n406), .A2(new_n413), .B1(new_n416), .B2(G475), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n451), .B(new_n453), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n542), .ZN(new_n684));
  OR4_X1    g498(.A1(new_n670), .A2(new_n678), .A3(new_n680), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  NAND3_X1  g500(.A1(new_n418), .A2(new_n635), .A3(new_n663), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n659), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n658), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  NOR2_X1   g504(.A1(new_n621), .A2(new_n636), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n520), .A2(new_n506), .A3(new_n533), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n530), .B1(new_n529), .B2(new_n319), .ZN(new_n693));
  AOI211_X1 g507(.A(KEYINPUT80), .B(new_n501), .C1(new_n485), .C2(new_n500), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n506), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n692), .B1(new_n695), .B2(new_n510), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n536), .A3(new_n464), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n697), .A2(new_n536), .A3(KEYINPUT94), .A4(new_n464), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n371), .A2(new_n691), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n371), .A2(new_n642), .A3(new_n700), .A4(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NAND3_X1  g520(.A1(new_n463), .A2(new_n657), .A3(new_n649), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n697), .A2(new_n536), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(KEYINPUT95), .A3(new_n609), .A4(new_n464), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n697), .A2(new_n609), .A3(new_n536), .A4(new_n464), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT95), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n707), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n199), .ZN(G21));
  AND4_X1   g528(.A1(new_n455), .A2(new_n609), .A3(new_n418), .A4(new_n620), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n700), .A2(new_n715), .A3(new_n701), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT97), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n615), .A2(new_n718), .A3(G472), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n229), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n355), .B(new_n365), .C1(new_n357), .C2(new_n362), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n327), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT96), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n327), .A3(KEYINPUT96), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n329), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n341), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n720), .A2(new_n721), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n716), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT98), .B(G122), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G24));
  AOI21_X1  g546(.A(new_n718), .B1(new_n615), .B2(G472), .ZN(new_n733));
  INV_X1    g547(.A(G472), .ZN(new_n734));
  AOI211_X1 g548(.A(KEYINPUT97), .B(new_n734), .C1(new_n340), .C2(new_n221), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n728), .B(new_n649), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT99), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT99), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n720), .A2(new_n738), .A3(new_n649), .A4(new_n728), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n687), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n710), .A2(new_n711), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n710), .A2(new_n711), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT100), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n687), .B1(new_n709), .B2(new_n712), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n737), .A2(new_n739), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT100), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  AND3_X1   g565(.A1(new_n599), .A2(new_n542), .A3(new_n608), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n541), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n687), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT101), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n343), .A2(new_n345), .B1(G472), .B2(new_n369), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n229), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n657), .A2(KEYINPUT101), .A3(new_n721), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT42), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n657), .A2(new_n541), .A3(new_n721), .A4(new_n752), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n687), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  XNOR2_X1  g578(.A(new_n664), .B(KEYINPUT102), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT103), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT102), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n664), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n536), .A2(new_n540), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n769), .A2(new_n464), .A3(new_n752), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT103), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n371), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  OR2_X1    g588(.A1(new_n539), .A2(KEYINPUT45), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n539), .A2(KEYINPUT45), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT104), .ZN(new_n782));
  INV_X1    g596(.A(new_n536), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n779), .B2(new_n780), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n465), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n668), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT105), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n617), .A2(new_n649), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT107), .Z(new_n789));
  NAND2_X1  g603(.A1(new_n635), .A2(new_n681), .ZN(new_n790));
  NAND2_X1  g604(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT44), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n796), .B1(new_n795), .B2(KEYINPUT44), .ZN(new_n798));
  INV_X1    g612(.A(new_n752), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n795), .B2(KEYINPUT44), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n787), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NAND3_X1  g617(.A1(new_n741), .A2(new_n229), .A3(new_n752), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n782), .A2(new_n784), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n805), .B1(new_n806), .B2(new_n465), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n657), .B(new_n804), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n188), .ZN(G42));
  NAND3_X1  g624(.A1(new_n721), .A2(new_n542), .A3(new_n464), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT109), .ZN(new_n812));
  INV_X1    g626(.A(new_n708), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n790), .B(new_n812), .C1(KEYINPUT49), .C2(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT110), .Z(new_n815));
  INV_X1    g629(.A(new_n677), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n680), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n807), .B(new_n808), .C1(new_n464), .C2(new_n813), .ZN(new_n820));
  INV_X1    g634(.A(new_n458), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n794), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n729), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n752), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n822), .A2(new_n698), .A3(new_n799), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n747), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n698), .A2(new_n799), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n816), .A2(new_n827), .A3(new_n721), .A4(new_n821), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n418), .A2(new_n635), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n542), .B1(KEYINPUT115), .B2(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n464), .A2(new_n680), .A3(new_n708), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(KEYINPUT50), .ZN(new_n836));
  AOI211_X1 g650(.A(KEYINPUT115), .B(new_n831), .C1(new_n823), .C2(new_n833), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT116), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n830), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n824), .B1(new_n840), .B2(KEYINPUT117), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n819), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n757), .A2(new_n758), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n825), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT48), .ZN(new_n847));
  OAI211_X1 g661(.A(G952), .B(new_n214), .C1(new_n828), .C2(new_n636), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n709), .A2(new_n712), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n823), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n830), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n836), .A2(new_n837), .A3(new_n819), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n830), .A2(new_n852), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n851), .B1(new_n824), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n843), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n541), .A2(new_n683), .A3(new_n609), .A4(new_n663), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n666), .B(new_n689), .C1(new_n678), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(KEYINPUT52), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n702), .A2(new_n705), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n730), .A3(new_n713), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n759), .A2(new_n762), .B1(new_n766), .B2(new_n772), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n414), .A2(new_n417), .A3(new_n682), .A4(new_n663), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT112), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n681), .A2(KEYINPUT112), .A3(new_n682), .A4(new_n663), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n752), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT113), .A4(new_n752), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n657), .A2(new_n541), .A3(new_n649), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n741), .A2(new_n541), .A3(new_n752), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n737), .B2(new_n739), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n621), .B2(new_n641), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n541), .A3(new_n618), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n621), .A2(new_n887), .A3(new_n641), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n652), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n372), .A2(new_n610), .B1(new_n619), .B2(new_n637), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n872), .A2(new_n873), .A3(new_n886), .A4(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n860), .B1(new_n870), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g710(.A(KEYINPUT53), .B(new_n894), .C1(new_n868), .C2(new_n869), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n859), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT52), .B1(new_n750), .B2(new_n863), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n867), .B(new_n862), .C1(new_n745), .C2(new_n749), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT53), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n870), .A2(new_n860), .A3(new_n895), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(KEYINPUT54), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n898), .A2(new_n904), .A3(KEYINPUT114), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n896), .A2(new_n897), .A3(new_n859), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT54), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n858), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n818), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n214), .A2(G952), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n557), .A2(new_n568), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n566), .ZN(new_n915));
  XOR2_X1   g729(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n896), .A2(new_n897), .A3(new_n221), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n917), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n920), .A4(new_n917), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n913), .B(new_n921), .C1(new_n924), .C2(new_n925), .ZN(G51));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  INV_X1    g741(.A(new_n913), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n898), .A2(new_n904), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n778), .B(KEYINPUT57), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n534), .B(KEYINPUT121), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR4_X1   g747(.A1(new_n896), .A2(new_n897), .A3(new_n221), .A4(new_n777), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n927), .B(new_n928), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n931), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT122), .B1(new_n936), .B2(new_n913), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(G54));
  NAND3_X1  g752(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(new_n411), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n411), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n913), .ZN(G60));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n909), .A2(new_n905), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n946), .A2(KEYINPUT123), .A3(new_n632), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT123), .B1(new_n946), .B2(new_n632), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n632), .A2(new_n944), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n929), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n928), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n902), .A2(new_n903), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n220), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n913), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n902), .A2(new_n647), .A3(new_n903), .A4(new_n954), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(KEYINPUT61), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n957), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n963), .A2(KEYINPUT125), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT125), .B1(new_n963), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n959), .B1(new_n965), .B2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n460), .B2(new_n563), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n872), .A2(new_n893), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n968), .B1(new_n971), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n914), .B1(G898), .B2(new_n214), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G69));
  AOI21_X1  g788(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n809), .B1(new_n787), .B2(new_n801), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n787), .A2(new_n609), .A3(new_n683), .A4(new_n845), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n750), .A2(new_n666), .A3(new_n689), .A4(new_n873), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n214), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n323), .B1(new_n336), .B2(KEYINPUT30), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n403), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n660), .B2(new_n214), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n685), .A2(new_n750), .A3(new_n666), .A4(new_n689), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n799), .B1(new_n636), .B2(new_n641), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(new_n371), .A3(new_n541), .A4(new_n668), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n977), .A2(new_n986), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n990), .A2(new_n214), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n976), .B1(new_n981), .B2(new_n984), .C1(new_n991), .C2(new_n983), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n981), .A2(new_n984), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n983), .B1(new_n990), .B2(new_n214), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n975), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n672), .A2(new_n367), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n902), .A2(new_n903), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n999), .B1(new_n1002), .B2(new_n971), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n366), .B(KEYINPUT127), .Z(new_n1004));
  OAI211_X1 g818(.A(new_n928), .B(new_n1001), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n672), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n990), .A2(new_n970), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n998), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1005), .A2(new_n1008), .ZN(G57));
endmodule


