

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U322 ( .A1(n495), .A2(n557), .ZN(n497) );
  INV_X1 U323 ( .A(KEYINPUT108), .ZN(n496) );
  INV_X1 U324 ( .A(KEYINPUT110), .ZN(n499) );
  XNOR2_X1 U325 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U326 ( .A(n502), .B(n501), .ZN(n510) );
  XNOR2_X1 U327 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U328 ( .A(n343), .B(n342), .ZN(n346) );
  NOR2_X1 U329 ( .A1(n548), .A2(n547), .ZN(n560) );
  XNOR2_X1 U330 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n290) );
  XNOR2_X1 U331 ( .A(n290), .B(KEYINPUT90), .ZN(n291) );
  XOR2_X1 U332 ( .A(n291), .B(KEYINPUT2), .Z(n293) );
  XNOR2_X1 U333 ( .A(G141GAT), .B(G162GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n396) );
  XOR2_X1 U335 ( .A(G85GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U336 ( .A(G29GAT), .B(G1GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U338 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n297) );
  XNOR2_X1 U339 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(n299), .B(n298), .Z(n309) );
  XOR2_X1 U342 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n301) );
  XNOR2_X1 U343 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT78), .Z(n349) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G127GAT), .Z(n303) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n407) );
  XOR2_X1 U349 ( .A(n349), .B(n407), .Z(n305) );
  NAND2_X1 U350 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n396), .B(n310), .ZN(n565) );
  XOR2_X1 U355 ( .A(G1GAT), .B(KEYINPUT70), .Z(n312) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(G22GAT), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n374) );
  XOR2_X1 U358 ( .A(G169GAT), .B(G8GAT), .Z(n420) );
  XOR2_X1 U359 ( .A(n374), .B(n420), .Z(n314) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U362 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n316) );
  XNOR2_X1 U363 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U365 ( .A(n318), .B(n317), .Z(n327) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n319), .B(G29GAT), .ZN(n320) );
  XOR2_X1 U368 ( .A(n320), .B(KEYINPUT8), .Z(n322) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G50GAT), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n363) );
  XOR2_X1 U371 ( .A(KEYINPUT68), .B(G197GAT), .Z(n324) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n363), .B(n325), .ZN(n326) );
  XOR2_X1 U375 ( .A(n327), .B(n326), .Z(n493) );
  XOR2_X1 U376 ( .A(KEYINPUT72), .B(n493), .Z(n549) );
  XOR2_X1 U377 ( .A(KEYINPUT74), .B(G57GAT), .Z(n329) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U380 ( .A(KEYINPUT73), .B(n330), .Z(n382) );
  XOR2_X1 U381 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n332) );
  XNOR2_X1 U382 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n382), .B(n333), .ZN(n348) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  INV_X1 U386 ( .A(G92GAT), .ZN(n334) );
  NAND2_X1 U387 ( .A1(n334), .A2(G64GAT), .ZN(n337) );
  INV_X1 U388 ( .A(G64GAT), .ZN(n335) );
  NAND2_X1 U389 ( .A1(n335), .A2(G92GAT), .ZN(n336) );
  NAND2_X1 U390 ( .A1(n337), .A2(n336), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n428) );
  XOR2_X1 U392 ( .A(G99GAT), .B(G85GAT), .Z(n358) );
  XNOR2_X1 U393 ( .A(n428), .B(n358), .ZN(n343) );
  AND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  INV_X1 U395 ( .A(KEYINPUT31), .ZN(n340) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n344), .B(G148GAT), .ZN(n386) );
  XNOR2_X1 U398 ( .A(n386), .B(KEYINPUT76), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n574) );
  NAND2_X1 U401 ( .A1(n549), .A2(n574), .ZN(n461) );
  XOR2_X1 U402 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n351) );
  XOR2_X1 U403 ( .A(G190GAT), .B(KEYINPUT79), .Z(n419) );
  XNOR2_X1 U404 ( .A(n419), .B(n349), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U406 ( .A(n352), .B(KEYINPUT65), .Z(n357) );
  XOR2_X1 U407 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n354) );
  XNOR2_X1 U408 ( .A(G162GAT), .B(KEYINPUT77), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U410 ( .A(G218GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U412 ( .A(G92GAT), .B(n358), .Z(n360) );
  NAND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U415 ( .A(n362), .B(n361), .Z(n365) );
  XNOR2_X1 U416 ( .A(n363), .B(G106GAT), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n365), .B(n364), .ZN(n559) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G155GAT), .Z(n367) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(G127GAT), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U421 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n369) );
  XNOR2_X1 U422 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U424 ( .A(n371), .B(n370), .Z(n380) );
  XOR2_X1 U425 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n373) );
  XNOR2_X1 U426 ( .A(KEYINPUT83), .B(KEYINPUT80), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U428 ( .A(G183GAT), .B(G211GAT), .Z(n425) );
  XOR2_X1 U429 ( .A(n425), .B(n374), .Z(n376) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n503) );
  NOR2_X1 U435 ( .A1(n559), .A2(n503), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n383), .B(KEYINPUT16), .ZN(n448) );
  XOR2_X1 U437 ( .A(G204GAT), .B(G211GAT), .Z(n389) );
  XOR2_X1 U438 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n385) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U443 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n391) );
  XNOR2_X1 U444 ( .A(G197GAT), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n429) );
  XOR2_X1 U446 ( .A(KEYINPUT88), .B(n429), .Z(n393) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U449 ( .A(n395), .B(n394), .Z(n398) );
  XNOR2_X1 U450 ( .A(G50GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n542) );
  XOR2_X1 U452 ( .A(G176GAT), .B(KEYINPUT84), .Z(n400) );
  XNOR2_X1 U453 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n417) );
  XOR2_X1 U455 ( .A(G71GAT), .B(G134GAT), .Z(n402) );
  XNOR2_X1 U456 ( .A(G169GAT), .B(G43GAT), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U458 ( .A(G99GAT), .B(G190GAT), .Z(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n413) );
  XOR2_X1 U460 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n406) );
  XNOR2_X1 U461 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n421) );
  XNOR2_X1 U463 ( .A(n407), .B(n421), .ZN(n411) );
  XOR2_X1 U464 ( .A(KEYINPUT87), .B(KEYINPUT64), .Z(n409) );
  XNOR2_X1 U465 ( .A(G15GAT), .B(G183GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n415) );
  NAND2_X1 U469 ( .A1(G227GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n547) );
  INV_X1 U472 ( .A(n547), .ZN(n487) );
  NOR2_X1 U473 ( .A1(n542), .A2(n487), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n418), .B(KEYINPUT26), .ZN(n563) );
  XNOR2_X1 U475 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n434) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n433) );
  XOR2_X1 U477 ( .A(n421), .B(KEYINPUT94), .Z(n423) );
  NAND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U480 ( .A(n424), .B(KEYINPUT95), .Z(n427) );
  XNOR2_X1 U481 ( .A(G36GAT), .B(n425), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U483 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n538) );
  XNOR2_X1 U486 ( .A(n434), .B(n538), .ZN(n441) );
  NAND2_X1 U487 ( .A1(n563), .A2(n441), .ZN(n528) );
  XNOR2_X1 U488 ( .A(n528), .B(KEYINPUT97), .ZN(n439) );
  NAND2_X1 U489 ( .A1(n538), .A2(n487), .ZN(n435) );
  NAND2_X1 U490 ( .A1(n435), .A2(n542), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n436), .B(KEYINPUT25), .ZN(n437) );
  XNOR2_X1 U492 ( .A(KEYINPUT98), .B(n437), .ZN(n438) );
  NOR2_X1 U493 ( .A1(n439), .A2(n438), .ZN(n440) );
  NOR2_X1 U494 ( .A1(n440), .A2(n565), .ZN(n446) );
  INV_X1 U495 ( .A(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n542), .B(KEYINPUT67), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n442), .B(KEYINPUT28), .ZN(n489) );
  NOR2_X1 U498 ( .A1(n443), .A2(n489), .ZN(n444) );
  NAND2_X1 U499 ( .A1(n444), .A2(n565), .ZN(n513) );
  NOR2_X1 U500 ( .A1(n487), .A2(n513), .ZN(n445) );
  NOR2_X1 U501 ( .A1(n446), .A2(n445), .ZN(n447) );
  XNOR2_X1 U502 ( .A(KEYINPUT99), .B(n447), .ZN(n459) );
  NAND2_X1 U503 ( .A1(n448), .A2(n459), .ZN(n474) );
  NOR2_X1 U504 ( .A1(n461), .A2(n474), .ZN(n455) );
  NAND2_X1 U505 ( .A1(n565), .A2(n455), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n449), .B(KEYINPUT34), .ZN(n450) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(n450), .ZN(G1324GAT) );
  NAND2_X1 U508 ( .A1(n538), .A2(n455), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n451), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U510 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n453) );
  NAND2_X1 U511 ( .A1(n455), .A2(n487), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U513 ( .A(G15GAT), .B(n454), .ZN(G1326GAT) );
  NAND2_X1 U514 ( .A1(n455), .A2(n489), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U516 ( .A(n559), .B(KEYINPUT101), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT36), .ZN(n582) );
  INV_X1 U518 ( .A(n503), .ZN(n577) );
  NOR2_X1 U519 ( .A1(n582), .A2(n577), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n459), .A2(n458), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT37), .B(n460), .Z(n484) );
  OR2_X1 U522 ( .A1(n461), .A2(n484), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT38), .B(n462), .Z(n471) );
  NAND2_X1 U524 ( .A1(n565), .A2(n471), .ZN(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U527 ( .A(G29GAT), .B(n465), .ZN(G1328GAT) );
  NAND2_X1 U528 ( .A1(n471), .A2(n538), .ZN(n466) );
  XNOR2_X1 U529 ( .A(n466), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U530 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n468) );
  NAND2_X1 U532 ( .A1(n487), .A2(n471), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U535 ( .A(G50GAT), .B(KEYINPUT105), .Z(n473) );
  NAND2_X1 U536 ( .A1(n489), .A2(n471), .ZN(n472) );
  XNOR2_X1 U537 ( .A(n473), .B(n472), .ZN(G1331GAT) );
  XNOR2_X1 U538 ( .A(n574), .B(KEYINPUT41), .ZN(n554) );
  NAND2_X1 U539 ( .A1(n493), .A2(n554), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n483), .A2(n474), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n565), .A2(n480), .ZN(n477) );
  XNOR2_X1 U542 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n475) );
  XNOR2_X1 U543 ( .A(n475), .B(KEYINPUT106), .ZN(n476) );
  XNOR2_X1 U544 ( .A(n477), .B(n476), .ZN(G1332GAT) );
  NAND2_X1 U545 ( .A1(n538), .A2(n480), .ZN(n478) );
  XNOR2_X1 U546 ( .A(n478), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U547 ( .A1(n480), .A2(n487), .ZN(n479) );
  XNOR2_X1 U548 ( .A(n479), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U549 ( .A(G78GAT), .B(KEYINPUT43), .Z(n482) );
  NAND2_X1 U550 ( .A1(n480), .A2(n489), .ZN(n481) );
  XNOR2_X1 U551 ( .A(n482), .B(n481), .ZN(G1335GAT) );
  NOR2_X1 U552 ( .A1(n484), .A2(n483), .ZN(n490) );
  NAND2_X1 U553 ( .A1(n490), .A2(n565), .ZN(n485) );
  XNOR2_X1 U554 ( .A(G85GAT), .B(n485), .ZN(G1336GAT) );
  NAND2_X1 U555 ( .A1(n538), .A2(n490), .ZN(n486) );
  XNOR2_X1 U556 ( .A(n486), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U557 ( .A1(n490), .A2(n487), .ZN(n488) );
  XNOR2_X1 U558 ( .A(n488), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U559 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U560 ( .A(n491), .B(KEYINPUT44), .ZN(n492) );
  XNOR2_X1 U561 ( .A(G106GAT), .B(n492), .ZN(G1339GAT) );
  INV_X1 U562 ( .A(n493), .ZN(n569) );
  NAND2_X1 U563 ( .A1(n569), .A2(n554), .ZN(n494) );
  XOR2_X1 U564 ( .A(n494), .B(KEYINPUT46), .Z(n495) );
  XNOR2_X1 U565 ( .A(KEYINPUT107), .B(n503), .ZN(n557) );
  XNOR2_X1 U566 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X1 U567 ( .A1(n559), .A2(n498), .ZN(n502) );
  XNOR2_X1 U568 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n500) );
  NOR2_X1 U569 ( .A1(n582), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(KEYINPUT45), .B(n504), .ZN(n505) );
  NAND2_X1 U571 ( .A1(n505), .A2(n574), .ZN(n506) );
  XNOR2_X1 U572 ( .A(KEYINPUT111), .B(n506), .ZN(n508) );
  INV_X1 U573 ( .A(n549), .ZN(n507) );
  NAND2_X1 U574 ( .A1(n508), .A2(n507), .ZN(n509) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n539) );
  NOR2_X1 U578 ( .A1(n547), .A2(n513), .ZN(n514) );
  NAND2_X1 U579 ( .A1(n539), .A2(n514), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT113), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n549), .A2(n524), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U583 ( .A(G120GAT), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U584 ( .A1(n524), .A2(n554), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n520) );
  XNOR2_X1 U587 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n524), .A2(n557), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n521), .B(KEYINPUT114), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1342GAT) );
  XOR2_X1 U592 ( .A(G134GAT), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U593 ( .A1(n524), .A2(n559), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1343GAT) );
  XOR2_X1 U595 ( .A(G141GAT), .B(KEYINPUT117), .Z(n530) );
  NAND2_X1 U596 ( .A1(n539), .A2(n565), .ZN(n527) );
  NOR2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n536), .A2(n569), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(G1344GAT) );
  XNOR2_X1 U600 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n532) );
  NAND2_X1 U602 ( .A1(n536), .A2(n554), .ZN(n531) );
  XNOR2_X1 U603 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NAND2_X1 U605 ( .A1(n536), .A2(n577), .ZN(n535) );
  XNOR2_X1 U606 ( .A(n535), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U607 ( .A1(n536), .A2(n559), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n537), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U609 ( .A1(n539), .A2(n538), .ZN(n541) );
  XOR2_X1 U610 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(n567) );
  INV_X1 U612 ( .A(n542), .ZN(n543) );
  OR2_X1 U613 ( .A1(n565), .A2(n543), .ZN(n544) );
  OR2_X1 U614 ( .A1(n567), .A2(n544), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n560), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n550), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n552) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(n553), .Z(n556) );
  NAND2_X1 U623 ( .A1(n560), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT58), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n562), .ZN(G1351GAT) );
  INV_X1 U630 ( .A(n563), .ZN(n564) );
  OR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  OR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT123), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n569), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n578), .ZN(n583) );
  OR2_X1 U641 ( .A1(n583), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

