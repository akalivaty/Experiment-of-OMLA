

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730;

  XNOR2_X1 U370 ( .A(n421), .B(G146), .ZN(n505) );
  XNOR2_X2 U371 ( .A(n354), .B(KEYINPUT0), .ZN(n576) );
  XNOR2_X2 U372 ( .A(n518), .B(KEYINPUT75), .ZN(n626) );
  XNOR2_X2 U373 ( .A(n527), .B(KEYINPUT1), .ZN(n642) );
  XNOR2_X2 U374 ( .A(n478), .B(n477), .ZN(n527) );
  XNOR2_X1 U375 ( .A(n395), .B(n563), .ZN(n582) );
  XNOR2_X1 U376 ( .A(n394), .B(KEYINPUT19), .ZN(n560) );
  INV_X1 U377 ( .A(G125), .ZN(n421) );
  NOR2_X1 U378 ( .A1(n589), .A2(n586), .ZN(n621) );
  NOR2_X1 U379 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U380 ( .A(n358), .B(KEYINPUT41), .ZN(n679) );
  NAND2_X1 U381 ( .A1(n532), .A2(n525), .ZN(n394) );
  OR2_X1 U382 ( .A1(n647), .A2(n646), .ZN(n643) );
  NOR2_X1 U383 ( .A1(n691), .A2(G902), .ZN(n478) );
  XNOR2_X1 U384 ( .A(n400), .B(n501), .ZN(n701) );
  XNOR2_X1 U385 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U386 ( .A(n465), .B(n466), .ZN(n711) );
  NAND2_X1 U387 ( .A1(n470), .A2(n469), .ZN(n472) );
  INV_X1 U388 ( .A(n502), .ZN(n400) );
  XNOR2_X1 U389 ( .A(n505), .B(KEYINPUT10), .ZN(n450) );
  XNOR2_X1 U390 ( .A(n389), .B(n388), .ZN(n500) );
  XNOR2_X1 U391 ( .A(n441), .B(G143), .ZN(n504) );
  XNOR2_X1 U392 ( .A(G137), .B(G140), .ZN(n475) );
  INV_X2 U393 ( .A(G953), .ZN(n716) );
  XNOR2_X1 U394 ( .A(n504), .B(G134), .ZN(n465) );
  AND2_X1 U395 ( .A1(n530), .A2(n371), .ZN(n662) );
  INV_X1 U396 ( .A(n541), .ZN(n371) );
  NAND2_X1 U397 ( .A1(n366), .A2(n401), .ZN(n639) );
  XNOR2_X1 U398 ( .A(n606), .B(n367), .ZN(n366) );
  INV_X1 U399 ( .A(KEYINPUT80), .ZN(n367) );
  XNOR2_X1 U400 ( .A(G113), .B(G131), .ZN(n427) );
  NOR2_X1 U401 ( .A1(n621), .A2(n729), .ZN(n593) );
  XNOR2_X1 U402 ( .A(n462), .B(n422), .ZN(n647) );
  XNOR2_X1 U403 ( .A(n461), .B(KEYINPUT25), .ZN(n422) );
  XNOR2_X1 U404 ( .A(n543), .B(KEYINPUT101), .ZN(n666) );
  OR2_X1 U405 ( .A1(n660), .A2(n661), .ZN(n543) );
  XNOR2_X1 U406 ( .A(n711), .B(n387), .ZN(n386) );
  XOR2_X1 U407 ( .A(KEYINPUT5), .B(G101), .Z(n482) );
  XNOR2_X1 U408 ( .A(n356), .B(n458), .ZN(n698) );
  XNOR2_X1 U409 ( .A(n457), .B(n423), .ZN(n458) );
  XNOR2_X1 U410 ( .A(n713), .B(n453), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n368), .B(n455), .ZN(n457) );
  XNOR2_X1 U412 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n495) );
  XNOR2_X1 U413 ( .A(n496), .B(KEYINPUT18), .ZN(n497) );
  INV_X1 U414 ( .A(G128), .ZN(n441) );
  NAND2_X1 U415 ( .A1(G237), .A2(G234), .ZN(n491) );
  NOR2_X1 U416 ( .A1(n524), .A2(n661), .ZN(n378) );
  INV_X1 U417 ( .A(n530), .ZN(n542) );
  XNOR2_X1 U418 ( .A(n562), .B(KEYINPUT22), .ZN(n563) );
  NAND2_X1 U419 ( .A1(n398), .A2(n396), .ZN(n395) );
  INV_X1 U420 ( .A(n698), .ZN(n405) );
  XNOR2_X1 U421 ( .A(n377), .B(n375), .ZN(n696) );
  XNOR2_X1 U422 ( .A(n444), .B(n376), .ZN(n375) );
  XNOR2_X1 U423 ( .A(n448), .B(n446), .ZN(n377) );
  XNOR2_X1 U424 ( .A(n445), .B(KEYINPUT96), .ZN(n376) );
  XNOR2_X1 U425 ( .A(n411), .B(n410), .ZN(n691) );
  XNOR2_X1 U426 ( .A(n474), .B(n412), .ZN(n411) );
  XNOR2_X1 U427 ( .A(n475), .B(G146), .ZN(n412) );
  AND2_X1 U428 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U429 ( .A1(n683), .A2(n716), .ZN(n382) );
  XNOR2_X1 U430 ( .A(n545), .B(n546), .ZN(n547) );
  XNOR2_X1 U431 ( .A(n626), .B(n365), .ZN(n364) );
  INV_X1 U432 ( .A(KEYINPUT47), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n485), .B(n479), .ZN(n387) );
  XNOR2_X1 U434 ( .A(G146), .B(G137), .ZN(n479) );
  INV_X1 U435 ( .A(G104), .ZN(n468) );
  XNOR2_X1 U436 ( .A(n454), .B(n369), .ZN(n368) );
  INV_X1 U437 ( .A(KEYINPUT88), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n450), .B(n420), .ZN(n713) );
  INV_X1 U439 ( .A(n475), .ZN(n420) );
  XNOR2_X1 U440 ( .A(G128), .B(KEYINPUT24), .ZN(n451) );
  XOR2_X1 U441 ( .A(KEYINPUT89), .B(KEYINPUT67), .Z(n452) );
  XNOR2_X1 U442 ( .A(G140), .B(G143), .ZN(n429) );
  INV_X1 U443 ( .A(KEYINPUT44), .ZN(n360) );
  XNOR2_X1 U444 ( .A(n414), .B(n413), .ZN(n605) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n413) );
  AND2_X1 U446 ( .A1(n647), .A2(n397), .ZN(n514) );
  INV_X1 U447 ( .A(n576), .ZN(n398) );
  AND2_X1 U448 ( .A1(n662), .A2(n397), .ZN(n396) );
  AND2_X2 U449 ( .A1(n605), .A2(n384), .ZN(n715) );
  AND2_X1 U450 ( .A1(n635), .A2(n385), .ZN(n384) );
  INV_X1 U451 ( .A(n728), .ZN(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT16), .B(G122), .ZN(n389) );
  INV_X1 U453 ( .A(KEYINPUT70), .ZN(n388) );
  XNOR2_X1 U454 ( .A(G107), .B(G122), .ZN(n445) );
  XNOR2_X1 U455 ( .A(G116), .B(KEYINPUT95), .ZN(n442) );
  XOR2_X1 U456 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n443) );
  XNOR2_X1 U457 ( .A(n459), .B(KEYINPUT84), .ZN(n600) );
  XNOR2_X1 U458 ( .A(G902), .B(KEYINPUT15), .ZN(n459) );
  XNOR2_X1 U459 ( .A(G131), .B(KEYINPUT4), .ZN(n466) );
  XNOR2_X1 U460 ( .A(n499), .B(n473), .ZN(n474) );
  NOR2_X1 U461 ( .A1(n715), .A2(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U462 ( .A1(n666), .A2(n662), .ZN(n358) );
  AND2_X1 U463 ( .A1(n493), .A2(n515), .ZN(n494) );
  XNOR2_X1 U464 ( .A(n449), .B(G478), .ZN(n530) );
  XNOR2_X1 U465 ( .A(n701), .B(n399), .ZN(n685) );
  XNOR2_X1 U466 ( .A(n503), .B(n506), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n498), .B(n497), .ZN(n503) );
  NOR2_X1 U468 ( .A1(n551), .A2(n520), .ZN(n526) );
  XNOR2_X1 U469 ( .A(n372), .B(KEYINPUT97), .ZN(n725) );
  AND2_X1 U470 ( .A1(n642), .A2(n589), .ZN(n373) );
  INV_X1 U471 ( .A(KEYINPUT120), .ZN(n402) );
  NAND2_X1 U472 ( .A1(n404), .A2(n417), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n404) );
  NAND2_X1 U474 ( .A1(n418), .A2(n417), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n419), .B(n351), .ZN(n418) );
  INV_X1 U476 ( .A(KEYINPUT60), .ZN(n390) );
  NAND2_X1 U477 ( .A1(n392), .A2(n417), .ZN(n391) );
  XNOR2_X1 U478 ( .A(n393), .B(n352), .ZN(n392) );
  XNOR2_X1 U479 ( .A(n689), .B(n361), .ZN(n692) );
  XNOR2_X1 U480 ( .A(n691), .B(n690), .ZN(n361) );
  AND2_X1 U481 ( .A1(n383), .A2(n381), .ZN(n684) );
  NOR2_X1 U482 ( .A1(n678), .A2(n382), .ZN(n381) );
  XNOR2_X1 U483 ( .A(n641), .B(KEYINPUT79), .ZN(n383) );
  INV_X1 U484 ( .A(n547), .ZN(n726) );
  XOR2_X1 U485 ( .A(n508), .B(KEYINPUT86), .Z(n348) );
  XOR2_X1 U486 ( .A(KEYINPUT85), .B(KEYINPUT73), .Z(n349) );
  BUF_X1 U487 ( .A(n647), .Z(n357) );
  INV_X1 U488 ( .A(n357), .ZN(n589) );
  XOR2_X1 U489 ( .A(n578), .B(KEYINPUT74), .Z(n350) );
  XOR2_X1 U490 ( .A(n696), .B(n695), .Z(n351) );
  XOR2_X1 U491 ( .A(n694), .B(n693), .Z(n352) );
  XOR2_X1 U492 ( .A(n549), .B(KEYINPUT81), .Z(n353) );
  NOR2_X1 U493 ( .A1(G952), .A2(n716), .ZN(n699) );
  INV_X1 U494 ( .A(n699), .ZN(n417) );
  INV_X1 U495 ( .A(n577), .ZN(n407) );
  INV_X1 U496 ( .A(n711), .ZN(n410) );
  NOR2_X1 U497 ( .A1(n643), .A2(n642), .ZN(n565) );
  NAND2_X1 U498 ( .A1(n592), .A2(KEYINPUT44), .ZN(n579) );
  XNOR2_X2 U499 ( .A(n355), .B(n350), .ZN(n592) );
  XNOR2_X1 U500 ( .A(n483), .B(n386), .ZN(n609) );
  NOR2_X1 U501 ( .A1(n584), .A2(n522), .ZN(n516) );
  INV_X1 U502 ( .A(n646), .ZN(n397) );
  XNOR2_X1 U503 ( .A(n550), .B(n353), .ZN(n415) );
  NAND2_X1 U504 ( .A1(n560), .A2(n561), .ZN(n354) );
  XNOR2_X2 U505 ( .A(G110), .B(G101), .ZN(n471) );
  NAND2_X1 U506 ( .A1(n408), .A2(n407), .ZN(n355) );
  XNOR2_X2 U507 ( .A(n472), .B(n471), .ZN(n499) );
  NAND2_X1 U508 ( .A1(n359), .A2(n594), .ZN(n595) );
  XNOR2_X1 U509 ( .A(n593), .B(n360), .ZN(n359) );
  XNOR2_X1 U510 ( .A(n362), .B(n613), .ZN(G57) );
  NOR2_X2 U511 ( .A1(n612), .A2(n699), .ZN(n362) );
  NAND2_X1 U512 ( .A1(n363), .A2(n415), .ZN(n414) );
  XNOR2_X1 U513 ( .A(n538), .B(KEYINPUT64), .ZN(n363) );
  NAND2_X1 U514 ( .A1(n364), .A2(n519), .ZN(n529) );
  NAND2_X1 U515 ( .A1(n697), .A2(G210), .ZN(n687) );
  NOR2_X4 U516 ( .A1(n607), .A2(n608), .ZN(n697) );
  XNOR2_X1 U517 ( .A(n370), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U518 ( .A1(n688), .A2(n699), .ZN(n370) );
  NAND2_X1 U519 ( .A1(n374), .A2(n373), .ZN(n372) );
  XNOR2_X1 U520 ( .A(n588), .B(KEYINPUT82), .ZN(n374) );
  NAND2_X1 U521 ( .A1(n379), .A2(n378), .ZN(n551) );
  XNOR2_X1 U522 ( .A(n523), .B(n380), .ZN(n379) );
  INV_X1 U523 ( .A(KEYINPUT99), .ZN(n380) );
  XNOR2_X1 U524 ( .A(n391), .B(n390), .ZN(G60) );
  NAND2_X1 U525 ( .A1(n697), .A2(G475), .ZN(n393) );
  INV_X1 U526 ( .A(n532), .ZN(n520) );
  XNOR2_X2 U527 ( .A(n509), .B(n348), .ZN(n532) );
  NOR2_X2 U528 ( .A1(n582), .A2(n564), .ZN(n588) );
  NAND2_X1 U529 ( .A1(n401), .A2(n715), .ZN(n599) );
  NOR2_X1 U530 ( .A1(n401), .A2(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U531 ( .A1(n401), .A2(n716), .ZN(n706) );
  XNOR2_X2 U532 ( .A(n597), .B(KEYINPUT45), .ZN(n401) );
  XNOR2_X1 U533 ( .A(n403), .B(n402), .ZN(G66) );
  NAND2_X1 U534 ( .A1(n697), .A2(G217), .ZN(n406) );
  XNOR2_X1 U535 ( .A(n409), .B(KEYINPUT34), .ZN(n408) );
  NOR2_X1 U536 ( .A1(n680), .A2(n576), .ZN(n409) );
  XNOR2_X1 U537 ( .A(n416), .B(KEYINPUT119), .ZN(G63) );
  NAND2_X1 U538 ( .A1(n697), .A2(G478), .ZN(n419) );
  XNOR2_X1 U539 ( .A(n687), .B(n686), .ZN(n688) );
  AND2_X1 U540 ( .A1(n544), .A2(n679), .ZN(n545) );
  AND2_X1 U541 ( .A1(n456), .A2(G221), .ZN(n423) );
  XNOR2_X1 U542 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n424) );
  XNOR2_X1 U543 ( .A(KEYINPUT104), .B(KEYINPUT62), .ZN(n425) );
  INV_X1 U544 ( .A(KEYINPUT46), .ZN(n549) );
  INV_X1 U545 ( .A(n730), .ZN(n548) );
  INV_X1 U546 ( .A(KEYINPUT6), .ZN(n521) );
  XNOR2_X1 U547 ( .A(n609), .B(n425), .ZN(n610) );
  XNOR2_X1 U548 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X1 U549 ( .A1(G953), .A2(G237), .ZN(n484) );
  NAND2_X1 U550 ( .A1(G214), .A2(n484), .ZN(n426) );
  XOR2_X1 U551 ( .A(n426), .B(n450), .Z(n438) );
  XOR2_X1 U552 ( .A(G122), .B(G104), .Z(n428) );
  XNOR2_X1 U553 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U554 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n430) );
  XNOR2_X1 U555 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U556 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U557 ( .A(KEYINPUT91), .B(KEYINPUT94), .Z(n434) );
  XNOR2_X1 U558 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n433) );
  XNOR2_X1 U559 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U560 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U561 ( .A(n438), .B(n437), .ZN(n694) );
  NOR2_X1 U562 ( .A1(G902), .A2(n694), .ZN(n440) );
  XNOR2_X1 U563 ( .A(KEYINPUT13), .B(G475), .ZN(n439) );
  XNOR2_X1 U564 ( .A(n440), .B(n439), .ZN(n541) );
  INV_X1 U565 ( .A(n465), .ZN(n446) );
  XNOR2_X1 U566 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U567 ( .A1(G234), .A2(n716), .ZN(n447) );
  XOR2_X1 U568 ( .A(KEYINPUT8), .B(n447), .Z(n456) );
  NAND2_X1 U569 ( .A1(G217), .A2(n456), .ZN(n448) );
  NOR2_X1 U570 ( .A1(n696), .A2(G902), .ZN(n449) );
  NOR2_X1 U571 ( .A1(n541), .A2(n530), .ZN(n630) );
  XNOR2_X1 U572 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U573 ( .A(G119), .B(G110), .Z(n455) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n454) );
  NOR2_X1 U575 ( .A1(n698), .A2(G902), .ZN(n462) );
  NAND2_X1 U576 ( .A1(G234), .A2(n600), .ZN(n460) );
  XNOR2_X1 U577 ( .A(KEYINPUT20), .B(n460), .ZN(n463) );
  AND2_X1 U578 ( .A1(G217), .A2(n463), .ZN(n461) );
  NAND2_X1 U579 ( .A1(n463), .A2(G221), .ZN(n464) );
  XNOR2_X1 U580 ( .A(n464), .B(KEYINPUT21), .ZN(n646) );
  INV_X1 U581 ( .A(G107), .ZN(n467) );
  NAND2_X1 U582 ( .A1(n467), .A2(G104), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n468), .A2(G107), .ZN(n469) );
  NAND2_X1 U584 ( .A1(G227), .A2(n716), .ZN(n473) );
  XNOR2_X1 U585 ( .A(G469), .B(KEYINPUT65), .ZN(n476) );
  XOR2_X1 U586 ( .A(n476), .B(KEYINPUT66), .Z(n477) );
  NOR2_X1 U587 ( .A1(n643), .A2(n527), .ZN(n568) );
  XOR2_X1 U588 ( .A(G113), .B(G116), .Z(n481) );
  XNOR2_X1 U589 ( .A(G119), .B(KEYINPUT3), .ZN(n480) );
  XNOR2_X1 U590 ( .A(n481), .B(n480), .ZN(n502) );
  XNOR2_X1 U591 ( .A(n502), .B(n482), .ZN(n483) );
  AND2_X1 U592 ( .A1(n484), .A2(G210), .ZN(n485) );
  NOR2_X1 U593 ( .A1(n609), .A2(G902), .ZN(n486) );
  XNOR2_X2 U594 ( .A(n486), .B(G472), .ZN(n584) );
  NOR2_X1 U595 ( .A1(G902), .A2(G237), .ZN(n487) );
  XOR2_X1 U596 ( .A(KEYINPUT72), .B(n487), .Z(n507) );
  NAND2_X1 U597 ( .A1(G214), .A2(n507), .ZN(n488) );
  XNOR2_X1 U598 ( .A(n488), .B(KEYINPUT87), .ZN(n661) );
  NOR2_X1 U599 ( .A1(n584), .A2(n661), .ZN(n489) );
  XNOR2_X1 U600 ( .A(KEYINPUT30), .B(n489), .ZN(n493) );
  AND2_X1 U601 ( .A1(n716), .A2(G952), .ZN(n557) );
  NAND2_X1 U602 ( .A1(G953), .A2(G902), .ZN(n555) );
  NOR2_X1 U603 ( .A1(G900), .A2(n555), .ZN(n490) );
  NOR2_X1 U604 ( .A1(n557), .A2(n490), .ZN(n492) );
  XOR2_X1 U605 ( .A(KEYINPUT14), .B(n491), .Z(n675) );
  NOR2_X1 U606 ( .A1(n492), .A2(n675), .ZN(n515) );
  NAND2_X1 U607 ( .A1(n568), .A2(n494), .ZN(n531) );
  XNOR2_X1 U608 ( .A(n349), .B(n495), .ZN(n498) );
  NAND2_X1 U609 ( .A1(G224), .A2(n716), .ZN(n496) );
  XNOR2_X1 U610 ( .A(n504), .B(n505), .ZN(n506) );
  NAND2_X1 U611 ( .A1(n685), .A2(n600), .ZN(n509) );
  NAND2_X1 U612 ( .A1(n507), .A2(G210), .ZN(n508) );
  INV_X1 U613 ( .A(KEYINPUT38), .ZN(n510) );
  XNOR2_X1 U614 ( .A(n520), .B(n510), .ZN(n660) );
  NOR2_X1 U615 ( .A1(n531), .A2(n660), .ZN(n512) );
  INV_X1 U616 ( .A(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n512), .B(n511), .ZN(n539) );
  NAND2_X1 U618 ( .A1(n630), .A2(n539), .ZN(n513) );
  XNOR2_X1 U619 ( .A(KEYINPUT103), .B(n513), .ZN(n728) );
  NAND2_X1 U620 ( .A1(n515), .A2(n514), .ZN(n522) );
  XOR2_X1 U621 ( .A(KEYINPUT28), .B(n516), .Z(n517) );
  NOR2_X1 U622 ( .A1(n527), .A2(n517), .ZN(n544) );
  INV_X1 U623 ( .A(n661), .ZN(n525) );
  NAND2_X1 U624 ( .A1(n544), .A2(n560), .ZN(n518) );
  NAND2_X1 U625 ( .A1(n530), .A2(n541), .ZN(n524) );
  INV_X1 U626 ( .A(n524), .ZN(n628) );
  NOR2_X1 U627 ( .A1(n628), .A2(n630), .ZN(n664) );
  XOR2_X1 U628 ( .A(KEYINPUT77), .B(n664), .Z(n571) );
  NAND2_X1 U629 ( .A1(n626), .A2(n571), .ZN(n519) );
  INV_X1 U630 ( .A(n584), .ZN(n652) );
  XNOR2_X2 U631 ( .A(n652), .B(n521), .ZN(n564) );
  INV_X1 U632 ( .A(n564), .ZN(n573) );
  NOR2_X1 U633 ( .A1(n573), .A2(n522), .ZN(n523) );
  XNOR2_X1 U634 ( .A(KEYINPUT36), .B(n526), .ZN(n528) );
  INV_X1 U635 ( .A(n642), .ZN(n587) );
  NAND2_X1 U636 ( .A1(n528), .A2(n587), .ZN(n634) );
  NAND2_X1 U637 ( .A1(n529), .A2(n634), .ZN(n537) );
  NAND2_X1 U638 ( .A1(n664), .A2(KEYINPUT47), .ZN(n534) );
  NAND2_X1 U639 ( .A1(n542), .A2(n541), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n577), .A2(n531), .ZN(n533) );
  NAND2_X1 U641 ( .A1(n533), .A2(n532), .ZN(n624) );
  NAND2_X1 U642 ( .A1(n534), .A2(n624), .ZN(n535) );
  XNOR2_X1 U643 ( .A(KEYINPUT76), .B(n535), .ZN(n536) );
  NOR2_X1 U644 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U645 ( .A1(n628), .A2(n539), .ZN(n540) );
  XNOR2_X1 U646 ( .A(KEYINPUT40), .B(n540), .ZN(n730) );
  XOR2_X1 U647 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n546) );
  NAND2_X1 U648 ( .A1(n548), .A2(n547), .ZN(n550) );
  XOR2_X1 U649 ( .A(n551), .B(KEYINPUT100), .Z(n552) );
  NAND2_X1 U650 ( .A1(n552), .A2(n642), .ZN(n553) );
  XNOR2_X1 U651 ( .A(KEYINPUT43), .B(n553), .ZN(n554) );
  NAND2_X1 U652 ( .A1(n554), .A2(n520), .ZN(n635) );
  NOR2_X1 U653 ( .A1(G898), .A2(n555), .ZN(n556) );
  OR2_X1 U654 ( .A1(n557), .A2(n556), .ZN(n559) );
  INV_X1 U655 ( .A(n675), .ZN(n558) );
  AND2_X1 U656 ( .A1(n559), .A2(n558), .ZN(n561) );
  XOR2_X1 U657 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n562) );
  INV_X1 U658 ( .A(n576), .ZN(n567) );
  XNOR2_X1 U659 ( .A(n565), .B(KEYINPUT71), .ZN(n574) );
  NOR2_X1 U660 ( .A1(n584), .A2(n574), .ZN(n655) );
  NAND2_X1 U661 ( .A1(n567), .A2(n655), .ZN(n566) );
  XNOR2_X1 U662 ( .A(n566), .B(KEYINPUT31), .ZN(n631) );
  NAND2_X1 U663 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U664 ( .A1(n652), .A2(n569), .ZN(n616) );
  NOR2_X1 U665 ( .A1(n631), .A2(n616), .ZN(n570) );
  NOR2_X1 U666 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U667 ( .A1(n725), .A2(n572), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n575), .B(KEYINPUT33), .ZN(n680) );
  INV_X1 U670 ( .A(KEYINPUT35), .ZN(n578) );
  NAND2_X1 U671 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U672 ( .A(n581), .B(KEYINPUT83), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n583), .B(KEYINPUT98), .ZN(n585) );
  NAND2_X1 U674 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U675 ( .A1(n588), .A2(n587), .ZN(n590) );
  NOR2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U677 ( .A(n591), .B(KEYINPUT32), .ZN(n729) );
  NAND2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U680 ( .A(KEYINPUT2), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n602) );
  INV_X1 U682 ( .A(n600), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n598), .A2(n728), .ZN(n603) );
  AND2_X1 U685 ( .A1(n635), .A2(n603), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U687 ( .A(n639), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n697), .A2(G472), .ZN(n611) );
  XNOR2_X1 U689 ( .A(KEYINPUT63), .B(KEYINPUT105), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n616), .A2(n628), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(KEYINPUT106), .ZN(n615) );
  XNOR2_X1 U692 ( .A(G104), .B(n615), .ZN(G6) );
  XOR2_X1 U693 ( .A(KEYINPUT26), .B(KEYINPUT107), .Z(n618) );
  NAND2_X1 U694 ( .A1(n616), .A2(n630), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n618), .B(n617), .ZN(n620) );
  XOR2_X1 U696 ( .A(G107), .B(KEYINPUT27), .Z(n619) );
  XNOR2_X1 U697 ( .A(n620), .B(n619), .ZN(G9) );
  XOR2_X1 U698 ( .A(G110), .B(n621), .Z(G12) );
  XOR2_X1 U699 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U700 ( .A1(n626), .A2(n630), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n623), .B(n622), .ZN(G30) );
  XNOR2_X1 U702 ( .A(G143), .B(KEYINPUT108), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(n624), .ZN(G45) );
  NAND2_X1 U704 ( .A1(n626), .A2(n628), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n627), .B(G146), .ZN(G48) );
  NAND2_X1 U706 ( .A1(n631), .A2(n628), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n629), .B(G113), .ZN(G15) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(G116), .ZN(G18) );
  XOR2_X1 U710 ( .A(G125), .B(KEYINPUT37), .Z(n633) );
  XNOR2_X1 U711 ( .A(n634), .B(n633), .ZN(G27) );
  XNOR2_X1 U712 ( .A(G140), .B(n635), .ZN(G42) );
  XNOR2_X1 U713 ( .A(n636), .B(KEYINPUT78), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n640) );
  XOR2_X1 U715 ( .A(KEYINPUT50), .B(KEYINPUT109), .Z(n645) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n357), .A2(n646), .ZN(n648) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(n648), .Z(n649) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT110), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U724 ( .A(n656), .B(KEYINPUT51), .Z(n657) );
  XNOR2_X1 U725 ( .A(KEYINPUT111), .B(n657), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n679), .A2(n658), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT112), .B(n659), .Z(n672) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n668) );
  INV_X1 U730 ( .A(n664), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT113), .B(n669), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n680), .A2(n670), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U736 ( .A(n673), .B(KEYINPUT52), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n676), .A2(G952), .ZN(n677) );
  XOR2_X1 U739 ( .A(KEYINPUT114), .B(n677), .Z(n678) );
  INV_X1 U740 ( .A(n679), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U742 ( .A(n682), .B(KEYINPUT115), .ZN(n683) );
  XNOR2_X1 U743 ( .A(n684), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U744 ( .A(n685), .B(n424), .ZN(n686) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n690) );
  NAND2_X1 U746 ( .A1(n697), .A2(G469), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n699), .A2(n692), .ZN(G54) );
  XOR2_X1 U748 ( .A(KEYINPUT116), .B(KEYINPUT59), .Z(n693) );
  XOR2_X1 U749 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n695) );
  NOR2_X1 U750 ( .A1(G898), .A2(n716), .ZN(n700) );
  NOR2_X1 U751 ( .A1(n701), .A2(n700), .ZN(n709) );
  XOR2_X1 U752 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n703) );
  NAND2_X1 U753 ( .A1(G224), .A2(G953), .ZN(n702) );
  XNOR2_X1 U754 ( .A(n703), .B(n702), .ZN(n704) );
  NAND2_X1 U755 ( .A1(G898), .A2(n704), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n705), .B(KEYINPUT122), .ZN(n707) );
  NAND2_X1 U757 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U758 ( .A(n709), .B(n708), .ZN(G69) );
  XOR2_X1 U759 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n710) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U761 ( .A(n713), .B(n712), .ZN(n718) );
  INV_X1 U762 ( .A(n718), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(n716), .ZN(n723) );
  XNOR2_X1 U765 ( .A(G227), .B(n718), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n719), .A2(G900), .ZN(n720) );
  NAND2_X1 U767 ( .A1(G953), .A2(n720), .ZN(n721) );
  XOR2_X1 U768 ( .A(KEYINPUT125), .B(n721), .Z(n722) );
  NAND2_X1 U769 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U770 ( .A(KEYINPUT126), .B(n724), .ZN(G72) );
  XOR2_X1 U771 ( .A(n725), .B(G101), .Z(G3) );
  XNOR2_X1 U772 ( .A(G137), .B(n726), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n727), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U774 ( .A(G134), .B(n728), .Z(G36) );
  XOR2_X1 U775 ( .A(n592), .B(G122), .Z(G24) );
  XOR2_X1 U776 ( .A(G119), .B(n729), .Z(G21) );
  XOR2_X1 U777 ( .A(G131), .B(n730), .Z(G33) );
endmodule

