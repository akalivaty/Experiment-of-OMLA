//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G140), .Z(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT76), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT71), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n195), .A2(G227), .ZN(new_n196));
  XOR2_X1   g010(.A(new_n190), .B(new_n196), .Z(new_n197));
  AND2_X1   g011(.A1(KEYINPUT77), .A2(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT77), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(G107), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT77), .A2(G104), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n202), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT3), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n210), .B2(KEYINPUT3), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n198), .A2(new_n199), .A3(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT78), .B1(new_n217), .B2(new_n201), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT3), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT79), .A3(new_n205), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(G101), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n223), .B(new_n205), .C1(new_n212), .C2(new_n213), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT4), .A4(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT65), .B1(new_n232), .B2(G143), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n230), .A3(G146), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G128), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n232), .A2(G143), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(KEYINPUT0), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n231), .A2(new_n239), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(new_n238), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(KEYINPUT0), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT79), .B1(new_n220), .B2(new_n205), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n215), .B(new_n204), .C1(new_n218), .C2(new_n219), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT81), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .A4(G101), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n216), .A2(new_n221), .A3(new_n249), .A4(G101), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT81), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n229), .A2(new_n244), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n202), .A2(G104), .ZN(new_n255));
  OAI21_X1  g069(.A(G101), .B1(new_n217), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n224), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT82), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n261), .A2(new_n263), .A3(new_n230), .A4(G146), .ZN(new_n264));
  INV_X1    g078(.A(new_n240), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n233), .A2(new_n235), .ZN(new_n266));
  INV_X1    g080(.A(new_n231), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n263), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n266), .A2(G128), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n236), .A2(new_n271), .A3(G128), .A4(new_n268), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n265), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n259), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT10), .ZN(new_n275));
  INV_X1    g089(.A(new_n257), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n272), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n238), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n236), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT10), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n254), .A2(new_n275), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G137), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(KEYINPUT11), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(KEYINPUT11), .ZN(new_n287));
  INV_X1    g101(.A(G137), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n286), .B(new_n287), .C1(G134), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n289), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n283), .A2(KEYINPUT85), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n292), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n254), .A2(new_n275), .A3(new_n298), .A4(new_n282), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n197), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n299), .A2(new_n197), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n277), .A2(new_n240), .A3(new_n264), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n276), .A2(new_n302), .A3(KEYINPUT83), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n280), .A2(KEYINPUT83), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n276), .A2(new_n302), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n303), .B(new_n292), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT12), .B1(new_n292), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n306), .B(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n187), .B(new_n188), .C1(new_n300), .C2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n197), .B1(new_n309), .B2(new_n299), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n297), .B2(new_n301), .ZN(new_n313));
  OAI21_X1  g127(.A(G469), .B1(new_n313), .B2(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G221), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT9), .B(G234), .Z(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n188), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(new_n322), .A3(KEYINPUT72), .A4(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n324), .B(new_n326), .C1(new_n325), .C2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(G146), .ZN(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n195), .A2(G214), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(G143), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n290), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n290), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n331), .B(new_n336), .C1(new_n337), .C2(KEYINPUT17), .ZN(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(new_n207), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(KEYINPUT18), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT18), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n334), .B1(new_n342), .B2(new_n290), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n329), .A2(G146), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT73), .ZN(new_n345));
  INV_X1    g159(.A(new_n329), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n232), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n340), .A3(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n330), .A2(new_n232), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n329), .B(KEYINPUT19), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(G146), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT92), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n337), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(new_n348), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n349), .B1(new_n357), .B2(new_n340), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n359));
  INV_X1    g173(.A(G475), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n188), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n338), .A2(new_n348), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(new_n340), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n349), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n188), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G475), .ZN(new_n368));
  INV_X1    g182(.A(new_n349), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n340), .B1(new_n356), .B2(new_n348), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n360), .B(new_n188), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT93), .B1(new_n371), .B2(KEYINPUT20), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n361), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G234), .ZN(new_n376));
  OAI211_X1 g190(.A(G952), .B(new_n191), .C1(new_n376), .C2(new_n332), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT96), .ZN(new_n378));
  INV_X1    g192(.A(new_n195), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G902), .C1(new_n376), .C2(new_n332), .ZN(new_n380));
  XOR2_X1   g194(.A(KEYINPUT21), .B(G898), .Z(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G122), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT14), .B1(new_n383), .B2(G116), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n384), .A2(new_n385), .B1(G116), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n385), .B2(new_n384), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n383), .A2(KEYINPUT14), .A3(G116), .ZN(new_n388));
  OAI21_X1  g202(.A(G107), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G116), .B(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n202), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n238), .A2(G143), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n230), .A2(G128), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n284), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n389), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n393), .B1(KEYINPUT13), .B2(new_n392), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(KEYINPUT13), .B2(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G134), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n390), .B(new_n202), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n284), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n317), .A2(G217), .A3(new_n191), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT95), .A3(new_n188), .ZN(new_n406));
  INV_X1    g220(.A(G478), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n406), .B(new_n408), .Z(new_n409));
  NAND3_X1  g223(.A1(new_n375), .A2(new_n382), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n320), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n412));
  INV_X1    g226(.A(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G116), .ZN(new_n414));
  INV_X1    g228(.A(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G119), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT2), .B(G113), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n417), .B(KEYINPUT69), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n418), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n250), .B2(new_n252), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n229), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n419), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G113), .B1(new_n414), .B2(KEYINPUT5), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n259), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(G110), .B(G122), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n429), .B1(new_n229), .B2(new_n422), .ZN(new_n435));
  INV_X1    g249(.A(new_n432), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  MUX2_X1   g252(.A(new_n244), .B(new_n302), .S(new_n327), .Z(new_n439));
  NAND2_X1  g253(.A1(new_n191), .A2(G224), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n436), .B1(new_n423), .B2(new_n430), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  NOR4_X1   g258(.A1(new_n435), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n436), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n438), .B(new_n441), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n431), .A2(new_n434), .A3(new_n432), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT86), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n443), .A2(new_n442), .A3(new_n434), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n441), .A4(new_n438), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n439), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n440), .A2(KEYINPUT7), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT89), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n439), .A2(new_n458), .A3(KEYINPUT7), .A4(new_n440), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n417), .A2(new_n425), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT88), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n424), .B1(new_n461), .B2(new_n427), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n276), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n432), .B(KEYINPUT8), .Z(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(new_n464), .C1(new_n428), .C2(new_n276), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n457), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n435), .A2(new_n436), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n455), .A2(new_n456), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n188), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(KEYINPUT90), .A3(new_n188), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n454), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n454), .A2(new_n476), .A3(new_n474), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n412), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI221_X4 g296(.A(new_n477), .B1(new_n473), .B2(new_n472), .C1(new_n447), .C2(new_n453), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n476), .B1(new_n454), .B2(new_n474), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n412), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n411), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT97), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n490));
  XNOR2_X1  g304(.A(G119), .B(G128), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT24), .B(G110), .Z(new_n492));
  AOI21_X1  g306(.A(new_n331), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n413), .A2(G128), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n496), .C1(G119), .C2(new_n238), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G110), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  OAI22_X1  g313(.A1(new_n497), .A2(G110), .B1(new_n491), .B2(new_n492), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n350), .A3(new_n345), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT22), .Z(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n288), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n502), .B(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n490), .B1(new_n507), .B2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n502), .B(new_n505), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G217), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(G234), .B2(new_n188), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(KEYINPUT74), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n509), .B(KEYINPUT75), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n519), .A2(G902), .A3(new_n513), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n195), .A2(G210), .A3(new_n332), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT27), .Z(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT26), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(new_n223), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n288), .A2(G134), .ZN(new_n526));
  OAI21_X1  g340(.A(G131), .B1(new_n526), .B2(new_n285), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n289), .A2(G131), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n302), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n292), .A2(new_n244), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT64), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT30), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT64), .B(new_n534), .C1(new_n529), .C2(new_n530), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n529), .A2(new_n421), .A3(new_n530), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n536), .A2(new_n421), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n421), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT70), .B(new_n540), .C1(new_n533), .C2(new_n535), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n525), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n421), .B1(new_n529), .B2(new_n530), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n531), .B2(new_n540), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n525), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n188), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(G472), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n527), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n273), .B2(new_n264), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n554), .A2(new_n528), .B1(new_n292), .B2(new_n244), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n534), .B1(new_n555), .B2(KEYINPUT64), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT30), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n421), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n538), .A2(new_n537), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n541), .B(new_n525), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n544), .A2(new_n546), .ZN(new_n561));
  INV_X1    g375(.A(new_n525), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT31), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n539), .A2(KEYINPUT31), .A3(new_n525), .A4(new_n541), .ZN(new_n565));
  INV_X1    g379(.A(G472), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n188), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n560), .B2(new_n563), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n570), .A2(KEYINPUT32), .A3(new_n566), .A4(new_n565), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n552), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n521), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT97), .B(new_n411), .C1(new_n482), .C2(new_n486), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n489), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT98), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G3));
  INV_X1    g392(.A(new_n481), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n478), .B2(new_n479), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n382), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n570), .A2(new_n565), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n567), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n521), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n320), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n405), .B(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(G478), .A3(new_n188), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n405), .A2(new_n188), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n407), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n374), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n582), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT99), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT34), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n207), .ZN(G6));
  AND2_X1   g413(.A1(new_n371), .A2(KEYINPUT20), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n361), .B1(new_n600), .B2(KEYINPUT100), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n371), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n602), .B1(G475), .B2(new_n367), .ZN(new_n603));
  INV_X1    g417(.A(new_n409), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n582), .A2(new_n588), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  OR2_X1    g422(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n502), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(G902), .A3(new_n513), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n518), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n586), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT101), .Z(new_n615));
  NAND3_X1  g429(.A1(new_n489), .A2(new_n575), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT37), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G110), .ZN(G12));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n572), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n318), .B1(new_n311), .B2(new_n314), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n378), .B1(new_n380), .B2(G900), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n603), .A2(new_n604), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n580), .A2(new_n620), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  XNOR2_X1  g440(.A(new_n622), .B(KEYINPUT103), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT39), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT40), .Z(new_n630));
  AOI21_X1  g444(.A(new_n562), .B1(new_n539), .B2(new_n541), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n538), .A2(new_n543), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n188), .B1(new_n633), .B2(new_n525), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n569), .A2(new_n571), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT102), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n569), .A2(new_n638), .A3(new_n571), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n375), .A2(new_n409), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n640), .A2(new_n481), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n480), .B(KEYINPUT38), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n630), .A2(new_n612), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT104), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT104), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n230), .ZN(G45));
  INV_X1    g462(.A(new_n622), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n594), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n580), .A2(new_n620), .A3(new_n621), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G146), .ZN(G48));
  AND3_X1   g466(.A1(new_n283), .A2(KEYINPUT85), .A3(new_n292), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT85), .B1(new_n283), .B2(new_n292), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n299), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n197), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n655), .A2(new_n656), .B1(new_n301), .B2(new_n309), .ZN(new_n657));
  OAI21_X1  g471(.A(G469), .B1(new_n657), .B2(G902), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n311), .A3(new_n319), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n573), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(new_n580), .A3(new_n382), .A4(new_n595), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT105), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT41), .B(G113), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  NAND4_X1  g478(.A1(new_n660), .A2(new_n580), .A3(new_n382), .A4(new_n605), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  OAI21_X1  g480(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT106), .B1(new_n667), .B2(new_n659), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n658), .A2(new_n319), .A3(new_n311), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n480), .A2(new_n669), .A3(new_n670), .A4(new_n481), .ZN(new_n671));
  AOI211_X1 g485(.A(new_n410), .B(new_n619), .C1(new_n668), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n413), .ZN(G21));
  NOR2_X1   g487(.A1(new_n659), .A2(new_n587), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n580), .A3(new_n382), .A4(new_n641), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  INV_X1    g490(.A(new_n650), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n614), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n668), .B2(new_n671), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n327), .ZN(G27));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT107), .B1(new_n567), .B2(new_n568), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n571), .A2(KEYINPUT108), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n571), .A2(KEYINPUT108), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OR3_X1    g500(.A1(new_n567), .A2(KEYINPUT108), .A3(new_n568), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n569), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n571), .A2(KEYINPUT108), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n686), .A2(new_n691), .A3(new_n552), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n521), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n621), .A2(new_n481), .A3(new_n478), .A4(new_n479), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n682), .B1(new_n695), .B2(new_n650), .ZN(new_n696));
  NOR4_X1   g510(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n573), .A4(new_n677), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G131), .ZN(G33));
  NOR3_X1   g513(.A1(new_n483), .A2(new_n484), .A3(new_n579), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n623), .A2(KEYINPUT109), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n574), .A3(new_n621), .A4(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n623), .A2(KEYINPUT109), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT110), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G134), .ZN(G36));
  XOR2_X1   g520(.A(new_n313), .B(KEYINPUT45), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND2_X1  g522(.A1(G469), .A2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(KEYINPUT46), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n711), .B(G469), .C1(new_n707), .C2(G902), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n311), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n319), .A3(new_n628), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT111), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n478), .A2(new_n481), .A3(new_n479), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n375), .A2(new_n593), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n717), .B1(KEYINPUT112), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n585), .A3(new_n613), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n716), .B1(new_n723), .B2(KEYINPUT44), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n713), .A2(new_n725), .A3(new_n319), .A4(new_n628), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n723), .A2(KEYINPUT44), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n715), .A2(new_n724), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G137), .ZN(G39));
  NAND2_X1  g543(.A1(new_n713), .A2(new_n319), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT47), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n716), .A2(new_n521), .A3(new_n572), .A4(new_n677), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT113), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(KEYINPUT47), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT114), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n322), .ZN(G42));
  OAI21_X1  g551(.A(new_n594), .B1(new_n409), .B2(new_n374), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n382), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n320), .A2(new_n587), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n482), .B2(new_n486), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n661), .A3(new_n665), .A4(new_n675), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n672), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n576), .A3(new_n616), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n668), .A2(new_n671), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n678), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n625), .A2(new_n651), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n481), .B(new_n641), .C1(new_n483), .C2(new_n484), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n621), .A2(new_n640), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n612), .A2(new_n622), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n625), .A2(new_n651), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n680), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT116), .A3(new_n752), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n650), .A2(new_n586), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n572), .A2(new_n409), .A3(new_n603), .A4(new_n622), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n612), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n700), .A3(new_n621), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n702), .B2(new_n703), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n696), .A2(new_n765), .A3(new_n697), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n753), .A2(KEYINPUT52), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n744), .A2(new_n760), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT53), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n576), .A2(new_n743), .A3(new_n616), .A4(new_n766), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT116), .B1(new_n758), .B2(new_n752), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n680), .A2(new_n757), .A3(new_n754), .A4(new_n751), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n771), .A3(new_n760), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT54), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n743), .A2(new_n766), .A3(new_n576), .A4(new_n616), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n772), .A2(new_n773), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n777), .B1(new_n756), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT53), .A4(new_n774), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n770), .A2(KEYINPUT53), .A3(new_n760), .A4(new_n774), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT117), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n768), .A2(new_n771), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n776), .B1(new_n785), .B2(KEYINPUT54), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n731), .A2(new_n734), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n658), .A2(new_n311), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n319), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n378), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n721), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n587), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n700), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n791), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n716), .A2(new_n659), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n614), .ZN(new_n797));
  INV_X1    g611(.A(new_n640), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n521), .A2(new_n795), .A3(new_n790), .A4(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n375), .A2(new_n799), .A3(new_n592), .A4(new_n590), .ZN(new_n800));
  INV_X1    g614(.A(new_n643), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n579), .A3(new_n674), .A4(new_n794), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n797), .B(new_n800), .C1(KEYINPUT50), .C2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n793), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT51), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n796), .A2(new_n693), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT119), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT119), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT48), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n799), .A2(new_n595), .B1(new_n745), .B2(new_n792), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n786), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n816));
  OAI211_X1 g630(.A(G952), .B(new_n191), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(G953), .B1(new_n815), .B2(KEYINPUT118), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  INV_X1    g635(.A(new_n717), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n521), .A3(new_n481), .A4(new_n319), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(new_n821), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n801), .A3(new_n798), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n817), .A2(new_n818), .A3(new_n826), .ZN(G75));
  AND3_X1   g641(.A1(new_n769), .A2(G902), .A3(new_n775), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n828), .B2(G210), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n451), .A2(new_n438), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(new_n441), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT55), .Z(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n833), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n195), .A2(G952), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G51));
  INV_X1    g651(.A(new_n776), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n769), .A2(KEYINPUT54), .A3(new_n775), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n709), .B(KEYINPUT57), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n840), .A2(new_n841), .B1(new_n300), .B2(new_n310), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n828), .A2(G469), .A3(new_n707), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n836), .B1(new_n842), .B2(new_n843), .ZN(G54));
  NAND3_X1  g658(.A1(new_n828), .A2(KEYINPUT58), .A3(G475), .ZN(new_n845));
  INV_X1    g659(.A(new_n358), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n847), .A2(new_n848), .A3(new_n836), .ZN(G60));
  INV_X1    g663(.A(new_n589), .ZN(new_n850));
  NAND2_X1  g664(.A1(G478), .A2(G902), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT59), .Z(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n786), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n838), .B2(new_n839), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n836), .B1(new_n856), .B2(new_n589), .ZN(new_n857));
  OAI211_X1 g671(.A(KEYINPUT120), .B(new_n850), .C1(new_n786), .C2(new_n852), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(G63));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n860));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n512), .A2(new_n188), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n769), .A2(new_n775), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT122), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n769), .A2(new_n866), .A3(new_n775), .A4(new_n863), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n519), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n836), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n610), .B1(new_n865), .B2(new_n867), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n871), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT61), .A3(new_n869), .A4(new_n868), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(G66));
  AOI21_X1  g689(.A(new_n191), .B1(new_n381), .B2(G224), .ZN(new_n876));
  INV_X1    g690(.A(new_n744), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n877), .B2(new_n195), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n830), .B1(G898), .B2(new_n195), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT123), .Z(new_n880));
  XNOR2_X1  g694(.A(new_n878), .B(new_n880), .ZN(G69));
  AOI21_X1  g695(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n758), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n647), .A2(new_n884), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n735), .A2(new_n728), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n645), .A2(new_n646), .A3(new_n758), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n574), .A2(new_n738), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n889), .A2(new_n629), .A3(new_n716), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n885), .A2(new_n886), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n195), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n536), .B(new_n351), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT124), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n379), .A2(G900), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n735), .A2(new_n698), .A3(new_n704), .ZN(new_n898));
  INV_X1    g712(.A(new_n693), .ZN(new_n899));
  INV_X1    g713(.A(new_n748), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n715), .A2(new_n899), .A3(new_n726), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n728), .A3(new_n758), .A4(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n897), .B(new_n893), .C1(new_n902), .C2(new_n379), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n896), .B1(new_n895), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n883), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n882), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(G72));
  NOR2_X1   g724(.A1(new_n902), .A2(new_n525), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n539), .A3(new_n541), .ZN(new_n912));
  INV_X1    g726(.A(new_n631), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n891), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n836), .B1(new_n914), .B2(new_n744), .ZN(new_n915));
  INV_X1    g729(.A(new_n542), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n560), .ZN(new_n917));
  NAND2_X1  g731(.A1(G472), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT63), .Z(new_n919));
  OR2_X1    g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  MUX2_X1   g734(.A(new_n917), .B(new_n916), .S(KEYINPUT127), .Z(new_n921));
  NAND3_X1  g735(.A1(new_n785), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n915), .A2(new_n920), .A3(new_n922), .ZN(G57));
endmodule


