//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n203), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n217), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G155gat), .B(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  INV_X1    g028(.A(G162gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT2), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(new_n220), .A3(new_n221), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n226), .A3(new_n217), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n202), .B1(new_n215), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n233), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(new_n232), .B2(new_n217), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT29), .B1(new_n211), .B2(new_n212), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n238), .B(KEYINPUT79), .C1(KEYINPUT3), .C2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT73), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n213), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n236), .B2(new_n237), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n214), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n213), .A2(new_n214), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n234), .B1(new_n250), .B2(new_n245), .ZN(new_n251));
  INV_X1    g050(.A(new_n213), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT3), .B1(new_n228), .B2(new_n233), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(KEYINPUT29), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(KEYINPUT78), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT78), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n256), .A3(new_n252), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n255), .A2(new_n257), .B1(G228gat), .B2(G233gat), .ZN(new_n258));
  OAI21_X1  g057(.A(G22gat), .B1(new_n249), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT80), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT77), .B(G50gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT31), .ZN(new_n262));
  XOR2_X1   g061(.A(G78gat), .B(G106gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(new_n257), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n265), .A2(new_n242), .B1(new_n248), .B2(new_n241), .ZN(new_n266));
  INV_X1    g065(.A(G22gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n260), .A2(new_n264), .B1(new_n268), .B2(new_n259), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270));
  AND4_X1   g069(.A1(new_n270), .A2(new_n268), .A3(new_n259), .A4(new_n264), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G169gat), .ZN(new_n276));
  INV_X1    g075(.A(G176gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n280), .B2(KEYINPUT23), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(KEYINPUT23), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT25), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n284), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n294), .B(new_n295), .C1(G183gat), .C2(G190gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n284), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n290), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n287), .A2(KEYINPUT27), .A3(new_n288), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(G190gat), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n304), .B1(new_n308), .B2(KEYINPUT28), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n278), .B1(KEYINPUT26), .B2(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n311), .A2(KEYINPUT26), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n312), .A2(new_n313), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n309), .A2(KEYINPUT67), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT67), .B1(new_n309), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n302), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G226gat), .ZN(new_n318));
  INV_X1    g117(.A(G233gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n283), .A2(new_n297), .B1(new_n300), .B2(new_n284), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n309), .B2(new_n314), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n320), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n322), .A2(new_n325), .A3(new_n244), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n290), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n290), .B1(new_n332), .B2(new_n306), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n313), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n292), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n327), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n309), .A2(KEYINPUT67), .A3(new_n314), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n320), .A3(new_n302), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n321), .B1(new_n342), .B2(new_n323), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n252), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n275), .B1(new_n326), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n320), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n343), .B1(new_n317), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n213), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n325), .A3(new_n244), .ZN(new_n349));
  INV_X1    g148(.A(new_n275), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(KEYINPUT30), .A3(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n317), .A2(new_n321), .B1(new_n324), .B2(new_n320), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n353), .A2(new_n244), .B1(new_n347), .B2(new_n213), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n350), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  OR2_X1    g156(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(G134gat), .A3(new_n359), .ZN(new_n360));
  OR2_X1    g159(.A1(G127gat), .A2(G134gat), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  INV_X1    g164(.A(G120gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(G113gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n364), .B2(G120gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n371), .B(new_n372), .C1(G113gat), .C2(new_n366), .ZN(new_n373));
  NAND2_X1  g172(.A1(G127gat), .A2(G134gat), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT1), .B1(new_n361), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n228), .A2(KEYINPUT3), .A3(new_n233), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n246), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n362), .A2(new_n368), .B1(new_n373), .B2(new_n375), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n381), .A2(new_n234), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n381), .B2(new_n234), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n379), .B(new_n380), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT75), .B(KEYINPUT5), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  INV_X1    g188(.A(G85gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n238), .A2(new_n377), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n381), .A2(new_n234), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n380), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n385), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n388), .B(new_n394), .C1(new_n400), .C2(new_n387), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n385), .A2(new_n387), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n387), .B1(new_n385), .B2(new_n399), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n393), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(KEYINPUT76), .B(KEYINPUT6), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n402), .A2(new_n403), .A3(new_n393), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n357), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n272), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT37), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n348), .A2(new_n349), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n275), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n348), .B2(new_n349), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT84), .B(KEYINPUT38), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT37), .B1(new_n326), .B2(new_n344), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n275), .A3(new_n414), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT84), .B1(new_n420), .B2(KEYINPUT38), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n350), .B1(new_n354), .B2(new_n413), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n353), .A2(new_n244), .B1(new_n347), .B2(new_n213), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT38), .B1(new_n424), .B2(KEYINPUT37), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n423), .A2(new_n425), .B1(new_n354), .B2(new_n350), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n402), .A2(new_n403), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n405), .B1(new_n427), .B2(new_n394), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT83), .B1(new_n428), .B2(new_n404), .ZN(new_n429));
  AND4_X1   g228(.A1(KEYINPUT83), .A2(new_n401), .A3(new_n404), .A4(new_n406), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(new_n409), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n260), .A2(new_n264), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n268), .A2(new_n259), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n268), .A2(new_n259), .A3(new_n270), .A4(new_n264), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n398), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(KEYINPUT39), .C1(new_n398), .C2(new_n397), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n441), .A3(new_n398), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n442), .A2(new_n443), .A3(new_n393), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n442), .B2(new_n393), .ZN(new_n445));
  OAI221_X1 g244(.A(new_n440), .B1(KEYINPUT82), .B2(KEYINPUT40), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n440), .B(new_n449), .C1(new_n444), .C2(new_n445), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n401), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n437), .B1(new_n453), .B2(new_n357), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n412), .B1(new_n432), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n317), .A2(new_n377), .ZN(new_n456));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n340), .A2(new_n381), .A3(new_n302), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT34), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n457), .B(KEYINPUT64), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT34), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(new_n465), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT71), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT70), .B(G15gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(G43gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G71gat), .B(G99gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n462), .B1(new_n456), .B2(new_n458), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(KEYINPUT33), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n458), .ZN(new_n478));
  AOI221_X4 g277(.A(new_n475), .B1(KEYINPUT33), .B2(new_n472), .C1(new_n478), .C2(new_n463), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n466), .B(new_n468), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n476), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n381), .B1(new_n340), .B2(new_n302), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n377), .B(new_n323), .C1(new_n338), .C2(new_n339), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n463), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n487), .A3(new_n472), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n460), .A2(new_n461), .A3(new_n465), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n461), .B1(new_n460), .B2(new_n465), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n481), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT36), .B1(new_n480), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT72), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n480), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n481), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(KEYINPUT72), .A3(new_n466), .A4(new_n468), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n497), .B2(KEYINPUT36), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT35), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n272), .B1(new_n494), .B2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(new_n411), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n437), .A2(new_n499), .A3(new_n357), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n491), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n428), .A2(KEYINPUT83), .A3(new_n404), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n407), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n505), .A2(new_n507), .B1(new_n408), .B2(new_n405), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n503), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  OAI22_X1  g308(.A1(new_n455), .A2(new_n498), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G176gat), .B(G204gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G230gat), .A2(G233gat), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516));
  INV_X1    g315(.A(G64gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(G57gat), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT89), .B1(new_n519), .B2(G64gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(G64gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT90), .ZN(new_n523));
  NAND2_X1  g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  OR2_X1    g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n524), .B(new_n525), .C1(new_n529), .C2(new_n526), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n532), .A2(new_n533), .B1(G85gat), .B2(G92gat), .ZN(new_n534));
  AOI211_X1 g333(.A(KEYINPUT91), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(G85gat), .B(G92gat), .C1(KEYINPUT91), .C2(KEYINPUT7), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(KEYINPUT91), .B2(KEYINPUT7), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT96), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  OR3_X1    g341(.A1(new_n536), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n536), .B2(new_n538), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT10), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n543), .A3(new_n544), .A4(new_n539), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n543), .A2(KEYINPUT92), .A3(new_n544), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT92), .B1(new_n543), .B2(new_n544), .ZN(new_n552));
  OAI211_X1 g351(.A(KEYINPUT10), .B(new_n531), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n515), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n514), .B1(new_n546), .B2(new_n548), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n513), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  INV_X1    g356(.A(new_n513), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT97), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  NOR4_X1   g359(.A1(new_n554), .A2(new_n560), .A3(new_n555), .A4(new_n513), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n556), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT16), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(G1gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n566), .B(new_n567), .C1(G1gat), .C2(new_n564), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(G8gat), .C1(new_n567), .C2(new_n566), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n564), .A2(G1gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n570), .B2(KEYINPUT88), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n571), .B(new_n572), .C1(KEYINPUT88), .C2(new_n566), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(G29gat), .A2(G36gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G43gat), .B(G50gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G43gat), .B(G50gat), .Z(new_n584));
  INV_X1    g383(.A(KEYINPUT15), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT86), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n578), .B(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n586), .A2(new_n577), .A3(new_n581), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n574), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n574), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(KEYINPUT17), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n574), .B(new_n590), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n595), .B(KEYINPUT13), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n596), .A2(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n594), .A2(KEYINPUT18), .A3(new_n595), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n604));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G169gat), .B(G197gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(new_n609), .A3(new_n602), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n563), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n531), .B1(KEYINPUT21), .B2(new_n574), .ZN(new_n615));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n286), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G211gat), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n574), .A2(KEYINPUT21), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n617), .A2(new_n620), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n621), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n621), .B2(new_n626), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n590), .B1(new_n551), .B2(new_n552), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(KEYINPUT41), .ZN(new_n639));
  INV_X1    g438(.A(new_n552), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n593), .A2(new_n640), .A3(new_n550), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n638), .B(new_n639), .C1(new_n641), .C2(KEYINPUT93), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n551), .A2(new_n552), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n593), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n637), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n638), .A2(new_n639), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(KEYINPUT93), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n643), .A3(new_n593), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n636), .ZN(new_n650));
  XNOR2_X1  g449(.A(G134gat), .B(G162gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n646), .B2(new_n650), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n635), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n634), .A3(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n614), .A2(new_n630), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n510), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n410), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(new_n357), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(KEYINPUT98), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(KEYINPUT98), .ZN(new_n674));
  OAI221_X1 g473(.A(new_n671), .B1(new_n572), .B2(new_n666), .C1(new_n673), .C2(new_n674), .ZN(G1325gat));
  INV_X1    g474(.A(new_n504), .ZN(new_n676));
  AOI21_X1  g475(.A(G15gat), .B1(new_n661), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n498), .A2(G15gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT100), .Z(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n661), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n272), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  AND2_X1   g482(.A1(new_n510), .A2(new_n659), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n614), .A2(new_n629), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(G29gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n662), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n455), .A2(new_n498), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n502), .B2(new_n509), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n508), .A2(new_n504), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n694), .A2(new_n499), .A3(new_n357), .A4(new_n437), .ZN(new_n695));
  AOI211_X1 g494(.A(new_n411), .B(new_n272), .C1(new_n494), .C2(new_n496), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n695), .B(KEYINPUT101), .C1(new_n696), .C2(new_n499), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n691), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n656), .A2(new_n658), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n690), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n702), .A2(new_n662), .A3(new_n685), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n689), .B1(new_n687), .B2(new_n703), .ZN(G1328gat));
  INV_X1    g503(.A(G36gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n686), .A2(new_n705), .A3(new_n665), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  AND3_X1   g506(.A1(new_n702), .A2(new_n665), .A3(new_n685), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n705), .B2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n686), .A2(new_n710), .A3(new_n676), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n702), .A2(new_n498), .A3(new_n685), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1330gat));
  NAND3_X1  g514(.A1(new_n702), .A2(new_n272), .A3(new_n685), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G50gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n437), .A2(G50gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n686), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n717), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT102), .B(KEYINPUT48), .Z(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(G1331gat));
  NAND2_X1  g524(.A1(new_n693), .A2(new_n697), .ZN(new_n726));
  INV_X1    g525(.A(new_n691), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n630), .A2(new_n659), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n611), .A2(new_n612), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n730), .A3(new_n562), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n410), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n519), .ZN(G1332gat));
  XOR2_X1   g534(.A(new_n357), .B(KEYINPUT105), .Z(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n698), .A2(KEYINPUT104), .A3(new_n731), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(G1333gat));
  NOR3_X1   g543(.A1(new_n733), .A2(G71gat), .A3(new_n504), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n738), .A2(new_n739), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n498), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(G71gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n272), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n699), .B1(new_n726), .B2(new_n727), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n629), .A2(new_n613), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n757), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n698), .A2(new_n699), .A3(new_n759), .A4(new_n754), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(new_n390), .A3(new_n662), .A4(new_n562), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n563), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n702), .A2(new_n662), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n390), .B2(new_n764), .ZN(G1336gat));
  NOR2_X1   g564(.A1(new_n737), .A2(G92gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n562), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n700), .A2(new_n701), .A3(new_n665), .A4(new_n763), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT107), .B1(new_n770), .B2(KEYINPUT52), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n772), .B(new_n773), .C1(new_n767), .C2(new_n769), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n700), .A2(new_n701), .A3(new_n736), .A4(new_n763), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(new_n776), .B2(G92gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n775), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n767), .A2(new_n775), .A3(new_n777), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n771), .A2(new_n774), .B1(new_n778), .B2(new_n779), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n702), .A2(new_n498), .A3(new_n763), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G99gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n504), .A2(G99gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n562), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n437), .A2(G106gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n761), .A2(new_n562), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n700), .A2(new_n701), .A3(new_n272), .A4(new_n763), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT109), .B(G106gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n792), .B(new_n793), .Z(G1339gat));
  NAND2_X1  g593(.A1(new_n549), .A2(new_n553), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n514), .ZN(new_n796));
  INV_X1    g595(.A(new_n555), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n797), .A3(new_n558), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n560), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n557), .A2(KEYINPUT97), .A3(new_n558), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n594), .A2(new_n595), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n598), .A2(new_n600), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n608), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n612), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n549), .A2(new_n553), .A3(new_n515), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n796), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n558), .B1(new_n554), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n807), .B2(new_n810), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n801), .B(new_n805), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n629), .B1(new_n813), .B2(new_n659), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n613), .B(new_n801), .C1(new_n811), .C2(new_n812), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n562), .A2(new_n805), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n699), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n730), .A2(new_n801), .A3(new_n556), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n729), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT111), .A3(new_n437), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n814), .A2(new_n817), .B1(new_n729), .B2(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(new_n272), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n736), .A2(new_n410), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n676), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n730), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n825), .A2(new_n410), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n500), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n736), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n364), .A3(new_n613), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n834), .ZN(G1340gat));
  OAI21_X1  g634(.A(G120gat), .B1(new_n829), .B2(new_n563), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n366), .A3(new_n562), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  AND2_X1   g637(.A1(new_n358), .A2(new_n359), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n829), .B2(new_n630), .ZN(new_n840));
  INV_X1    g639(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n833), .A2(new_n841), .A3(new_n629), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT112), .ZN(G1342gat));
  NOR4_X1   g643(.A1(new_n832), .A2(G134gat), .A3(new_n665), .A4(new_n699), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT56), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n829), .B2(new_n699), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1343gat));
  NOR3_X1   g647(.A1(new_n498), .A2(new_n410), .A3(new_n736), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n822), .B2(new_n272), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n825), .A2(new_n851), .A3(new_n437), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G141gat), .B1(new_n853), .B2(new_n730), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n498), .A2(new_n437), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n831), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n736), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n218), .A3(new_n613), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n853), .A2(KEYINPUT113), .ZN(new_n861));
  INV_X1    g660(.A(new_n849), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n272), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n851), .B1(new_n825), .B2(new_n437), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n730), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT114), .B1(new_n868), .B2(new_n218), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n865), .A2(new_n866), .ZN(new_n870));
  AOI211_X1 g669(.A(KEYINPUT113), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n613), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(G141gat), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n869), .A2(new_n874), .A3(new_n858), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n860), .B1(new_n875), .B2(new_n859), .ZN(G1344gat));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n219), .A3(new_n562), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n867), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n562), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n219), .A2(KEYINPUT59), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT116), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n852), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n849), .B(KEYINPUT115), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n883), .A2(new_n885), .A3(new_n562), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT117), .B(new_n877), .C1(new_n881), .C2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n879), .B2(new_n880), .ZN(new_n891));
  INV_X1    g690(.A(new_n877), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n893), .ZN(G1345gat));
  AOI21_X1  g693(.A(G155gat), .B1(new_n857), .B2(new_n629), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n630), .A2(new_n229), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n878), .B2(new_n896), .ZN(G1346gat));
  AOI21_X1  g696(.A(new_n699), .B1(new_n861), .B2(new_n867), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n659), .A2(new_n230), .A3(new_n357), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n898), .A2(new_n230), .B1(new_n856), .B2(new_n899), .ZN(G1347gat));
  NAND3_X1  g699(.A1(new_n676), .A2(new_n410), .A3(new_n665), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n827), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT119), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n827), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n730), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n825), .A2(new_n662), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(new_n500), .A3(new_n736), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n276), .A3(new_n613), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(G1348gat));
  NOR3_X1   g711(.A1(new_n907), .A2(new_n277), .A3(new_n563), .ZN(new_n913));
  AOI21_X1  g712(.A(G176gat), .B1(new_n910), .B2(new_n562), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n303), .A3(new_n629), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n904), .A2(new_n629), .A3(new_n906), .ZN(new_n919));
  INV_X1    g718(.A(new_n289), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(G1350gat));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n659), .A3(new_n906), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(G190gat), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n925), .B2(G190gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n925), .A2(G190gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(KEYINPUT61), .A3(new_n927), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n910), .A2(new_n290), .A3(new_n659), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(G1351gat));
  AND2_X1   g734(.A1(new_n883), .A2(new_n885), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n498), .A2(new_n662), .A3(new_n357), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n730), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n855), .A2(new_n736), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(KEYINPUT122), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n941), .A2(new_n909), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n613), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n939), .A2(new_n945), .ZN(G1352gat));
  XNOR2_X1  g745(.A(KEYINPUT123), .B(G204gat), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n563), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n562), .A3(new_n937), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n947), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n629), .A3(new_n937), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G211gat), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT126), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n957), .A2(new_n962), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n205), .A3(new_n629), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1354gat));
  AND2_X1   g765(.A1(new_n938), .A2(KEYINPUT127), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n659), .B1(new_n938), .B2(KEYINPUT127), .ZN(new_n968));
  OAI21_X1  g767(.A(G218gat), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n943), .A2(new_n206), .A3(new_n659), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1355gat));
endmodule


