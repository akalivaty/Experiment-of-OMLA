//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT75), .B1(new_n190), .B2(G125), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G140), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n194), .A2(new_n197), .B1(G125), .B2(new_n190), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n198), .B2(new_n192), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G140), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT19), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n191), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n204), .C1(new_n198), .C2(new_n203), .ZN(new_n205));
  NOR2_X1   g019(.A1(G237), .A2(G953), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(G143), .A3(G214), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(G143), .B1(new_n206), .B2(G214), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G237), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G214), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n207), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n205), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n191), .A2(new_n202), .A3(new_n201), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n198), .B2(new_n201), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n207), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT18), .A3(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT18), .A2(G131), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n215), .A2(new_n207), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G113), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n210), .A2(new_n233), .A3(new_n217), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n201), .B(new_n193), .C1(new_n198), .C2(new_n192), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n222), .A2(KEYINPUT17), .A3(G131), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n200), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n230), .A3(new_n226), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(G475), .A2(G902), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n189), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  AOI211_X1 g056(.A(KEYINPUT20), .B(new_n242), .C1(new_n232), .C2(new_n238), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT84), .B(G475), .Z(new_n245));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n226), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n231), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n238), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n230), .B1(new_n237), .B2(new_n226), .ZN(new_n250));
  AOI21_X1  g064(.A(G902), .B1(new_n250), .B2(KEYINPUT85), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n245), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT13), .B1(new_n255), .B2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G128), .B(G143), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G122), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G116), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT86), .ZN(new_n263));
  INV_X1    g077(.A(G107), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G122), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n263), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n260), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n262), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n266), .B(KEYINPUT14), .ZN(new_n272));
  OAI21_X1  g086(.A(G107), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n259), .B(new_n257), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT9), .B(G234), .ZN(new_n277));
  INV_X1    g091(.A(G217), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n277), .A2(new_n278), .A3(G953), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n269), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n269), .B2(new_n276), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n254), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G478), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT15), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G952), .ZN(new_n288));
  AOI211_X1 g102(.A(G953), .B(new_n288), .C1(G234), .C2(G237), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n254), .B(new_n212), .C1(G234), .C2(G237), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT21), .B(G898), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n253), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n297));
  INV_X1    g111(.A(G119), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(G116), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n265), .A2(KEYINPUT68), .A3(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n265), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G113), .ZN(new_n306));
  AND2_X1   g120(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n306), .B1(new_n309), .B2(new_n302), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n264), .A3(G104), .ZN(new_n314));
  INV_X1    g128(.A(G101), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n229), .A2(G107), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n229), .A2(G107), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n264), .A2(G104), .ZN(new_n319));
  OAI21_X1  g133(.A(G101), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G113), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n311), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n312), .A2(new_n314), .A3(new_n316), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G101), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n301), .A2(new_n303), .A3(new_n326), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n301), .B2(new_n303), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(G101), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n335), .A2(KEYINPUT4), .A3(new_n317), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n328), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G122), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n328), .B(new_n338), .C1(new_n334), .C2(new_n336), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n201), .A2(G143), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n214), .A2(G146), .ZN(new_n344));
  AND2_X1   g158(.A1(KEYINPUT0), .A2(G128), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G143), .B(G146), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT66), .A3(new_n345), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n214), .B2(G146), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n343), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT0), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n255), .A3(KEYINPUT64), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT64), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(KEYINPUT0), .B2(G128), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n345), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n196), .B1(new_n351), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n214), .A2(G146), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT65), .B1(new_n201), .B2(G143), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n352), .A2(new_n214), .A3(G146), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n255), .B1(new_n343), .B2(KEYINPUT1), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n364), .B(new_n196), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(G224), .B(new_n212), .C1(new_n362), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n360), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n348), .B(new_n350), .C1(new_n373), .C2(new_n368), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n212), .A2(G224), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n337), .A2(new_n379), .A3(new_n339), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n342), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT80), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n342), .A2(new_n383), .A3(new_n378), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n311), .A2(new_n327), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n317), .A2(new_n320), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n305), .A2(new_n310), .B1(new_n322), .B2(new_n326), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT81), .B1(new_n390), .B2(new_n321), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n332), .A2(new_n388), .ZN(new_n392));
  INV_X1    g206(.A(new_n322), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n310), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n338), .B(KEYINPUT8), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n398), .ZN(new_n402));
  INV_X1    g216(.A(new_n337), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n362), .B2(new_n371), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n375), .A2(new_n370), .A3(new_n404), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n403), .A2(new_n338), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n254), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n385), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n409), .B2(new_n254), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n296), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n254), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT83), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n416), .A2(new_n295), .A3(new_n385), .A4(new_n411), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n188), .B(new_n294), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT32), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n206), .A2(G210), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT27), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT26), .B(G101), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n257), .A2(G137), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n257), .A2(G137), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT67), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G137), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G134), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT11), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(KEYINPUT67), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n429), .A2(new_n435), .A3(G131), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n216), .B1(new_n431), .B2(new_n425), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT69), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n430), .A2(G134), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n431), .B2(new_n433), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n432), .A2(KEYINPUT11), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n426), .B1(new_n428), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n443), .A3(new_n216), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n445));
  INV_X1    g259(.A(new_n437), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n438), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n332), .A2(new_n333), .ZN(new_n449));
  OAI21_X1  g263(.A(G131), .B1(new_n429), .B2(new_n435), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n444), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n361), .A3(new_n351), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n449), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n216), .B1(new_n441), .B2(new_n443), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n436), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n374), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n439), .A2(new_n444), .A3(new_n446), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n456), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n448), .A2(KEYINPUT70), .A3(new_n449), .A4(new_n452), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n453), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n448), .B2(new_n452), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n452), .A2(new_n471), .A3(new_n460), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n456), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n423), .A3(new_n455), .A4(new_n463), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT31), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n455), .A2(new_n463), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(KEYINPUT31), .A3(new_n423), .A4(new_n475), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n424), .A2(new_n470), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(G472), .A2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n419), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n470), .A2(new_n424), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n482), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n448), .A2(new_n452), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT30), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n449), .B1(new_n490), .B2(new_n473), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n455), .A2(new_n463), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n424), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n424), .B(new_n468), .C1(new_n464), .C2(new_n465), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n489), .A2(new_n456), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n455), .A2(new_n463), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT28), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n469), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n423), .A2(KEYINPUT29), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n254), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G472), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n484), .A2(new_n488), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n278), .B1(G234), .B2(new_n254), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT76), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT73), .B1(new_n298), .B2(G128), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT73), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n255), .A3(G119), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n255), .A2(G119), .B1(KEYINPUT72), .B2(KEYINPUT23), .ZN(new_n512));
  AND2_X1   g326(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n509), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n255), .A2(KEYINPUT23), .A3(G119), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G119), .B(G128), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT24), .B(G110), .Z(new_n518));
  OAI22_X1  g332(.A1(new_n516), .A2(G110), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n220), .A3(new_n200), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n517), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n516), .B2(G110), .ZN(new_n523));
  INV_X1    g337(.A(G110), .ZN(new_n524));
  AOI211_X1 g338(.A(KEYINPUT74), .B(new_n524), .C1(new_n514), .C2(new_n515), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n200), .A2(new_n235), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n508), .B(new_n520), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n200), .A2(new_n235), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n533), .B(new_n521), .C1(new_n525), .C2(new_n523), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n508), .B1(new_n534), .B2(new_n520), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n508), .B(new_n531), .C1(new_n534), .C2(new_n520), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n254), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n520), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n528), .A3(new_n531), .ZN(new_n543));
  INV_X1    g357(.A(new_n537), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT25), .A3(new_n254), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n507), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n506), .A2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT77), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n549), .B2(new_n545), .ZN(new_n550));
  OAI21_X1  g364(.A(G221), .B1(new_n277), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n553), .A2(G128), .B1(new_n343), .B2(new_n344), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n363), .A2(new_n343), .A3(new_n344), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n317), .B(new_n320), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n321), .B2(new_n439), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n451), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT12), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n335), .A2(KEYINPUT4), .A3(new_n317), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n560), .A2(new_n351), .A3(new_n331), .A4(new_n361), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n321), .A2(new_n439), .A3(KEYINPUT10), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n561), .A2(new_n458), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n557), .A2(new_n566), .A3(new_n451), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n212), .A2(G227), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n361), .A2(new_n331), .A3(new_n348), .A4(new_n350), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n564), .B(new_n562), .C1(new_n573), .C2(new_n336), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n451), .ZN(new_n575));
  INV_X1    g389(.A(new_n571), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n565), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G469), .B1(new_n578), .B2(G902), .ZN(new_n579));
  INV_X1    g393(.A(G469), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n576), .B1(new_n575), .B2(new_n565), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT78), .ZN(new_n582));
  OAI22_X1  g396(.A1(new_n581), .A2(new_n582), .B1(new_n571), .B2(new_n568), .ZN(new_n583));
  AOI211_X1 g397(.A(KEYINPUT78), .B(new_n576), .C1(new_n575), .C2(new_n565), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n580), .B(new_n254), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n552), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n418), .A2(new_n505), .A3(new_n550), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  OAI21_X1  g402(.A(KEYINPUT33), .B1(new_n281), .B2(new_n282), .ZN(new_n589));
  INV_X1    g403(.A(new_n282), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n280), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n284), .A2(G902), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT89), .B(G478), .Z(new_n595));
  AOI22_X1  g409(.A1(new_n593), .A2(new_n594), .B1(new_n283), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n249), .A2(new_n251), .ZN(new_n598));
  INV_X1    g412(.A(new_n245), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n241), .B2(new_n243), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n292), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n414), .A2(new_n417), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT88), .B1(new_n604), .B2(new_n187), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT88), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n606), .B(new_n188), .C1(new_n414), .C2(new_n417), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT87), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n487), .B2(new_n254), .ZN(new_n612));
  AOI211_X1 g426(.A(G902), .B(new_n610), .C1(new_n485), .C2(new_n486), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n586), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n545), .A2(new_n549), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n615), .A2(new_n547), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  AOI211_X1 g435(.A(KEYINPUT90), .B(new_n189), .C1(new_n239), .C2(new_n240), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n244), .B2(KEYINPUT90), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT91), .B1(new_n598), .B2(new_n599), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n625), .B(new_n245), .C1(new_n249), .C2(new_n251), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(new_n627), .A3(new_n286), .A4(new_n293), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT92), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n605), .B2(new_n607), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n618), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  OR2_X1    g447(.A1(new_n531), .A2(KEYINPUT36), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n634), .A2(KEYINPUT94), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(KEYINPUT94), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n637), .A2(KEYINPUT93), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(KEYINPUT93), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n541), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n638), .A2(new_n534), .A3(new_n520), .A4(new_n639), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n641), .A2(new_n549), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n540), .A2(new_n546), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(new_n506), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n615), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n418), .A2(new_n614), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n290), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n289), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n623), .A2(new_n627), .A3(new_n286), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n645), .A2(new_n615), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n655), .B(new_n505), .C1(new_n605), .C2(new_n607), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XNOR2_X1  g471(.A(new_n653), .B(KEYINPUT39), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n586), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT40), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT97), .Z(new_n661));
  OAI21_X1  g475(.A(new_n423), .B1(new_n491), .B2(new_n492), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n662), .B(new_n254), .C1(new_n423), .C2(new_n499), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n484), .A2(new_n488), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT96), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT96), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n484), .A2(new_n488), .A3(new_n667), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n604), .B(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n645), .A2(new_n286), .A3(new_n601), .A4(new_n187), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  INV_X1    g489(.A(new_n653), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n253), .A2(new_n596), .A3(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n677), .B(new_n586), .C1(new_n547), .C2(new_n643), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n505), .B(new_n679), .C1(new_n605), .C2(new_n607), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(new_n254), .B1(new_n583), .B2(new_n584), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n551), .A3(new_n585), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT98), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n550), .A3(new_n505), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n608), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT41), .B(G113), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND2_X1  g503(.A1(new_n604), .A2(new_n187), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n606), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n188), .B1(new_n414), .B2(new_n417), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT88), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n505), .A2(new_n550), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n695), .A3(new_n629), .A4(new_n685), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT99), .B(G116), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G18));
  NOR2_X1   g512(.A1(new_n645), .A2(new_n294), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n694), .A2(new_n505), .A3(new_n685), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  NAND2_X1  g515(.A1(new_n501), .A2(new_n424), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n483), .B1(new_n702), .B2(new_n486), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n487), .A2(new_n254), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n703), .B1(new_n704), .B2(G472), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n550), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT100), .B1(new_n253), .B2(new_n287), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT100), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n601), .A2(new_n708), .A3(new_n286), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n292), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n694), .A2(new_n706), .A3(new_n685), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  OAI21_X1  g527(.A(new_n685), .B1(new_n605), .B2(new_n607), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT25), .B1(new_n545), .B2(new_n254), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n539), .B(G902), .C1(new_n543), .C2(new_n544), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n506), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n643), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n705), .A2(new_n719), .A3(new_n677), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n196), .ZN(G27));
  NAND3_X1  g536(.A1(new_n414), .A2(new_n187), .A3(new_n417), .ZN(new_n723));
  NAND2_X1  g537(.A1(G469), .A2(G902), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n572), .A2(KEYINPUT101), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n568), .A2(new_n726), .A3(new_n571), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(G469), .A3(new_n577), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n585), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n551), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n505), .A3(new_n550), .A4(new_n677), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  INV_X1    g551(.A(new_n654), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n731), .A2(new_n505), .A3(new_n550), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NOR2_X1   g554(.A1(new_n578), .A2(KEYINPUT45), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n580), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n577), .A4(new_n727), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n724), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n585), .ZN(new_n748));
  OR3_X1    g562(.A1(new_n745), .A2(KEYINPUT103), .A3(new_n746), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT103), .B1(new_n745), .B2(new_n746), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n552), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT104), .B1(new_n752), .B2(new_n658), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  INV_X1    g568(.A(new_n658), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n751), .A2(new_n754), .A3(new_n552), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n253), .A2(new_n597), .A3(KEYINPUT43), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n596), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n253), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n761), .A2(KEYINPUT106), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT106), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n614), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n719), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n723), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n765), .A2(KEYINPUT44), .A3(new_n766), .A4(new_n719), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n757), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n430), .ZN(G39));
  XOR2_X1   g588(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n752), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT47), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n752), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n677), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n505), .A2(new_n550), .A3(new_n780), .A4(new_n723), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT108), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT109), .B(G140), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G42));
  NAND2_X1  g599(.A1(new_n683), .A2(new_n585), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT49), .Z(new_n788));
  NOR4_X1   g602(.A1(new_n601), .A2(new_n596), .A3(new_n188), .A4(new_n552), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n671), .A2(new_n550), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n669), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n765), .A2(new_n289), .A3(new_n706), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n714), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n288), .A3(G953), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n685), .A2(new_n289), .A3(new_n770), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n765), .A2(new_n796), .A3(new_n695), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT48), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n550), .A3(new_n796), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n795), .B(new_n798), .C1(new_n602), .C2(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n787), .A2(new_n551), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n723), .B(new_n793), .C1(new_n779), .C2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n799), .A2(new_n601), .A3(new_n597), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n671), .A2(new_n188), .A3(new_n685), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT114), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n793), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n806), .A2(KEYINPUT114), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n807), .B(new_n809), .C1(new_n793), .C2(new_n805), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n765), .A2(new_n796), .A3(new_n719), .A4(new_n705), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n804), .A2(new_n808), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n800), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n813), .A2(new_n817), .A3(KEYINPUT51), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n817), .B1(new_n813), .B2(KEYINPUT51), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n710), .B1(new_n691), .B2(new_n693), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n719), .A2(new_n676), .A3(new_n730), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n822), .A2(new_n669), .A3(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n656), .B(new_n680), .C1(new_n714), .C2(new_n720), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT52), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n721), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n656), .A2(new_n680), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n669), .A3(new_n823), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n287), .A2(new_n623), .A3(new_n627), .A4(new_n653), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n505), .A2(new_n646), .A3(new_n770), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n719), .A2(new_n586), .A3(new_n833), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n505), .A4(new_n770), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n731), .A2(new_n719), .A3(new_n705), .A4(new_n677), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n739), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n736), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n601), .A2(new_n287), .A3(new_n292), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT111), .B1(new_n692), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n604), .A2(KEYINPUT111), .A3(new_n187), .A4(new_n844), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n614), .A3(new_n617), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n696), .A2(new_n700), .A3(new_n712), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n694), .A2(new_n695), .A3(new_n603), .A4(new_n685), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n614), .A2(new_n692), .A3(new_n603), .A4(new_n617), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n587), .A3(new_n647), .A4(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n843), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n832), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n826), .A2(new_n831), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n505), .A2(new_n699), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n630), .A2(new_n686), .B1(new_n714), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n711), .A2(new_n705), .A3(new_n550), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n614), .A2(new_n847), .A3(new_n617), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n714), .A2(new_n858), .B1(new_n859), .B2(new_n845), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n587), .A2(new_n851), .A3(new_n647), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n687), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n841), .B1(new_n838), .B2(new_n835), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n861), .A2(new_n736), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n855), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n821), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n832), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n855), .B2(new_n865), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n820), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n792), .B1(new_n873), .B2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n212), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n254), .B1(new_n869), .B2(new_n870), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n342), .A2(new_n380), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n378), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(G902), .B1(new_n854), .B2(new_n867), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n878), .A2(KEYINPUT116), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n296), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n883), .B1(new_n888), .B2(new_n890), .ZN(G51));
  XOR2_X1   g705(.A(new_n724), .B(KEYINPUT57), .Z(new_n892));
  NAND3_X1  g706(.A1(new_n868), .A2(new_n871), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n583), .A2(new_n584), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT117), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n744), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n886), .A2(new_n896), .A3(new_n887), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT117), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n877), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(KEYINPUT118), .B(new_n877), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(G54));
  NAND4_X1  g718(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT58), .A4(G475), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n232), .A2(new_n238), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n876), .ZN(G60));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT59), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n872), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n593), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n877), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n869), .B2(new_n870), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n918), .A2(new_n642), .A3(new_n641), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n877), .B1(new_n918), .B2(new_n545), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n919), .A2(new_n920), .B1(KEYINPUT119), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G66));
  INV_X1    g738(.A(G224), .ZN(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n291), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n849), .A2(new_n852), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n880), .B1(G898), .B2(new_n212), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G69));
  AOI21_X1  g744(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n822), .A2(new_n695), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n772), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n753), .B2(new_n756), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n779), .A2(new_n782), .ZN(new_n935));
  INV_X1    g749(.A(new_n825), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n736), .A2(new_n739), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n783), .A2(new_n825), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n940), .A2(new_n941), .A3(new_n934), .A4(new_n937), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n942), .A3(new_n212), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n204), .B1(new_n198), .B2(new_n203), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT120), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT121), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n472), .A2(new_n474), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G900), .A2(G953), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n659), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n602), .B1(new_n287), .B2(new_n601), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT123), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n695), .A2(new_n951), .A3(new_n770), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n757), .B2(new_n772), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(KEYINPUT124), .B(new_n954), .C1(new_n757), .C2(new_n772), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n674), .A2(new_n936), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  OR3_X1    g775(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT62), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n960), .B2(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n783), .B1(new_n960), .B2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n959), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n948), .B1(new_n966), .B2(new_n212), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n950), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n931), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n966), .A2(new_n212), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT125), .B1(new_n972), .B2(new_n948), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n967), .A2(new_n968), .ZN(new_n974));
  INV_X1    g788(.A(new_n931), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n950), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n971), .A2(new_n976), .ZN(G72));
  NAND3_X1  g791(.A1(new_n939), .A2(new_n942), .A3(new_n927), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT63), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n424), .A3(new_n479), .A4(new_n475), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n869), .A2(new_n870), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n493), .B2(new_n476), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n876), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n662), .ZN(new_n988));
  INV_X1    g802(.A(new_n927), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n981), .B1(new_n966), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(G57));
endmodule


