//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT66), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G137), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n462), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n478), .B2(G112), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n467), .A2(new_n468), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n462), .A2(KEYINPUT67), .A3(new_n478), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(new_n485), .B2(G136), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(KEYINPUT68), .B2(G114), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT68), .A2(G114), .ZN(new_n489));
  OAI211_X1 g064(.A(G2104), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n478), .C1(new_n467), .C2(new_n468), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n462), .A2(new_n495), .A3(G138), .A4(new_n478), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(G543), .B1(new_n498), .B2(KEYINPUT69), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT5), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(G543), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  XOR2_X1   g087(.A(new_n512), .B(KEYINPUT70), .Z(new_n513));
  AOI21_X1  g088(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n509), .A2(new_n514), .ZN(G166));
  INV_X1    g090(.A(new_n505), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  INV_X1    g092(.A(new_n508), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n505), .A2(new_n525), .B1(new_n526), .B2(new_n508), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n503), .A2(G64), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n510), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G171));
  NAND2_X1  g106(.A1(new_n518), .A2(G43), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(G81), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n499), .A2(new_n502), .A3(G56), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n510), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n532), .B1(new_n505), .B2(new_n533), .C1(new_n534), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n534), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(new_n516), .A2(G91), .ZN(new_n547));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT9), .B1(new_n508), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n504), .A2(new_n550), .A3(G53), .A4(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n499), .A2(new_n502), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n547), .A2(new_n552), .A3(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  NAND4_X1  g135(.A1(new_n504), .A2(G87), .A3(new_n499), .A4(new_n502), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n504), .A2(G49), .A3(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G74), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n510), .B1(new_n554), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n563), .A2(new_n565), .ZN(G288));
  NAND4_X1  g141(.A1(new_n504), .A2(G86), .A3(new_n499), .A4(new_n502), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n499), .A2(new_n502), .A3(G61), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G305));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n505), .A2(new_n575), .B1(new_n576), .B2(new_n508), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n503), .A2(G60), .ZN(new_n578));
  NAND2_X1  g153(.A1(G72), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n510), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n503), .A2(G92), .A3(new_n504), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n554), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n518), .B2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n583), .B1(new_n592), .B2(G868), .ZN(G321));
  XOR2_X1   g168(.A(G321), .B(KEYINPUT73), .Z(G284));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G168), .B2(new_n595), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(G168), .B2(new_n595), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  OAI21_X1  g175(.A(new_n595), .B1(new_n538), .B2(new_n540), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n591), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g179(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT12), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT74), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT13), .Z(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(G2100), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(G111), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(KEYINPUT75), .B1(new_n612), .B2(G2105), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT75), .B2(new_n611), .ZN(new_n614));
  INV_X1    g189(.A(G123), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n475), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G135), .B2(new_n485), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n609), .A2(new_n610), .A3(new_n618), .ZN(G156));
  INV_X1    g194(.A(G14), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2451), .B(G2454), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT16), .ZN(new_n622));
  XNOR2_X1  g197(.A(G1341), .B(G1348), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G2443), .B(G2446), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT76), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n620), .B1(new_n626), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n626), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT77), .Z(G401));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n639), .A2(new_n637), .A3(new_n640), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n637), .A3(new_n640), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT18), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2100), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n652), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n652), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT79), .Z(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G1981), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  NAND2_X1  g246(.A1(G290), .A2(G16), .ZN(new_n672));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G24), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT80), .ZN(new_n676));
  INV_X1    g251(.A(G1986), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n678), .A3(new_n674), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n676), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G25), .ZN(new_n683));
  INV_X1    g258(.A(G119), .ZN(new_n684));
  NOR2_X1   g259(.A1(G95), .A2(G2105), .ZN(new_n685));
  OAI21_X1  g260(.A(G2104), .B1(new_n478), .B2(G107), .ZN(new_n686));
  OAI22_X1  g261(.A1(new_n475), .A2(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n485), .B2(G131), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n683), .B1(new_n688), .B2(new_n682), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT35), .B(G1991), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n680), .A2(new_n681), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(G305), .A2(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n673), .A2(G6), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT82), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n673), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n673), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n698), .A2(new_n706), .A3(new_n699), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n701), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n673), .A2(G23), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G288), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  OAI21_X1  g288(.A(KEYINPUT33), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n710), .A2(new_n711), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT33), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n710), .A2(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G1976), .ZN(new_n720));
  INV_X1    g295(.A(G1976), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n714), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n708), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT81), .B(KEYINPUT34), .Z(new_n724));
  OAI21_X1  g299(.A(new_n692), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n708), .ZN(new_n726));
  INV_X1    g301(.A(new_n722), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n721), .B1(new_n714), .B2(new_n718), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n724), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT36), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n723), .A2(new_n724), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n692), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G301), .A2(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n673), .A2(G5), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G1961), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n738), .A2(new_n742), .A3(new_n739), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n682), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n485), .A2(G141), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n478), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G129), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n745), .A2(new_n749), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n744), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n741), .A2(new_n743), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  INV_X1    g335(.A(G127), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n482), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n762), .A2(G2105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n483), .A2(new_n484), .ZN(new_n768));
  INV_X1    g343(.A(G139), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(KEYINPUT84), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT84), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n682), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n682), .A2(G33), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n775), .A2(G2072), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(G2072), .B1(new_n775), .B2(new_n776), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n759), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(G164), .A2(G29), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G27), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2078), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n617), .A2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n473), .A2(G29), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT24), .ZN(new_n788));
  INV_X1    g363(.A(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G28), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(KEYINPUT30), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT86), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n793), .B2(KEYINPUT30), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT31), .B(G11), .Z(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n784), .A2(new_n785), .A3(new_n792), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n787), .A2(new_n786), .A3(new_n791), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT87), .Z(new_n802));
  AND2_X1   g377(.A1(new_n673), .A2(G21), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G286), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT85), .B(G1966), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n755), .A2(new_n756), .B1(new_n782), .B2(new_n783), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n800), .A2(new_n802), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT88), .B1(new_n780), .B2(new_n808), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n806), .A2(new_n800), .A3(new_n802), .A4(new_n807), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n758), .A2(new_n777), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT88), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n779), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n682), .A2(G35), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G162), .B2(new_n682), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT29), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G2090), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT89), .Z(new_n818));
  AND2_X1   g393(.A1(new_n673), .A2(G4), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n591), .B2(G16), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1348), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n673), .A2(G20), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT23), .Z(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1956), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n673), .A2(G19), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n541), .B2(new_n673), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n825), .B1(G1341), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n682), .A2(G26), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT28), .ZN(new_n830));
  INV_X1    g405(.A(G128), .ZN(new_n831));
  NOR2_X1   g406(.A1(G104), .A2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n475), .A2(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n485), .B2(G140), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n830), .B1(new_n835), .B2(new_n682), .ZN(new_n836));
  INV_X1    g411(.A(G2067), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n816), .B2(G2090), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n827), .A2(G1341), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n821), .A2(new_n828), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n809), .A2(new_n813), .A3(new_n818), .A4(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT90), .B1(new_n737), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT90), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n845), .B(new_n842), .C1(new_n732), .C2(new_n736), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n737), .A2(new_n843), .ZN(G150));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT92), .B(G55), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n505), .A2(new_n849), .B1(new_n508), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n503), .A2(G67), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n510), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT94), .B(G860), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n591), .A2(new_n599), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT93), .B1(new_n538), .B2(new_n540), .ZN(new_n862));
  INV_X1    g437(.A(new_n533), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n516), .A2(new_n863), .B1(G43), .B2(new_n518), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n537), .A2(new_n534), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n539), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n862), .A2(new_n855), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n855), .B1(new_n862), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n861), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n856), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n858), .B1(new_n873), .B2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n754), .A2(new_n835), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n749), .A2(new_n750), .A3(new_n753), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(G141), .B2(new_n485), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n485), .A2(G140), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n834), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n494), .A2(new_n496), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n490), .A2(new_n491), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n877), .A2(new_n881), .A3(G164), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n773), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n771), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n688), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n688), .A2(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n606), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(new_n606), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(G2104), .B1(new_n478), .B2(G118), .ZN(new_n901));
  INV_X1    g476(.A(G106), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n478), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT96), .ZN(new_n904));
  INV_X1    g479(.A(G130), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n475), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n748), .A2(KEYINPUT96), .A3(G130), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n485), .A2(G142), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n900), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n896), .A2(new_n899), .A3(new_n910), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT95), .B1(new_n770), .B2(new_n773), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n886), .B2(new_n888), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n891), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n913), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n770), .B1(new_n889), .B2(new_n773), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT98), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n891), .A2(new_n914), .A3(KEYINPUT99), .A4(new_n917), .ZN(new_n926));
  OAI211_X1 g501(.A(KEYINPUT98), .B(new_n921), .C1(new_n922), .C2(new_n916), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n920), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n617), .B(new_n473), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(G162), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n933), .B2(new_n918), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n931), .A2(KEYINPUT40), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT40), .B1(new_n931), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(G395));
  OAI21_X1  g512(.A(new_n870), .B1(G559), .B2(new_n591), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n547), .A2(new_n557), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n591), .A2(new_n552), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(G299), .A2(new_n586), .A3(new_n590), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(KEYINPUT41), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n602), .B1(new_n868), .B2(new_n869), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n938), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n942), .B(KEYINPUT100), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n938), .B2(new_n947), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n951));
  OR3_X1    g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n581), .B(G305), .ZN(new_n953));
  XNOR2_X1  g528(.A(G166), .B(G288), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n953), .B(new_n954), .Z(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n948), .B2(new_n950), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n952), .B2(new_n956), .ZN(new_n958));
  OAI21_X1  g533(.A(G868), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n855), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n595), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(G295));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n961), .ZN(G331));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  XNOR2_X1  g539(.A(G286), .B(G171), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n868), .B2(new_n869), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n862), .A2(new_n867), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n960), .ZN(new_n968));
  XNOR2_X1  g543(.A(G301), .B(G286), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n862), .A2(new_n855), .A3(new_n867), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT102), .B(new_n965), .C1(new_n868), .C2(new_n869), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n946), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n955), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n966), .A2(new_n971), .A3(new_n942), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G37), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n964), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT41), .B1(new_n940), .B2(new_n941), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT103), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n945), .B(KEYINPUT104), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n984), .A2(new_n985), .B1(new_n966), .B2(new_n971), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n949), .B1(new_n973), .B2(new_n974), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n955), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(KEYINPUT43), .A3(new_n979), .A4(new_n978), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT44), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n980), .B2(new_n981), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n988), .A2(new_n964), .A3(new_n979), .A4(new_n978), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n996), .ZN(G397));
  AOI21_X1  g572(.A(new_n478), .B1(new_n463), .B2(new_n464), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT105), .B(G40), .Z(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(new_n471), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n883), .B2(new_n884), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n837), .ZN(new_n1002));
  INV_X1    g577(.A(new_n999), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n466), .A2(new_n472), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n885), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1008), .A3(KEYINPUT110), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n885), .A2(new_n1007), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1004), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1002), .B1(new_n1013), .B2(G1348), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n592), .ZN(new_n1015));
  NAND2_X1  g590(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G299), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT119), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(G299), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1004), .B1(new_n1010), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1025), .A2(KEYINPUT120), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(new_n1026), .A3(new_n1000), .A4(new_n1027), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1005), .A2(new_n1008), .A3(new_n1000), .ZN(new_n1033));
  INV_X1    g608(.A(G1956), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND4_X1   g610(.A1(new_n1023), .A2(new_n1028), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1015), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1028), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT121), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1031), .A2(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n1028), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1023), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n591), .B(new_n1002), .C1(new_n1013), .C2(G1348), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1015), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT60), .ZN(new_n1047));
  INV_X1    g622(.A(G1996), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1025), .A2(new_n1048), .A3(new_n1026), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1025), .A2(KEYINPUT122), .A3(new_n1048), .A4(new_n1026), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT58), .B(G1341), .Z(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1010), .B2(new_n1004), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n541), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT59), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(KEYINPUT59), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT59), .A4(new_n541), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1047), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1023), .B1(new_n1040), .B2(new_n1028), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1036), .B2(new_n1064), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1014), .A2(KEYINPUT60), .A3(new_n591), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1040), .A2(new_n1023), .A3(new_n1028), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT61), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1065), .B(new_n1066), .C1(new_n1043), .C2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1044), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(G171), .B(KEYINPUT54), .Z(new_n1071));
  NAND3_X1  g646(.A1(new_n1029), .A2(G40), .A3(G160), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT125), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1029), .A2(new_n1074), .A3(G40), .A4(G160), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1026), .A2(KEYINPUT53), .A3(new_n783), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1071), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1029), .A2(new_n1026), .A3(new_n783), .A4(new_n1000), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1078), .B(new_n1081), .C1(G1961), .C2(new_n1013), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1025), .A2(KEYINPUT53), .A3(new_n783), .A4(new_n1026), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1081), .B(new_n1083), .C1(new_n1013), .C2(G1961), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1071), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT111), .B(G8), .Z(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G286), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  AOI211_X1 g665(.A(G2084), .B(new_n1004), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1966), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n786), .A3(new_n1000), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1092), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1089), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(KEYINPUT51), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT51), .B1(G286), .B2(new_n1088), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n509), .B2(new_n514), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT55), .Z(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1971), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n1107));
  AOI21_X1  g682(.A(G2090), .B1(new_n1033), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1005), .A2(new_n1008), .A3(KEYINPUT115), .A4(new_n1000), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1110), .B2(new_n1087), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n721), .B1(new_n563), .B2(new_n565), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1087), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1116));
  OR3_X1    g691(.A1(new_n563), .A2(new_n721), .A3(new_n565), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1112), .A2(new_n1118), .A3(new_n1113), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT49), .ZN(new_n1121));
  INV_X1    g696(.A(G1981), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n569), .B2(new_n573), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n567), .A2(new_n568), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n510), .B1(new_n570), .B2(new_n571), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(new_n1125), .A3(G1981), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1121), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n569), .A2(new_n1122), .A3(new_n573), .ZN(new_n1128));
  OAI21_X1  g703(.A(G1981), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT49), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1116), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1120), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1116), .A2(KEYINPUT112), .A3(new_n1117), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT112), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(new_n1113), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1004), .A2(G2090), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1104), .B(G8), .C1(new_n1106), .C2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1111), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1086), .A2(new_n1102), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1070), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(KEYINPUT63), .ZN(new_n1143));
  OAI211_X1 g718(.A(G168), .B(new_n1088), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(G8), .B1(new_n1138), .B2(new_n1106), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1105), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1147), .A2(new_n1136), .A3(KEYINPUT116), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT116), .B1(new_n1147), .B2(new_n1136), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1145), .B(KEYINPUT117), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT62), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1084), .A2(G171), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1158), .A2(new_n1111), .A3(new_n1136), .A4(new_n1139), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1098), .A2(KEYINPUT62), .A3(new_n1101), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1139), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1136), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1131), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1116), .B1(new_n1165), .B2(new_n1126), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT114), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT114), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1160), .A2(new_n1161), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1142), .A2(new_n1156), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n879), .B(new_n1048), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1029), .A2(new_n1004), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT106), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n880), .A2(G2067), .A3(new_n834), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n835), .A2(new_n837), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(G2067), .B1(new_n880), .B2(new_n834), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n835), .A2(new_n837), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(KEYINPUT106), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1182), .A3(new_n1174), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT107), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1175), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT108), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(KEYINPUT108), .B(new_n1175), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1190));
  INV_X1    g765(.A(new_n688), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1191), .A2(new_n690), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n690), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1174), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n581), .B(new_n677), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1174), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1189), .A2(new_n1190), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT109), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1172), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1174), .A2(new_n677), .A3(new_n581), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1189), .A2(new_n1190), .A3(new_n1194), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1174), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1204), .A2(G1996), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT46), .Z(new_n1206));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1204), .B1(new_n1208), .B2(new_n879), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1206), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT47), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1205), .B(KEYINPUT46), .ZN(new_n1213));
  OAI21_X1  g788(.A(KEYINPUT127), .B1(new_n1213), .B2(new_n1209), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1212), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1203), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT126), .B1(new_n1218), .B2(new_n1181), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1219), .A2(new_n1204), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1218), .A2(KEYINPUT126), .A3(new_n1181), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1200), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g798(.A(new_n460), .ZN(new_n1225));
  NAND4_X1  g799(.A1(new_n670), .A2(new_n1225), .A3(new_n635), .A4(new_n649), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n1226), .B1(new_n931), .B2(new_n934), .ZN(new_n1227));
  AND2_X1   g801(.A1(new_n1227), .A2(new_n994), .ZN(G308));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n994), .ZN(G225));
endmodule


