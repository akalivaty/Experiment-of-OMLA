

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U558 ( .A(n785), .B(KEYINPUT32), .ZN(n812) );
  AND2_X2 U559 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X2 U560 ( .A1(G2104), .A2(n548), .ZN(n896) );
  XOR2_X1 U561 ( .A(KEYINPUT65), .B(n536), .Z(G160) );
  XNOR2_X1 U562 ( .A(KEYINPUT17), .B(n531), .ZN(n524) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n736) );
  OR2_X1 U564 ( .A1(n792), .A2(n791), .ZN(n813) );
  INV_X1 U565 ( .A(KEYINPUT107), .ZN(n807) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n655) );
  INV_X1 U567 ( .A(n524), .ZN(n900) );
  NOR2_X1 U568 ( .A1(G651), .A2(n651), .ZN(n661) );
  INV_X1 U569 ( .A(G2105), .ZN(n548) );
  AND2_X1 U570 ( .A1(G2104), .A2(G101), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n548), .A2(n525), .ZN(n526) );
  XNOR2_X1 U572 ( .A(n526), .B(KEYINPUT66), .ZN(n528) );
  INV_X1 U573 ( .A(KEYINPUT23), .ZN(n527) );
  XNOR2_X1 U574 ( .A(n528), .B(n527), .ZN(n530) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n895) );
  NAND2_X1 U576 ( .A1(G113), .A2(n895), .ZN(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n535) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  NAND2_X1 U579 ( .A1(G137), .A2(n900), .ZN(n533) );
  NAND2_X1 U580 ( .A1(G125), .A2(n896), .ZN(n532) );
  NAND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n536) );
  AND2_X1 U583 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U584 ( .A(G120), .ZN(G236) );
  INV_X1 U585 ( .A(G69), .ZN(G235) );
  INV_X1 U586 ( .A(G108), .ZN(G238) );
  INV_X1 U587 ( .A(G132), .ZN(G219) );
  INV_X1 U588 ( .A(G82), .ZN(G220) );
  NAND2_X1 U589 ( .A1(G90), .A2(n655), .ZN(n538) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n651) );
  INV_X1 U591 ( .A(G651), .ZN(n542) );
  NOR2_X1 U592 ( .A1(n651), .A2(n542), .ZN(n656) );
  NAND2_X1 U593 ( .A1(G77), .A2(n656), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U595 ( .A(n539), .B(KEYINPUT9), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G52), .A2(n661), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n547) );
  NOR2_X1 U598 ( .A1(G543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U599 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n543) );
  XNOR2_X1 U600 ( .A(n544), .B(n543), .ZN(n654) );
  NAND2_X1 U601 ( .A1(n654), .A2(G64), .ZN(n545) );
  XOR2_X1 U602 ( .A(KEYINPUT68), .B(n545), .Z(n546) );
  NOR2_X1 U603 ( .A1(n547), .A2(n546), .ZN(G171) );
  NAND2_X1 U604 ( .A1(G138), .A2(n900), .ZN(n550) );
  AND2_X1 U605 ( .A1(n548), .A2(G2104), .ZN(n903) );
  NAND2_X1 U606 ( .A1(G102), .A2(n903), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U608 ( .A1(G114), .A2(n895), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G126), .A2(n896), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n554), .A2(n553), .ZN(G164) );
  NAND2_X1 U612 ( .A1(G63), .A2(n654), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G51), .A2(n661), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(KEYINPUT75), .Z(n557) );
  XNOR2_X1 U616 ( .A(n558), .B(n557), .ZN(n565) );
  NAND2_X1 U617 ( .A1(G89), .A2(n655), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(KEYINPUT74), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G76), .A2(n656), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT5), .B(n563), .Z(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n568) );
  XNOR2_X1 U624 ( .A(KEYINPUT77), .B(KEYINPUT7), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT76), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n568), .B(n567), .ZN(G168) );
  XOR2_X1 U627 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G567), .ZN(n689) );
  NOR2_X1 U631 ( .A1(n689), .A2(G223), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n570), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n572) );
  NAND2_X1 U634 ( .A1(G56), .A2(n654), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n572), .B(n571), .ZN(n579) );
  XNOR2_X1 U636 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n655), .A2(G81), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G68), .A2(n656), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n661), .A2(G43), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n1002) );
  INV_X1 U645 ( .A(G860), .ZN(n603) );
  OR2_X1 U646 ( .A1(n1002), .A2(n603), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G301), .A2(G868), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n582), .B(KEYINPUT72), .ZN(n592) );
  INV_X1 U650 ( .A(G868), .ZN(n608) );
  NAND2_X1 U651 ( .A1(G66), .A2(n654), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G92), .A2(n655), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G79), .A2(n656), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G54), .A2(n661), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n589), .Z(n590) );
  XNOR2_X1 U659 ( .A(KEYINPUT73), .B(n590), .ZN(n985) );
  NAND2_X1 U660 ( .A1(n608), .A2(n985), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G78), .A2(n656), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G53), .A2(n661), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G65), .A2(n654), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G91), .A2(n655), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U670 ( .A1(G299), .A2(n608), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT78), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U675 ( .A(n985), .ZN(n921) );
  NAND2_X1 U676 ( .A1(n604), .A2(n921), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT16), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n606) );
  XNOR2_X1 U679 ( .A(n607), .B(n606), .ZN(G148) );
  NOR2_X1 U680 ( .A1(n985), .A2(n608), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT82), .B(n609), .Z(n610) );
  NOR2_X1 U682 ( .A1(G559), .A2(n610), .ZN(n613) );
  NOR2_X1 U683 ( .A1(G868), .A2(n1002), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT81), .B(n611), .Z(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U686 ( .A1(G135), .A2(n900), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G111), .A2(n895), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n896), .A2(G123), .ZN(n616) );
  XOR2_X1 U690 ( .A(KEYINPUT18), .B(n616), .Z(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n903), .A2(G99), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n940) );
  XNOR2_X1 U694 ( .A(n940), .B(G2096), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT83), .ZN(n623) );
  INV_X1 U696 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G559), .A2(n921), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n1002), .B(n624), .ZN(n670) );
  NOR2_X1 U700 ( .A1(n670), .A2(G860), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G67), .A2(n654), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G55), .A2(n661), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G93), .A2(n655), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G80), .A2(n656), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n673) );
  XNOR2_X1 U708 ( .A(n631), .B(n673), .ZN(G145) );
  NAND2_X1 U709 ( .A1(n654), .A2(G62), .ZN(n632) );
  XOR2_X1 U710 ( .A(KEYINPUT85), .B(n632), .Z(n634) );
  NAND2_X1 U711 ( .A1(n661), .A2(G50), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U713 ( .A(KEYINPUT86), .B(n635), .Z(n639) );
  NAND2_X1 U714 ( .A1(G88), .A2(n655), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G75), .A2(n656), .ZN(n636) );
  AND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(G303) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G73), .A2(n656), .ZN(n640) );
  XNOR2_X1 U720 ( .A(n640), .B(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G61), .A2(n654), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G48), .A2(n661), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n655), .A2(G86), .ZN(n643) );
  XOR2_X1 U725 ( .A(KEYINPUT84), .B(n643), .Z(n644) );
  NOR2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U728 ( .A1(G49), .A2(n661), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U731 ( .A1(n654), .A2(n650), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n651), .A2(G87), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(G288) );
  AND2_X1 U734 ( .A1(n654), .A2(G60), .ZN(n660) );
  NAND2_X1 U735 ( .A1(G85), .A2(n655), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G72), .A2(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n661), .A2(G47), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(G290) );
  INV_X1 U741 ( .A(G299), .ZN(n988) );
  XNOR2_X1 U742 ( .A(KEYINPUT87), .B(G305), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(G288), .ZN(n665) );
  XNOR2_X1 U744 ( .A(KEYINPUT19), .B(n665), .ZN(n667) );
  XNOR2_X1 U745 ( .A(G290), .B(n673), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U747 ( .A(G166), .B(n668), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n988), .B(n669), .ZN(n920) );
  XOR2_X1 U749 ( .A(n920), .B(n670), .Z(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G868), .ZN(n672) );
  XOR2_X1 U751 ( .A(KEYINPUT88), .B(n672), .Z(n675) );
  NOR2_X1 U752 ( .A1(n673), .A2(G868), .ZN(n674) );
  NOR2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U754 ( .A(KEYINPUT89), .B(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n677) );
  XNOR2_X1 U757 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U764 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G96), .A2(n684), .ZN(n856) );
  NAND2_X1 U766 ( .A1(G2106), .A2(n856), .ZN(n685) );
  XNOR2_X1 U767 ( .A(n685), .B(KEYINPUT91), .ZN(n691) );
  NOR2_X1 U768 ( .A1(G235), .A2(G236), .ZN(n686) );
  XNOR2_X1 U769 ( .A(KEYINPUT92), .B(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n687), .A2(G57), .ZN(n688) );
  NOR2_X1 U771 ( .A1(G238), .A2(n688), .ZN(n858) );
  NOR2_X1 U772 ( .A1(n689), .A2(n858), .ZN(n690) );
  NOR2_X1 U773 ( .A1(n691), .A2(n690), .ZN(G319) );
  INV_X1 U774 ( .A(G319), .ZN(n693) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U776 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U777 ( .A(KEYINPUT93), .B(n694), .Z(n855) );
  NAND2_X1 U778 ( .A1(G36), .A2(n855), .ZN(n695) );
  XNOR2_X1 U779 ( .A(n695), .B(KEYINPUT94), .ZN(G176) );
  XNOR2_X1 U780 ( .A(G1986), .B(G290), .ZN(n998) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n727) );
  NAND2_X1 U782 ( .A1(G160), .A2(G40), .ZN(n696) );
  NOR2_X1 U783 ( .A1(n727), .A2(n696), .ZN(n837) );
  NAND2_X1 U784 ( .A1(n998), .A2(n837), .ZN(n825) );
  XNOR2_X1 U785 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  NAND2_X1 U786 ( .A1(n903), .A2(G104), .ZN(n697) );
  XOR2_X1 U787 ( .A(KEYINPUT95), .B(n697), .Z(n699) );
  NAND2_X1 U788 ( .A1(n900), .A2(G140), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U790 ( .A(KEYINPUT34), .B(n700), .ZN(n706) );
  NAND2_X1 U791 ( .A1(G116), .A2(n895), .ZN(n702) );
  NAND2_X1 U792 ( .A1(G128), .A2(n896), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U794 ( .A(KEYINPUT35), .B(n703), .Z(n704) );
  XNOR2_X1 U795 ( .A(KEYINPUT96), .B(n704), .ZN(n705) );
  NOR2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U797 ( .A(KEYINPUT36), .B(n707), .ZN(n916) );
  OR2_X1 U798 ( .A1(n835), .A2(n916), .ZN(n708) );
  XNOR2_X1 U799 ( .A(KEYINPUT97), .B(n708), .ZN(n947) );
  NAND2_X1 U800 ( .A1(n837), .A2(n947), .ZN(n833) );
  NAND2_X1 U801 ( .A1(G141), .A2(n900), .ZN(n710) );
  NAND2_X1 U802 ( .A1(G117), .A2(n895), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n903), .A2(G105), .ZN(n711) );
  XOR2_X1 U805 ( .A(KEYINPUT38), .B(n711), .Z(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n896), .A2(G129), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n893) );
  NAND2_X1 U809 ( .A1(G1996), .A2(n893), .ZN(n723) );
  NAND2_X1 U810 ( .A1(G131), .A2(n900), .ZN(n717) );
  NAND2_X1 U811 ( .A1(G107), .A2(n895), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U813 ( .A1(G95), .A2(n903), .ZN(n719) );
  NAND2_X1 U814 ( .A1(G119), .A2(n896), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n720) );
  OR2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n913) );
  NAND2_X1 U817 ( .A1(G1991), .A2(n913), .ZN(n722) );
  NAND2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U819 ( .A(KEYINPUT98), .B(n724), .Z(n936) );
  INV_X1 U820 ( .A(n936), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n837), .A2(n725), .ZN(n826) );
  NAND2_X1 U822 ( .A1(n833), .A2(n826), .ZN(n726) );
  XOR2_X1 U823 ( .A(KEYINPUT99), .B(n726), .Z(n823) );
  AND2_X1 U824 ( .A1(n727), .A2(G40), .ZN(n728) );
  NAND2_X1 U825 ( .A1(n728), .A2(G160), .ZN(n729) );
  XNOR2_X2 U826 ( .A(n729), .B(KEYINPUT64), .ZN(n776) );
  NAND2_X1 U827 ( .A1(n776), .A2(G8), .ZN(n816) );
  NOR2_X1 U828 ( .A1(G1981), .A2(G305), .ZN(n730) );
  XOR2_X1 U829 ( .A(n730), .B(KEYINPUT24), .Z(n731) );
  NOR2_X1 U830 ( .A1(n816), .A2(n731), .ZN(n821) );
  INV_X1 U831 ( .A(n776), .ZN(n761) );
  NAND2_X1 U832 ( .A1(G2072), .A2(n761), .ZN(n733) );
  XOR2_X1 U833 ( .A(KEYINPUT101), .B(KEYINPUT27), .Z(n732) );
  XNOR2_X1 U834 ( .A(n733), .B(n732), .ZN(n735) );
  INV_X1 U835 ( .A(G1956), .ZN(n1010) );
  NOR2_X1 U836 ( .A1(n761), .A2(n1010), .ZN(n734) );
  NOR2_X1 U837 ( .A1(n735), .A2(n734), .ZN(n738) );
  NOR2_X1 U838 ( .A1(n738), .A2(n988), .ZN(n737) );
  XNOR2_X1 U839 ( .A(n737), .B(n736), .ZN(n757) );
  NAND2_X1 U840 ( .A1(n738), .A2(n988), .ZN(n755) );
  XNOR2_X1 U841 ( .A(KEYINPUT26), .B(KEYINPUT102), .ZN(n745) );
  NOR2_X1 U842 ( .A1(G1996), .A2(n745), .ZN(n739) );
  NOR2_X1 U843 ( .A1(n1002), .A2(n739), .ZN(n743) );
  NAND2_X1 U844 ( .A1(G2067), .A2(n761), .ZN(n741) );
  NAND2_X1 U845 ( .A1(n776), .A2(G1348), .ZN(n740) );
  NAND2_X1 U846 ( .A1(n741), .A2(n740), .ZN(n751) );
  NAND2_X1 U847 ( .A1(n985), .A2(n751), .ZN(n742) );
  NAND2_X1 U848 ( .A1(n743), .A2(n742), .ZN(n750) );
  INV_X1 U849 ( .A(G1341), .ZN(n1011) );
  NAND2_X1 U850 ( .A1(n1011), .A2(n745), .ZN(n744) );
  NAND2_X1 U851 ( .A1(n744), .A2(n776), .ZN(n748) );
  AND2_X1 U852 ( .A1(n761), .A2(G1996), .ZN(n746) );
  NAND2_X1 U853 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U854 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U855 ( .A1(n750), .A2(n749), .ZN(n753) );
  NOR2_X1 U856 ( .A1(n751), .A2(n985), .ZN(n752) );
  NOR2_X1 U857 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U858 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U859 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U860 ( .A(n758), .B(KEYINPUT29), .ZN(n759) );
  XNOR2_X1 U861 ( .A(n759), .B(KEYINPUT103), .ZN(n765) );
  XOR2_X1 U862 ( .A(G2078), .B(KEYINPUT25), .Z(n962) );
  NOR2_X1 U863 ( .A1(n776), .A2(n962), .ZN(n760) );
  XNOR2_X1 U864 ( .A(n760), .B(KEYINPUT100), .ZN(n763) );
  NOR2_X1 U865 ( .A1(n761), .A2(G1961), .ZN(n762) );
  NOR2_X1 U866 ( .A1(n763), .A2(n762), .ZN(n771) );
  OR2_X1 U867 ( .A1(G301), .A2(n771), .ZN(n764) );
  NAND2_X1 U868 ( .A1(n765), .A2(n764), .ZN(n787) );
  INV_X1 U869 ( .A(G168), .ZN(n770) );
  NOR2_X1 U870 ( .A1(G1966), .A2(n816), .ZN(n789) );
  NOR2_X1 U871 ( .A1(n776), .A2(G2084), .ZN(n788) );
  NOR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n766) );
  NAND2_X1 U873 ( .A1(G8), .A2(n766), .ZN(n767) );
  XNOR2_X1 U874 ( .A(KEYINPUT104), .B(n767), .ZN(n768) );
  XOR2_X1 U875 ( .A(KEYINPUT30), .B(n768), .Z(n769) );
  NAND2_X1 U876 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U877 ( .A1(n771), .A2(G301), .ZN(n772) );
  NAND2_X1 U878 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U879 ( .A(n774), .B(KEYINPUT31), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n775) );
  NAND2_X1 U881 ( .A1(n775), .A2(G286), .ZN(n784) );
  INV_X1 U882 ( .A(G8), .ZN(n782) );
  NOR2_X1 U883 ( .A1(n776), .A2(G2090), .ZN(n778) );
  NOR2_X1 U884 ( .A1(G1971), .A2(n816), .ZN(n777) );
  NOR2_X1 U885 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U886 ( .A(KEYINPUT105), .B(n779), .Z(n780) );
  NAND2_X1 U887 ( .A1(n780), .A2(G303), .ZN(n781) );
  OR2_X1 U888 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U889 ( .A1(n787), .A2(n786), .ZN(n792) );
  AND2_X1 U890 ( .A1(G8), .A2(n788), .ZN(n790) );
  OR2_X1 U891 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U892 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U893 ( .A(KEYINPUT33), .ZN(n793) );
  NAND2_X1 U894 ( .A1(n992), .A2(n793), .ZN(n799) );
  INV_X1 U895 ( .A(n799), .ZN(n794) );
  AND2_X1 U896 ( .A1(n813), .A2(n794), .ZN(n795) );
  NAND2_X1 U897 ( .A1(n812), .A2(n795), .ZN(n801) );
  NOR2_X1 U898 ( .A1(G1976), .A2(G288), .ZN(n991) );
  NOR2_X1 U899 ( .A1(G1971), .A2(G303), .ZN(n796) );
  XNOR2_X1 U900 ( .A(KEYINPUT106), .B(n796), .ZN(n797) );
  NOR2_X1 U901 ( .A1(n991), .A2(n797), .ZN(n798) );
  OR2_X1 U902 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U903 ( .A1(n801), .A2(n800), .ZN(n802) );
  INV_X1 U904 ( .A(n816), .ZN(n803) );
  NAND2_X1 U905 ( .A1(n802), .A2(n803), .ZN(n806) );
  NAND2_X1 U906 ( .A1(n991), .A2(n803), .ZN(n804) );
  NAND2_X1 U907 ( .A1(n804), .A2(KEYINPUT33), .ZN(n805) );
  NAND2_X1 U908 ( .A1(n806), .A2(n805), .ZN(n808) );
  XNOR2_X1 U909 ( .A(n808), .B(n807), .ZN(n809) );
  XOR2_X1 U910 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U911 ( .A1(n809), .A2(n982), .ZN(n819) );
  NOR2_X1 U912 ( .A1(G2090), .A2(G303), .ZN(n810) );
  XNOR2_X1 U913 ( .A(n810), .B(KEYINPUT108), .ZN(n811) );
  NAND2_X1 U914 ( .A1(n811), .A2(G8), .ZN(n815) );
  NAND2_X1 U915 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U916 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U917 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n840) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n893), .ZN(n934) );
  INV_X1 U923 ( .A(n826), .ZN(n830) );
  NOR2_X1 U924 ( .A1(G1991), .A2(n913), .ZN(n939) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n827) );
  XOR2_X1 U926 ( .A(n827), .B(KEYINPUT109), .Z(n828) );
  NOR2_X1 U927 ( .A1(n939), .A2(n828), .ZN(n829) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U929 ( .A1(n934), .A2(n831), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n832), .B(KEYINPUT39), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n835), .A2(n916), .ZN(n944) );
  NAND2_X1 U933 ( .A1(n836), .A2(n944), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U937 ( .A(G2454), .B(G2451), .ZN(n850) );
  XNOR2_X1 U938 ( .A(G2430), .B(G2446), .ZN(n848) );
  XOR2_X1 U939 ( .A(G2435), .B(G2427), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT110), .B(G2438), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(n844), .B(G2443), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1341), .B(G1348), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U947 ( .A1(n851), .A2(G14), .ZN(n926) );
  XNOR2_X1 U948 ( .A(KEYINPUT111), .B(n926), .ZN(G401) );
  INV_X1 U949 ( .A(G223), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G2106), .A2(n852), .ZN(G217) );
  AND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G661), .A2(n853), .ZN(G259) );
  NAND2_X1 U953 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(G188) );
  INV_X1 U956 ( .A(G96), .ZN(G221) );
  INV_X1 U957 ( .A(G57), .ZN(G237) );
  INV_X1 U958 ( .A(n856), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(G261) );
  INV_X1 U960 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U961 ( .A(G1966), .B(KEYINPUT41), .ZN(n868) );
  XOR2_X1 U962 ( .A(G1981), .B(G1961), .Z(n860) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1956), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U965 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U967 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U968 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT112), .B(G2474), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(G229) );
  XOR2_X1 U972 ( .A(G2100), .B(G2096), .Z(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT42), .B(G2678), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U975 ( .A(KEYINPUT43), .B(G2090), .Z(n872) );
  XNOR2_X1 U976 ( .A(G2067), .B(G2072), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U978 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U979 ( .A(G2078), .B(G2084), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(G227) );
  NAND2_X1 U981 ( .A1(G124), .A2(n896), .ZN(n877) );
  XOR2_X1 U982 ( .A(KEYINPUT113), .B(n877), .Z(n878) );
  XNOR2_X1 U983 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G112), .A2(n895), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G136), .A2(n900), .ZN(n882) );
  NAND2_X1 U987 ( .A1(G100), .A2(n903), .ZN(n881) );
  NAND2_X1 U988 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U989 ( .A1(n884), .A2(n883), .ZN(G162) );
  NAND2_X1 U990 ( .A1(G118), .A2(n895), .ZN(n886) );
  NAND2_X1 U991 ( .A1(G130), .A2(n896), .ZN(n885) );
  NAND2_X1 U992 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U993 ( .A(KEYINPUT114), .B(n887), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G142), .A2(n900), .ZN(n889) );
  NAND2_X1 U995 ( .A1(G106), .A2(n903), .ZN(n888) );
  NAND2_X1 U996 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U997 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U998 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U999 ( .A(n894), .B(n893), .ZN(n910) );
  XOR2_X1 U1000 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n908) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n895), .ZN(n898) );
  NAND2_X1 U1002 ( .A1(G127), .A2(n896), .ZN(n897) );
  NAND2_X1 U1003 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U1004 ( .A(n899), .B(KEYINPUT47), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n900), .ZN(n901) );
  NAND2_X1 U1006 ( .A1(n902), .A2(n901), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n903), .ZN(n904) );
  XNOR2_X1 U1008 ( .A(KEYINPUT115), .B(n904), .ZN(n905) );
  NOR2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n949) );
  XNOR2_X1 U1010 ( .A(n949), .B(KEYINPUT116), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1012 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1013 ( .A(G164), .B(G162), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(n912), .B(n911), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(G160), .B(n913), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(n914), .B(n940), .ZN(n915) );
  XOR2_X1 U1017 ( .A(n916), .B(n915), .Z(n917) );
  XNOR2_X1 U1018 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n919), .ZN(G395) );
  XNOR2_X1 U1020 ( .A(G286), .B(n920), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n921), .B(G171), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(n1002), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(G37), .A2(n925), .ZN(G397) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n926), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1032 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1042) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n956) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G162), .ZN(n932) );
  XNOR2_X1 U1035 ( .A(n932), .B(KEYINPUT117), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n935), .Z(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n943) );
  XOR2_X1 U1039 ( .A(G160), .B(G2084), .Z(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT118), .B(n948), .ZN(n954) );
  XOR2_X1 U1046 ( .A(G2072), .B(n949), .Z(n951) );
  XOR2_X1 U1047 ( .A(G164), .B(G2078), .Z(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(KEYINPUT50), .B(n952), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n956), .B(n955), .ZN(n957) );
  INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n978) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n978), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(G29), .ZN(n1040) );
  XOR2_X1 U1055 ( .A(G2067), .B(G26), .Z(n959) );
  NAND2_X1 U1056 ( .A1(n959), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G1996), .B(G32), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G1991), .B(G25), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(G27), .B(n962), .ZN(n963) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1065 ( .A(n969), .B(KEYINPUT53), .Z(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT121), .B(n970), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT54), .B(G2084), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G34), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1070 ( .A(G2090), .B(KEYINPUT120), .Z(n974) );
  XNOR2_X1 U1071 ( .A(G35), .B(n974), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(n978), .B(n977), .ZN(n980) );
  INV_X1 U1074 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n981), .ZN(n1038) );
  XNOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(KEYINPUT57), .B(n984), .ZN(n1006) );
  XNOR2_X1 U1081 ( .A(n985), .B(G1348), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(G301), .B(G1961), .ZN(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G166), .B(G1971), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(n988), .B(G1956), .ZN(n989) );
  NAND2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n995) );
  XOR2_X1 U1087 ( .A(n991), .B(KEYINPUT122), .Z(n993) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(KEYINPUT123), .B(n996), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT124), .B(n1001), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(n1011), .B(n1002), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1036) );
  INV_X1 U1098 ( .A(G16), .ZN(n1034) );
  XNOR2_X1 U1099 ( .A(KEYINPUT125), .B(G1961), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(G5), .ZN(n1029) );
  XNOR2_X1 U1101 ( .A(n1010), .B(G20), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(n1011), .B(G19), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(G1981), .B(G6), .Z(n1012) );
  XNOR2_X1 U1104 ( .A(KEYINPUT126), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1107 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1110 ( .A(n1020), .B(KEYINPUT60), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1114 ( .A(G1986), .B(G24), .Z(n1023) );
  NAND2_X1 U1115 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1116 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(G21), .B(G1966), .ZN(n1030) );
  NOR2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1126 ( .A(n1042), .B(n1041), .ZN(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

