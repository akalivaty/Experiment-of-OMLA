//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT67), .B(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G120gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n202), .B(new_n204), .C1(new_n207), .C2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G113gat), .B(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n203), .B1(KEYINPUT1), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n217), .B(new_n220), .C1(new_n221), .C2(KEYINPUT2), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G148gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G141gat), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT79), .B(G148gat), .Z(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G141gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n222), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n229), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT80), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n216), .ZN(new_n234));
  INV_X1    g033(.A(new_n229), .ZN(new_n235));
  OR3_X1    g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT80), .ZN(new_n236));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n230), .B(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n216), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n237), .ZN(new_n247));
  OAI211_X1 g046(.A(KEYINPUT5), .B(new_n239), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT82), .B(G1gat), .Z(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G57gat), .B(G85gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G29gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n251), .B(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n241), .A2(new_n245), .A3(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n248), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n254), .B1(new_n248), .B2(new_n256), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT6), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n260));
  AOI211_X1 g059(.A(new_n260), .B(new_n254), .C1(new_n248), .C2(new_n256), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT71), .B(G211gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT72), .B(G218gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT22), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n267), .A2(new_n268), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n264), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n265), .A2(new_n266), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT73), .B1(new_n278), .B2(KEYINPUT22), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n267), .A2(new_n268), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n274), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n285), .ZN(new_n292));
  OR3_X1    g091(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n289), .A2(new_n292), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  INV_X1    g099(.A(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n304), .A3(new_n294), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n297), .A2(KEYINPUT24), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT65), .A4(new_n294), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(G183gat), .A3(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n297), .A2(KEYINPUT24), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n320), .A2(new_n305), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n299), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n284), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n315), .B2(new_n316), .ZN(new_n326));
  OAI211_X1 g125(.A(G226gat), .B(G233gat), .C1(new_n326), .C2(new_n299), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT75), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n326), .B2(new_n299), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n284), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n283), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n283), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n325), .A3(new_n327), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT77), .Z(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n335), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n341), .B1(new_n333), .B2(new_n335), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n345), .A2(KEYINPUT30), .ZN(new_n346));
  INV_X1    g145(.A(new_n341), .ZN(new_n347));
  AND4_X1   g146(.A1(KEYINPUT78), .A2(new_n336), .A3(KEYINPUT30), .A4(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT78), .B1(new_n345), .B2(KEYINPUT30), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n344), .B(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT85), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n345), .A2(KEYINPUT30), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n335), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n333), .B2(new_n335), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n356), .B2(new_n342), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n336), .A2(KEYINPUT30), .A3(new_n347), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT78), .A3(KEYINPUT30), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n352), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n263), .B1(new_n351), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G22gat), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n276), .B2(new_n282), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n229), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n372));
  INV_X1    g171(.A(G228gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n243), .A2(new_n330), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n334), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n372), .A2(new_n377), .A3(KEYINPUT84), .A4(new_n375), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n330), .B1(new_n281), .B2(new_n273), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n273), .B(new_n264), .C1(new_n269), .C2(new_n270), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n242), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n229), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n375), .B1(new_n387), .B2(new_n377), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n370), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  AOI211_X1 g189(.A(G22gat), .B(new_n388), .C1(new_n380), .C2(new_n381), .ZN(new_n391));
  OAI211_X1 g190(.A(KEYINPUT83), .B(new_n369), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n324), .A2(new_n216), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n234), .B1(new_n326), .B2(new_n299), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n393), .A2(new_n394), .B1(G227gat), .B2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(KEYINPUT68), .A3(KEYINPUT34), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT34), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n399), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT69), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT69), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n395), .A2(new_n404), .A3(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G15gat), .B(G43gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G71gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G99gat), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n393), .A2(G227gat), .A3(G233gat), .A4(new_n394), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(KEYINPUT32), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n411), .B(KEYINPUT32), .C1(new_n412), .C2(new_n410), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n401), .A2(new_n406), .A3(new_n415), .A4(new_n416), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT89), .B1(new_n418), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT83), .B1(new_n390), .B2(new_n391), .ZN(new_n423));
  INV_X1    g222(.A(new_n369), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n392), .A2(new_n422), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n350), .A2(KEYINPUT85), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n362), .A2(new_n352), .A3(new_n344), .A4(new_n346), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(KEYINPUT88), .A3(new_n263), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n366), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n417), .A3(KEYINPUT70), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n419), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(KEYINPUT70), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n425), .A2(new_n392), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n262), .A2(new_n350), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT35), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n433), .B(KEYINPUT36), .C1(new_n434), .C2(KEYINPUT70), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(KEYINPUT36), .B2(new_n434), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n392), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n233), .A2(new_n236), .ZN(new_n444));
  OR3_X1    g243(.A1(new_n444), .A2(KEYINPUT86), .A3(new_n238), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n246), .A2(new_n238), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT86), .B1(new_n444), .B2(new_n238), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(KEYINPUT39), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(KEYINPUT39), .ZN(new_n449));
  INV_X1    g248(.A(new_n254), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(KEYINPUT87), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(new_n258), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(KEYINPUT87), .A3(new_n453), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n428), .A3(new_n429), .A4(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n442), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n347), .B1(new_n356), .B2(KEYINPUT37), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n336), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(KEYINPUT38), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n325), .A2(new_n327), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n283), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n328), .A2(new_n332), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT37), .B(new_n464), .C1(new_n465), .C2(new_n283), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n466), .A3(new_n342), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  INV_X1    g267(.A(new_n345), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n262), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n458), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n432), .A2(new_n439), .B1(new_n443), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(G1gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(G1gat), .B2(new_n475), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G8gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(KEYINPUT92), .A3(G8gat), .ZN(new_n482));
  AOI21_X1  g281(.A(G8gat), .B1(new_n478), .B2(KEYINPUT93), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(G43gat), .B(G50gat), .Z(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR3_X1    g288(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n490), .A2(new_n491), .B1(G29gat), .B2(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n487), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n493), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT17), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(KEYINPUT15), .A3(new_n494), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n489), .A2(new_n495), .A3(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n478), .A2(KEYINPUT93), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n485), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT92), .B1(new_n478), .B2(G8gat), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n478), .A2(KEYINPUT92), .A3(G8gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n500), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT94), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n503), .A2(new_n510), .A3(KEYINPUT18), .A4(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT96), .B1(new_n486), .B2(new_n496), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n509), .A2(new_n517), .A3(new_n500), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT97), .B1(new_n509), .B2(new_n500), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n486), .A2(new_n521), .A3(new_n496), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n512), .B(KEYINPUT13), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n515), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n510), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(new_n512), .ZN(new_n530));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT12), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n527), .B(new_n530), .C1(KEYINPUT95), .C2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n516), .A2(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n530), .B(new_n514), .C1(new_n539), .C2(new_n525), .ZN(new_n540));
  OAI211_X1 g339(.A(KEYINPUT95), .B(new_n514), .C1(new_n539), .C2(new_n525), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G183gat), .B(G211gat), .ZN(new_n545));
  INV_X1    g344(.A(G127gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n218), .ZN(new_n548));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT98), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G57gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G64gat), .ZN(new_n560));
  INV_X1    g359(.A(G64gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G57gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n555), .B(new_n558), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n562), .A2(KEYINPUT100), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n562), .A2(KEYINPUT100), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT101), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n573), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n486), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT103), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT103), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n567), .B1(new_n564), .B2(new_n565), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n582), .A2(new_n554), .A3(new_n557), .ZN(new_n583));
  INV_X1    g382(.A(new_n576), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n581), .B1(new_n586), .B2(new_n486), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n553), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(KEYINPUT103), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n581), .A3(new_n486), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n552), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n577), .A2(new_n578), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT102), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n588), .B2(new_n591), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n551), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT7), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(G85gat), .A3(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n599), .A2(new_n601), .B1(KEYINPUT8), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT104), .B(G92gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(G85gat), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n497), .A2(new_n502), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n605), .B(new_n606), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n500), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT105), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n614), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(KEYINPUT105), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n615), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n615), .A2(new_n618), .ZN(new_n624));
  INV_X1    g423(.A(new_n621), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n617), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n588), .A2(new_n591), .ZN(new_n627));
  INV_X1    g426(.A(new_n593), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n550), .A3(new_n594), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n597), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n597), .A2(new_n626), .A3(new_n630), .A4(KEYINPUT106), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n610), .A2(new_n568), .A3(new_n576), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n607), .B1(new_n583), .B2(new_n584), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT107), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n635), .A2(new_n636), .A3(new_n641), .A4(new_n637), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT108), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n635), .A2(new_n636), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(G230gat), .A3(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n643), .A2(new_n644), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n648), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n633), .A2(new_n634), .A3(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n474), .A2(new_n544), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n262), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NOR4_X1   g460(.A1(new_n474), .A2(new_n544), .A3(new_n430), .A4(new_n658), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n476), .A2(new_n505), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n476), .A2(new_n505), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n662), .A2(new_n505), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n662), .A2(KEYINPUT42), .A3(new_n664), .A4(new_n665), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT109), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n668), .A2(new_n673), .A3(new_n669), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1325gat));
  AOI21_X1  g474(.A(G15gat), .B1(new_n659), .B2(new_n422), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT110), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n441), .A2(G15gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n659), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n659), .A2(new_n442), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n432), .A2(new_n439), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n473), .A2(new_n443), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n626), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n597), .A2(new_n630), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n653), .A2(new_n656), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n685), .A2(new_n543), .A3(new_n686), .A4(new_n690), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n691), .A2(G29gat), .A3(new_n263), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n474), .B2(new_n626), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT35), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n425), .A2(new_n392), .A3(new_n435), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n437), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT88), .B1(new_n430), .B2(new_n263), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n365), .B(new_n262), .C1(new_n428), .C2(new_n429), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n698), .B1(new_n701), .B2(new_n427), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n473), .A2(new_n443), .ZN(new_n703));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n686), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n538), .A2(KEYINPUT111), .A3(new_n542), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT111), .B1(new_n538), .B2(new_n542), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n695), .A2(new_n704), .A3(new_n707), .A4(new_n690), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n263), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n709), .ZN(G1328gat));
  OR3_X1    g509(.A1(new_n691), .A2(G36gat), .A3(new_n430), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n708), .B2(new_n430), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n422), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n691), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n441), .A2(G43gat), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n718), .B(new_n720), .C1(new_n708), .C2(new_n721), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n719), .A2(KEYINPUT47), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n708), .B2(new_n458), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n691), .A2(G50gat), .A3(new_n458), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  AOI21_X1  g529(.A(new_n657), .B1(new_n683), .B2(new_n684), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n633), .B(new_n634), .C1(new_n705), .C2(new_n706), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n263), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n559), .ZN(G1332gat));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n731), .B2(new_n733), .ZN(new_n738));
  NOR4_X1   g537(.A1(new_n474), .A2(KEYINPUT113), .A3(new_n657), .A4(new_n732), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n430), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n740), .A2(new_n741), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n441), .B1(new_n738), .B2(new_n739), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G71gat), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n717), .A2(G71gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n747), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(KEYINPUT50), .B(new_n751), .C1(new_n748), .C2(G71gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n442), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g556(.A1(new_n705), .A2(new_n706), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(KEYINPUT114), .A3(new_n687), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n707), .B2(new_n688), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n689), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT115), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n695), .A2(new_n704), .A3(new_n262), .A4(new_n764), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(G85gat), .A3(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n686), .B(new_n762), .C1(new_n702), .C2(new_n703), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT51), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n685), .A2(new_n771), .A3(new_n686), .A4(new_n762), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n263), .A2(G85gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n770), .A2(new_n689), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n774), .ZN(G1336gat));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n430), .A2(G92gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n770), .A2(new_n689), .A3(new_n772), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(KEYINPUT117), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n695), .A2(new_n704), .A3(new_n764), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n604), .B1(new_n780), .B2(new_n430), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n778), .C1(KEYINPUT117), .C2(new_n776), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1337gat));
  NAND4_X1  g584(.A1(new_n695), .A2(new_n704), .A3(new_n441), .A4(new_n764), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G99gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n717), .A2(G99gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n689), .A3(new_n772), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1338gat));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n695), .A2(new_n704), .A3(new_n442), .A4(new_n764), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n458), .A2(G106gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n770), .A2(new_n689), .A3(new_n772), .A4(new_n794), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n791), .B(KEYINPUT53), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n798));
  AND4_X1   g597(.A1(new_n797), .A2(new_n793), .A3(new_n798), .A4(new_n795), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(G1339gat));
  NOR2_X1   g599(.A1(new_n732), .A2(new_n689), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  INV_X1    g601(.A(new_n645), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n639), .A2(new_n803), .A3(new_n640), .A4(new_n642), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n643), .A2(new_n806), .A3(new_n645), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n652), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n652), .A4(new_n807), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n809), .A2(new_n811), .A3(new_n656), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n540), .A2(new_n536), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n539), .A2(new_n525), .B1(new_n512), .B2(new_n529), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n535), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(new_n686), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n689), .A2(new_n816), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n812), .B2(new_n707), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(new_n686), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n801), .B1(new_n821), .B2(new_n687), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n442), .A3(new_n717), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n741), .A2(new_n263), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT119), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n544), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n822), .A2(new_n263), .A3(new_n741), .A4(new_n436), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n758), .A2(new_n205), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT120), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n826), .B2(new_n657), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n206), .A3(new_n689), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1341gat));
  NOR3_X1   g634(.A1(new_n826), .A2(new_n546), .A3(new_n687), .ZN(new_n836));
  AOI21_X1  g635(.A(G127gat), .B1(new_n828), .B2(new_n688), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n826), .B2(new_n626), .ZN(new_n839));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n828), .A2(new_n840), .A3(new_n686), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT56), .Z(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(G1343gat));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n809), .A2(new_n543), .A3(new_n656), .A4(new_n811), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n818), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n626), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n817), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n687), .ZN(new_n849));
  INV_X1    g648(.A(new_n801), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n844), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(KEYINPUT121), .A3(new_n442), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n844), .B1(new_n822), .B2(new_n458), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n688), .B1(new_n847), .B2(new_n817), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n801), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n856), .B2(new_n458), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n441), .A2(new_n263), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n430), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n543), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT58), .B1(new_n862), .B2(G141gat), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n821), .A2(new_n687), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n442), .B(new_n859), .C1(new_n864), .C2(new_n801), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n822), .A2(new_n458), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT122), .A3(new_n859), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n867), .A2(new_n430), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n544), .A2(G141gat), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n707), .A3(new_n861), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n822), .A2(new_n458), .A3(new_n860), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n875), .A2(G141gat), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n873), .B1(new_n874), .B2(new_n877), .ZN(G1344gat));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n822), .B2(new_n458), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n658), .A2(new_n543), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n844), .B(new_n442), .C1(new_n855), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n689), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G148gat), .B1(new_n882), .B2(new_n860), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT59), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n858), .A2(new_n689), .A3(new_n861), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n887), .B2(new_n227), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n867), .A2(new_n869), .A3(new_n227), .A4(new_n430), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n657), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(KEYINPUT123), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n889), .A2(new_n892), .A3(new_n657), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n891), .B2(new_n893), .ZN(G1345gat));
  AOI21_X1  g693(.A(G155gat), .B1(new_n870), .B2(new_n688), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n858), .A2(new_n861), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n687), .A2(new_n218), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n870), .B2(new_n686), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n626), .A2(new_n219), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n896), .B2(new_n900), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n741), .A2(new_n263), .ZN(new_n902));
  NOR4_X1   g701(.A1(new_n822), .A2(new_n442), .A3(new_n717), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n300), .B1(new_n903), .B2(new_n543), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT125), .Z(new_n905));
  NAND2_X1  g704(.A1(new_n697), .A2(new_n741), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n908));
  NOR4_X1   g707(.A1(new_n822), .A2(new_n907), .A3(new_n908), .A4(new_n262), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n300), .A3(new_n707), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n910), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n909), .B2(new_n689), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n657), .A2(new_n301), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n903), .B2(new_n913), .ZN(G1349gat));
  NAND2_X1  g713(.A1(new_n903), .A2(new_n688), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G183gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n909), .A2(new_n290), .A3(new_n688), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g718(.A(new_n285), .B1(new_n903), .B2(new_n686), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT61), .Z(new_n921));
  NAND3_X1  g720(.A1(new_n909), .A2(new_n285), .A3(new_n686), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1351gat));
  NOR4_X1   g722(.A1(new_n822), .A2(new_n458), .A3(new_n441), .A4(new_n902), .ZN(new_n924));
  INV_X1    g723(.A(G197gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n707), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n902), .A2(KEYINPUT126), .A3(new_n441), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n902), .B2(new_n441), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n879), .A2(new_n881), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(new_n543), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n931), .B2(new_n925), .ZN(G1352gat));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n924), .A2(new_n933), .A3(new_n689), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n882), .B1(new_n927), .B2(new_n928), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n936), .B(new_n937), .C1(new_n933), .C2(new_n938), .ZN(G1353gat));
  INV_X1    g738(.A(new_n265), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n940), .A3(new_n688), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n879), .A2(new_n688), .A3(new_n881), .A4(new_n929), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n941), .B(KEYINPUT127), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n924), .B2(new_n686), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n686), .A2(new_n266), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n930), .B2(new_n951), .ZN(G1355gat));
endmodule


