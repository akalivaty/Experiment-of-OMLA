//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  XNOR2_X1  g0004(.A(KEYINPUT66), .B(G244), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n204), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n204), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT65), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n224), .B1(G58), .B2(G68), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n225), .A3(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n214), .B(new_n217), .C1(new_n220), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G294), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT81), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT81), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n251), .A3(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT80), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(new_n248), .B2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(new_n263), .B2(G250), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n247), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n255), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT94), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT94), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n271), .A3(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n273), .A2(new_n274), .A3(G1), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT86), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(new_n266), .A3(KEYINPUT5), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT5), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(KEYINPUT86), .B2(G41), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n275), .A2(new_n267), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n273), .A2(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n282), .A2(G264), .A3(new_n267), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n270), .A2(new_n272), .A3(new_n280), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G169), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n287), .B(new_n283), .C1(new_n265), .C2(new_n268), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n280), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n218), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n248), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT70), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n248), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT22), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n301), .A2(new_n302), .A3(new_n219), .A4(G87), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n252), .A2(new_n219), .A3(new_n254), .A4(new_n256), .ZN(new_n305));
  INV_X1    g0105(.A(G87), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT22), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT93), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n254), .A2(new_n256), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n310), .A2(new_n219), .A3(G87), .A4(new_n252), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT93), .A3(KEYINPUT22), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n304), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G107), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT23), .B1(new_n314), .B2(G20), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(KEYINPUT23), .A3(G20), .ZN(new_n317));
  INV_X1    g0117(.A(G116), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n255), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n316), .A2(new_n317), .B1(new_n319), .B2(new_n219), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT24), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n311), .A2(KEYINPUT93), .A3(KEYINPUT22), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT93), .B1(new_n311), .B2(KEYINPUT22), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n303), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT24), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n320), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n293), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G13), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n329), .A2(new_n219), .A3(G1), .ZN(new_n330));
  INV_X1    g0130(.A(G1), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n292), .B(new_n330), .C1(new_n331), .C2(G33), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT25), .B1(new_n330), .B2(new_n314), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(KEYINPUT25), .A3(new_n314), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n332), .A2(G107), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n290), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n313), .A2(KEYINPUT24), .A3(new_n321), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n326), .B1(new_n325), .B2(new_n320), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n292), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n247), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n249), .A2(new_n251), .A3(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n254), .A2(new_n256), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G250), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(new_n258), .B2(new_n259), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n342), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n280), .B(new_n284), .C1(new_n351), .C2(new_n267), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n285), .B2(G190), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n341), .A2(new_n336), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n338), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT8), .B(G58), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n255), .A2(G20), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n359), .A2(new_n221), .A3(KEYINPUT8), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G50), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n221), .A3(new_n222), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G20), .A2(G33), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(G20), .B1(G150), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n293), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n330), .A2(new_n364), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n292), .B1(new_n331), .B2(G20), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(new_n364), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT9), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OR3_X1    g0175(.A1(new_n368), .A2(new_n372), .A3(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT69), .B(G45), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n331), .B(G274), .C1(new_n379), .C2(G41), .ZN(new_n380));
  INV_X1    g0180(.A(G226), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n331), .B1(G41), .B2(G45), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n267), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n259), .B1(new_n296), .B2(new_n300), .ZN(new_n385));
  INV_X1    g0185(.A(new_n300), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n299), .B1(new_n297), .B2(new_n298), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n385), .A2(G223), .B1(new_n388), .B2(G77), .ZN(new_n389));
  INV_X1    g0189(.A(G222), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n301), .A2(new_n263), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n384), .B1(new_n392), .B2(new_n268), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G190), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n378), .B(new_n394), .C1(new_n353), .C2(new_n393), .ZN(new_n395));
  XOR2_X1   g0195(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT75), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(KEYINPUT10), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(new_n268), .ZN(new_n399));
  INV_X1    g0199(.A(new_n384), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n377), .B1(new_n401), .B2(G200), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  INV_X1    g0203(.A(new_n396), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n394), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n398), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n401), .A2(G179), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n373), .B1(new_n393), .B2(G169), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n361), .A2(G77), .ZN(new_n412));
  INV_X1    g0212(.A(new_n366), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n412), .B1(new_n219), .B2(G68), .C1(new_n364), .C2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(new_n292), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n330), .A2(new_n222), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT12), .B1(new_n417), .B2(KEYINPUT79), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(KEYINPUT79), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n370), .A2(G68), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT78), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n416), .A2(new_n420), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n267), .A2(KEYINPUT76), .A3(new_n382), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G238), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT76), .B1(new_n267), .B2(new_n382), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n380), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT77), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT77), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n380), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n385), .A2(G232), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n301), .A2(G226), .A3(new_n263), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n268), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT13), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT13), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(G179), .A3(new_n441), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n432), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n445), .B2(KEYINPUT14), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n441), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(G169), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n424), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(G200), .B1(new_n443), .B2(new_n444), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n439), .A2(G190), .A3(new_n441), .ZN(new_n452));
  INV_X1    g0252(.A(new_n424), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(G58), .B(G68), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G20), .B1(G159), .B2(new_n366), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n296), .A2(new_n219), .A3(new_n300), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT7), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n298), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n248), .A2(KEYINPUT82), .A3(G33), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(G33), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n459), .A2(G20), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n458), .A2(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n457), .B1(new_n466), .B2(new_n222), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT16), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n257), .A2(new_n459), .A3(new_n219), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G68), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n459), .B1(new_n257), .B2(new_n219), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT16), .B(new_n457), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n474), .A2(new_n292), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT83), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n467), .A2(new_n476), .A3(new_n468), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n360), .A2(new_n362), .ZN(new_n479));
  INV_X1    g0279(.A(new_n330), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n479), .B2(new_n370), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT84), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n380), .B1(new_n230), .B2(new_n383), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G87), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n263), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n257), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n487), .B2(new_n268), .ZN(new_n488));
  INV_X1    g0288(.A(G190), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n488), .A2(G200), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n483), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n489), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(KEYINPUT84), .C1(G200), .C2(new_n488), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n478), .A2(new_n482), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n482), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n476), .B1(new_n467), .B2(new_n468), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n474), .A2(new_n292), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n501), .B2(new_n477), .ZN(new_n502));
  INV_X1    g0302(.A(G169), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n488), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(G179), .B2(new_n488), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT18), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n492), .A2(new_n494), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n507), .A3(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n478), .A2(new_n482), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT18), .ZN(new_n510));
  INV_X1    g0310(.A(new_n505), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n497), .A2(new_n506), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n358), .A2(new_n413), .B1(new_n219), .B2(new_n206), .ZN(new_n514));
  XOR2_X1   g0314(.A(KEYINPUT15), .B(G87), .Z(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(new_n361), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n293), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n330), .A2(new_n206), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n371), .B2(new_n206), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n380), .B1(new_n205), .B2(new_n383), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n385), .A2(G238), .B1(new_n388), .B2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n230), .B2(new_n391), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n524), .B2(new_n268), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n521), .B1(new_n525), .B2(G169), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n287), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(KEYINPUT73), .A3(new_n287), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(G190), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n520), .C1(new_n353), .C2(new_n525), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR4_X1   g0335(.A1(new_n411), .A2(new_n455), .A3(new_n513), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n282), .A2(new_n267), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n280), .B1(new_n537), .B2(new_n258), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT85), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n346), .A2(G244), .A3(new_n347), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n343), .A2(new_n344), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n385), .B2(G250), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  INV_X1    g0346(.A(G244), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n301), .A2(new_n263), .A3(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n261), .A2(new_n262), .A3(new_n547), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n550), .A2(new_n252), .A3(new_n254), .A4(new_n256), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n542), .A2(new_n545), .A3(new_n549), .A4(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n538), .B1(new_n553), .B2(new_n268), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT87), .B1(new_n554), .B2(new_n353), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT87), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT85), .B1(new_n551), .B2(new_n546), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n549), .A2(new_n560), .A3(new_n543), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n267), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n556), .B(G200), .C1(new_n562), .C2(new_n538), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n554), .A2(G190), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n480), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n332), .B2(G97), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  INV_X1    g0367(.A(G97), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n567), .A2(new_n568), .A3(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(G97), .B(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n571), .A2(new_n219), .B1(new_n206), .B2(new_n413), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n458), .A2(new_n459), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n464), .A2(new_n465), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n575), .B2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n566), .B1(new_n576), .B2(new_n293), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n555), .A2(new_n563), .A3(new_n564), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n554), .A2(new_n287), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n577), .C1(G169), .C2(new_n554), .ZN(new_n581));
  INV_X1    g0381(.A(new_n275), .ZN(new_n582));
  OAI21_X1  g0382(.A(G250), .B1(new_n273), .B2(G1), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n268), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n263), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n585), .A2(new_n257), .B1(new_n255), .B2(new_n318), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n584), .B1(new_n586), .B2(new_n268), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G169), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n287), .B2(new_n587), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n345), .A2(KEYINPUT89), .A3(new_n219), .A4(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT89), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n305), .B2(new_n222), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT19), .B1(new_n361), .B2(G97), .ZN(new_n593));
  NAND3_X1  g0393(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n219), .ZN(new_n595));
  NOR3_X1   g0395(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT88), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n219), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT88), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n568), .A2(new_n314), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(G87), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n593), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n590), .A2(new_n592), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n292), .ZN(new_n604));
  INV_X1    g0404(.A(new_n515), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n330), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n332), .A2(new_n515), .ZN(new_n607));
  AND4_X1   g0407(.A1(KEYINPUT90), .A2(new_n604), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n603), .A2(new_n292), .B1(new_n330), .B2(new_n605), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT90), .B1(new_n609), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n589), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n332), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n306), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n587), .A2(G190), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n353), .B2(new_n587), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n579), .A2(new_n581), .A3(new_n611), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n282), .A2(G270), .A3(new_n267), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n280), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT91), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT91), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n621), .A3(new_n280), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n296), .A2(G303), .A3(new_n300), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT92), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n263), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n624), .B(new_n625), .C1(new_n257), .C2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n624), .B1(new_n257), .B2(new_n626), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n267), .B1(new_n628), .B2(KEYINPUT92), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n543), .B(new_n219), .C1(G33), .C2(new_n568), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n292), .C1(new_n219), .C2(G116), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT20), .Z(new_n633));
  NOR2_X1   g0433(.A1(new_n480), .A2(G116), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n332), .B2(G116), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n630), .A2(G179), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(G169), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT21), .B1(new_n638), .B2(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n628), .A2(KEYINPUT92), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n268), .A3(new_n627), .ZN(new_n641));
  INV_X1    g0441(.A(new_n622), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n621), .B1(new_n618), .B2(new_n280), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(G169), .A4(new_n636), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n637), .B1(new_n639), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n636), .B1(new_n645), .B2(G200), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n489), .B2(new_n645), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n357), .A2(new_n536), .A3(new_n617), .A4(new_n651), .ZN(G372));
  AND2_X1   g0452(.A1(new_n506), .A2(new_n512), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n448), .A2(new_n447), .A3(G169), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n442), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n656), .A2(new_n424), .B1(new_n531), .B2(new_n454), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n497), .A2(new_n508), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT95), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n398), .A2(new_n405), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n659), .A2(new_n660), .B1(new_n397), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n409), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n611), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n577), .B1(new_n554), .B2(G169), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n562), .A2(G179), .A3(new_n538), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n611), .A3(new_n616), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n668), .A2(new_n611), .A3(new_n616), .A4(KEYINPUT26), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n665), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n338), .A2(new_n648), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n617), .A2(new_n356), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n536), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n664), .A2(new_n677), .ZN(G369));
  NAND3_X1  g0478(.A1(new_n331), .A2(new_n219), .A3(G13), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n636), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n651), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n648), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n341), .A2(new_n336), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n684), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n357), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n338), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n648), .A2(new_n684), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n357), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n690), .A2(new_n290), .A3(new_n692), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  NAND2_X1  g0500(.A1(new_n215), .A2(new_n266), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n596), .A2(new_n318), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n226), .B2(new_n701), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n675), .B1(new_n673), .B2(new_n707), .ZN(new_n708));
  AOI211_X1 g0508(.A(KEYINPUT97), .B(new_n665), .C1(new_n671), .C2(new_n672), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT29), .B(new_n692), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n676), .A2(new_n692), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n617), .A2(new_n357), .A3(new_n651), .A4(new_n692), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(new_n584), .ZN(new_n716));
  INV_X1    g0516(.A(G238), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n348), .A2(new_n717), .B1(new_n547), .B2(new_n259), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n319), .B1(new_n345), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n719), .B2(new_n267), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n352), .A2(new_n287), .A3(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n554), .A2(new_n630), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n553), .A2(new_n268), .ZN(new_n723));
  INV_X1    g0523(.A(new_n538), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n641), .A2(new_n288), .A3(new_n587), .A4(new_n644), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT30), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n269), .A2(G179), .A3(new_n284), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n720), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n554), .A2(new_n729), .A3(new_n630), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n722), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT96), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n684), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(KEYINPUT96), .B(new_n722), .C1(new_n727), .C2(new_n731), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n715), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n722), .ZN(new_n737));
  AND4_X1   g0537(.A1(new_n288), .A2(new_n641), .A3(new_n587), .A4(new_n644), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n730), .B1(new_n738), .B2(new_n554), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n730), .A2(new_n554), .A3(new_n630), .A4(new_n729), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n714), .A2(new_n736), .A3(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n710), .A2(new_n713), .B1(G330), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n706), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(new_n701), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n329), .A2(new_n273), .A3(G20), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT98), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT98), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(G1), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n215), .A2(new_n301), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n215), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n242), .A2(G45), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n215), .A2(new_n257), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n226), .A2(new_n379), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT99), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n218), .B1(G20), .B2(new_n503), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n759), .B2(new_n760), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n751), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n219), .A2(G190), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT103), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n770), .A2(G179), .A3(new_n353), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n219), .A2(new_n489), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n287), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT100), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n775), .A2(new_n287), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n776), .A2(new_n769), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n388), .B1(new_n785), .B2(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(KEYINPUT33), .A2(G317), .ZN(new_n792));
  AND2_X1   g0592(.A1(KEYINPUT33), .A2(G317), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n219), .B1(new_n796), .B2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n790), .A2(new_n489), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n794), .B1(new_n795), .B2(new_n797), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NOR4_X1   g0601(.A1(new_n774), .A2(new_n784), .A3(new_n789), .A4(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n770), .A2(G179), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT104), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT104), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G329), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n808), .A2(G159), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT32), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n771), .A2(G107), .ZN(new_n817));
  INV_X1    g0617(.A(new_n786), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n388), .B1(G87), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n797), .A2(new_n568), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n791), .B2(G68), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n816), .A2(new_n817), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n782), .ZN(new_n823));
  INV_X1    g0623(.A(new_n788), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n823), .A2(G58), .B1(G77), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(KEYINPUT101), .B1(G50), .B2(new_n799), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(KEYINPUT101), .B2(new_n825), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT102), .Z(new_n828));
  OAI21_X1  g0628(.A(new_n814), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n768), .B1(new_n829), .B2(new_n765), .ZN(new_n830));
  INV_X1    g0630(.A(new_n764), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n687), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n687), .A2(G330), .ZN(new_n833));
  INV_X1    g0633(.A(new_n751), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n688), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(G396));
  NAND3_X1  g0636(.A1(new_n532), .A2(new_n534), .A3(new_n692), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n613), .A2(new_n615), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n609), .A2(new_n607), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT90), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n609), .A2(KEYINPUT90), .A3(new_n607), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n839), .B1(new_n844), .B2(new_n589), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT26), .B1(new_n845), .B2(new_n668), .ZN(new_n846));
  INV_X1    g0646(.A(new_n672), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n611), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n845), .A2(new_n356), .A3(new_n579), .A4(new_n581), .ZN(new_n849));
  INV_X1    g0649(.A(new_n674), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n838), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n711), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n532), .B(new_n534), .C1(new_n520), .C2(new_n692), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n531), .A2(new_n521), .A3(new_n684), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n743), .A2(G330), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n751), .B1(new_n857), .B2(new_n858), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n854), .A2(new_n855), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n762), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n765), .A2(new_n762), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT106), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n751), .B1(G77), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n824), .A2(G159), .B1(G137), .B2(new_n799), .ZN(new_n867));
  INV_X1    g0667(.A(G150), .ZN(new_n868));
  INV_X1    g0668(.A(new_n791), .ZN(new_n869));
  INV_X1    g0669(.A(G143), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n867), .B1(new_n868), .B2(new_n869), .C1(new_n782), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(KEYINPUT108), .B(KEYINPUT34), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n772), .A2(new_n222), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n345), .B1(new_n364), .B2(new_n786), .C1(new_n221), .C2(new_n797), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n872), .B2(new_n873), .ZN(new_n878));
  INV_X1    g0678(.A(G132), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n812), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n812), .A2(new_n787), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n772), .A2(new_n306), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G294), .B2(new_n823), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n869), .A2(new_n773), .B1(new_n800), .B2(new_n785), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n820), .B(new_n884), .C1(G116), .C2(new_n824), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n301), .B1(G107), .B2(new_n818), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT107), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n878), .A2(new_n880), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n866), .B1(new_n889), .B2(new_n765), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n860), .A2(new_n861), .B1(new_n863), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  INV_X1    g0692(.A(new_n571), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n893), .A2(KEYINPUT35), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(KEYINPUT35), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(G116), .A3(new_n220), .A4(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT36), .Z(new_n897));
  OAI211_X1 g0697(.A(new_n227), .B(G77), .C1(new_n221), .C2(new_n222), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n364), .A2(G68), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n331), .B(G13), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n457), .B1(new_n472), .B2(new_n473), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n468), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n482), .B1(new_n903), .B2(new_n500), .ZN(new_n904));
  INV_X1    g0704(.A(new_n682), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n513), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n509), .A2(new_n511), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n509), .A2(new_n905), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n495), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n904), .B1(new_n511), .B2(new_n905), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n495), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n909), .A3(new_n495), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  INV_X1    g0718(.A(new_n909), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n911), .B1(new_n513), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n916), .B1(new_n920), .B2(KEYINPUT38), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n656), .A2(new_n424), .A3(new_n692), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT112), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n907), .A2(new_n915), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n923), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n916), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n454), .A2(new_n654), .A3(new_n442), .A4(new_n655), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n453), .A2(new_n692), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT110), .ZN(new_n937));
  INV_X1    g0737(.A(new_n935), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n450), .A2(new_n454), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT110), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n940), .A3(new_n935), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT109), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n531), .A2(new_n692), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n943), .B1(new_n852), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n837), .B1(new_n673), .B2(new_n675), .ZN(new_n946));
  INV_X1    g0746(.A(new_n944), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n946), .A2(KEYINPUT109), .A3(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n933), .B(new_n942), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n653), .A2(new_n905), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n932), .B1(new_n952), .B2(KEYINPUT111), .ZN(new_n953));
  INV_X1    g0753(.A(new_n942), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n852), .A2(new_n943), .A3(new_n944), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT109), .B1(new_n946), .B2(new_n947), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n950), .B1(new_n957), .B2(new_n933), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT111), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n710), .A2(new_n536), .A3(new_n713), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n664), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(G330), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n918), .A2(new_n911), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n513), .A2(new_n919), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT38), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n732), .A2(new_n733), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n971), .A2(KEYINPUT31), .A3(new_n684), .A4(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n714), .A2(new_n736), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n942), .A2(new_n974), .A3(new_n856), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT40), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT40), .B1(new_n929), .B2(new_n916), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n942), .A2(new_n974), .A3(new_n856), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n536), .A2(new_n974), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n965), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n980), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n964), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(G1), .B1(new_n329), .B2(G20), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n964), .A2(new_n983), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n901), .B1(new_n986), .B2(new_n987), .ZN(G367));
  NOR2_X1   g0788(.A1(new_n237), .A2(new_n756), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n766), .B1(new_n215), .B2(new_n605), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n772), .A2(new_n568), .B1(new_n785), .B2(new_n782), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n786), .A2(new_n318), .ZN(new_n992));
  INV_X1    g0792(.A(new_n797), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n992), .A2(KEYINPUT46), .B1(G107), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n787), .B2(new_n800), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n257), .B1(new_n773), .B2(new_n788), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n992), .A2(KEYINPUT46), .B1(new_n795), .B2(new_n869), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n991), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(G317), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n807), .ZN(new_n1000));
  INV_X1    g0800(.A(G137), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n807), .A2(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n301), .B1(new_n364), .B2(new_n788), .C1(new_n221), .C2(new_n786), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G150), .B2(new_n823), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n797), .A2(new_n222), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n800), .A2(new_n870), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G159), .C2(new_n791), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n771), .A2(G77), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1000), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  INV_X1    g0811(.A(new_n765), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n751), .B1(new_n989), .B2(new_n990), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT114), .Z(new_n1014));
  AND2_X1   g0814(.A1(new_n613), .A2(new_n684), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n665), .A2(new_n839), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n665), .A2(new_n1015), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n764), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n579), .B(new_n581), .C1(new_n578), .C2(new_n692), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n668), .A2(new_n684), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n699), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n699), .A2(new_n1022), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n695), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1024), .A2(new_n695), .A3(new_n1027), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n697), .B1(new_n694), .B2(new_n696), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(new_n689), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n744), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n744), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n750), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1022), .A2(new_n357), .A3(new_n696), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT42), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n581), .B1(new_n1020), .B2(new_n338), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n692), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(KEYINPUT42), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT113), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT43), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1048), .A2(KEYINPUT43), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1029), .B(new_n1022), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1022), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1050), .B1(new_n695), .B2(new_n1055), .C1(new_n1052), .C2(new_n1047), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1019), .B1(new_n1039), .B2(new_n1057), .ZN(G387));
  OR2_X1    g0858(.A1(new_n694), .A2(new_n831), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n752), .A2(new_n703), .B1(G107), .B2(new_n215), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n233), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n379), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT115), .Z(new_n1063));
  NOR2_X1   g0863(.A1(new_n358), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  AOI211_X1 g0865(.A(G45), .B(new_n702), .C1(G68), .C2(G77), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n756), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1060), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n766), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n751), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G159), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n800), .A2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n772), .A2(new_n568), .B1(KEYINPUT117), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n605), .A2(new_n797), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n345), .B1(new_n222), .B2(new_n788), .C1(new_n206), .C2(new_n786), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n782), .B2(new_n364), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n479), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n791), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT116), .B(G150), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1076), .B(new_n1080), .C1(new_n807), .C2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n786), .A2(new_n795), .B1(new_n797), .B2(new_n773), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n824), .A2(G303), .B1(G311), .B2(new_n791), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n783), .B2(new_n800), .C1(new_n782), .C2(new_n999), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT48), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT49), .Z(new_n1089));
  OAI221_X1 g0889(.A(new_n257), .B1(new_n318), .B2(new_n772), .C1(new_n807), .C2(new_n798), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1070), .B1(new_n1091), .B2(new_n765), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1034), .A2(new_n750), .B1(new_n1059), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1035), .A2(new_n746), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1034), .A2(new_n744), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(G393));
  INV_X1    g0896(.A(KEYINPUT118), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n746), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n746), .A4(new_n1098), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1055), .A2(new_n764), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n245), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n766), .B1(new_n568), .B2(new_n215), .C1(new_n1106), .C2(new_n756), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n751), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n786), .A2(new_n222), .B1(new_n788), .B2(new_n358), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n993), .A2(G77), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n869), .B2(new_n364), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n882), .A2(new_n257), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n870), .B2(new_n807), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n782), .A2(new_n1071), .B1(new_n868), .B2(new_n800), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT51), .Z(new_n1115));
  AOI22_X1  g0915(.A1(new_n818), .A2(G283), .B1(new_n824), .B2(G294), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n993), .A2(G116), .B1(G303), .B2(new_n791), .ZN(new_n1117));
  AND4_X1   g0917(.A1(new_n388), .A2(new_n817), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n807), .B2(new_n783), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n782), .A2(new_n787), .B1(new_n999), .B2(new_n800), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT52), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n1113), .A2(new_n1115), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1108), .B1(new_n1122), .B2(new_n765), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1105), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n750), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1032), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1104), .A2(new_n1127), .ZN(G390));
  NAND2_X1  g0928(.A1(new_n955), .A2(new_n956), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n974), .A2(G330), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n939), .A2(new_n941), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n862), .B1(new_n1132), .B2(new_n937), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n743), .A2(G330), .A3(new_n856), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1131), .A2(new_n1133), .B1(new_n1134), .B2(new_n954), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n974), .A2(G330), .A3(new_n856), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n954), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n942), .A2(new_n743), .A3(G330), .A4(new_n856), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n692), .B(new_n856), .C1(new_n708), .C2(new_n709), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n944), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1130), .A2(new_n1135), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1131), .A2(new_n536), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n962), .A2(new_n664), .A3(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1143), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n942), .A2(new_n974), .A3(G330), .A4(new_n856), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n923), .A2(new_n930), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n957), .B2(new_n926), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n921), .A2(new_n925), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1141), .B2(new_n942), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1141), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n954), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1152), .B(new_n1138), .C1(new_n1158), .C2(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1148), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1159), .B(new_n1156), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n746), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n811), .A2(G125), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT54), .B(G143), .Z(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT120), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n771), .A2(G50), .B1(new_n1166), .B2(new_n824), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n786), .A2(new_n1081), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n879), .C2(new_n782), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n301), .B1(new_n869), .B2(new_n1001), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n800), .A2(new_n1172), .B1(new_n797), .B2(new_n1071), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n811), .A2(G294), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n782), .A2(new_n318), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n388), .B1(new_n306), .B2(new_n786), .C1(new_n568), .C2(new_n788), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1110), .B1(new_n800), .B2(new_n773), .C1(new_n314), .C2(new_n869), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n875), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1164), .A2(new_n1174), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n751), .B1(new_n1079), .B2(new_n865), .C1(new_n1180), .C2(new_n1012), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1151), .B2(new_n762), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT121), .Z(new_n1183));
  NAND3_X1  g0983(.A1(new_n1156), .A2(new_n750), .A3(new_n1159), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1163), .A2(new_n1183), .A3(new_n1184), .ZN(G378));
  NOR3_X1   g0985(.A1(new_n765), .A2(G50), .A3(new_n762), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n869), .A2(new_n568), .B1(new_n800), .B2(new_n318), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1187), .A2(new_n345), .A3(new_n1005), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n772), .A2(new_n221), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n782), .A2(new_n314), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n266), .B1(new_n786), .B2(new_n206), .C1(new_n605), .C2(new_n788), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1188), .B(new_n1192), .C1(new_n812), .C2(new_n773), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n823), .A2(G128), .B1(new_n818), .B2(new_n1166), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n824), .A2(G137), .B1(new_n993), .B2(G150), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n791), .A2(G132), .B1(new_n799), .B2(G125), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n808), .A2(G124), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n771), .C2(G159), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n266), .B1(new_n257), .B2(new_n255), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n364), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1195), .A2(new_n1196), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n834), .B(new_n1186), .C1(new_n1209), .C2(new_n765), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n373), .A2(new_n905), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n411), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n406), .A2(new_n410), .A3(new_n1211), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n762), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1210), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n931), .B1(new_n958), .B2(new_n959), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n952), .A2(KEYINPUT111), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1218), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n980), .B2(G330), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n965), .B(new_n1218), .C1(new_n976), .C2(new_n979), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1222), .A2(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1133), .A2(new_n921), .A3(new_n974), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1228), .A2(KEYINPUT40), .B1(new_n977), .B2(new_n978), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1218), .B1(new_n1229), .B2(new_n965), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n980), .A2(G330), .A3(new_n1224), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n953), .A2(new_n960), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1227), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1221), .B1(new_n1233), .B2(new_n750), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1162), .A2(new_n1145), .B1(new_n1232), .B2(new_n1227), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n746), .B1(new_n1235), .B2(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1162), .A2(new_n1145), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1237), .A2(KEYINPUT57), .A3(new_n1233), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1236), .B2(new_n1238), .ZN(G375));
  XNOR2_X1  g1039(.A(new_n750), .B(KEYINPUT122), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n954), .A2(new_n762), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n751), .B1(G68), .B2(new_n865), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n812), .A2(new_n1172), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1189), .B1(new_n791), .B2(new_n1166), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n800), .A2(new_n879), .B1(new_n797), .B2(new_n364), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n786), .A2(new_n1071), .B1(new_n788), .B2(new_n868), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n257), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1245), .B(new_n1248), .C1(new_n1001), .C2(new_n782), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n812), .A2(new_n785), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n823), .A2(G283), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n818), .A2(G97), .B1(new_n824), .B2(G107), .ZN(new_n1252));
  AND4_X1   g1052(.A1(new_n388), .A2(new_n1251), .A3(new_n1008), .A4(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1074), .B1(new_n799), .B2(G294), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n318), .C2(new_n869), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1244), .A2(new_n1249), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1243), .B1(new_n1256), .B2(new_n765), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1142), .A2(new_n1241), .B1(new_n1242), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(new_n1037), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1148), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(G381));
  INV_X1    g1063(.A(G387), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1126), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1262), .A4(new_n1266), .ZN(new_n1267));
  OR3_X1    g1067(.A1(G375), .A2(new_n1267), .A3(G378), .ZN(G407));
  AND3_X1   g1068(.A1(new_n1163), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n683), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  OAI211_X1 g1073(.A(G378), .B(new_n1234), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1233), .A2(new_n1241), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT123), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1220), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1237), .A2(new_n1038), .A3(new_n1233), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1240), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT123), .B1(new_n1279), .B2(new_n1221), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1269), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1270), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1134), .A2(new_n954), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1149), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1285), .A2(new_n1157), .B1(new_n1129), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n962), .A2(new_n664), .A3(new_n1144), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT119), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1142), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(KEYINPUT60), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1260), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n701), .B1(new_n1260), .B2(KEYINPUT60), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n891), .B1(new_n1299), .B2(new_n1259), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1297), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(G384), .A3(new_n1258), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1271), .A2(G2897), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1300), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1298), .B1(new_n1301), .B2(KEYINPUT124), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n891), .B(new_n1259), .C1(new_n1309), .C2(new_n1303), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1304), .B2(new_n1258), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G2897), .B(new_n1271), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1300), .A2(new_n1313), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1284), .A2(new_n1308), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1283), .A2(new_n1317), .A3(new_n1270), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1283), .A2(new_n1317), .A3(new_n1320), .A4(new_n1270), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1315), .A2(new_n1316), .A3(new_n1319), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G390), .A2(new_n1264), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1265), .A2(G387), .ZN(new_n1324));
  XOR2_X1   g1124(.A(G393), .B(G396), .Z(new_n1325));
  AND4_X1   g1125(.A1(KEYINPUT126), .A2(new_n1323), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1265), .B2(G387), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n1328), .A2(new_n1325), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1322), .A2(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1283), .A2(new_n1317), .A3(KEYINPUT63), .A4(new_n1270), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1318), .A2(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1334), .A2(new_n1316), .A3(new_n1315), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1332), .A2(new_n1337), .ZN(G405));
  OR2_X1    g1138(.A1(new_n1330), .A2(KEYINPUT127), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1330), .A2(KEYINPUT127), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(G375), .A2(new_n1269), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1274), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1342), .A2(new_n1317), .ZN(new_n1343));
  AOI211_X1 g1143(.A(new_n1311), .B(new_n1310), .C1(new_n1341), .C2(new_n1274), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1339), .B(new_n1340), .C1(new_n1343), .C2(new_n1344), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1343), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(KEYINPUT127), .A3(new_n1330), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1345), .A2(new_n1347), .ZN(G402));
endmodule


