//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n590, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT70), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n458), .A2(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(KEYINPUT71), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n466), .ZN(new_n482));
  INV_X1    g057(.A(G137), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n478), .A2(new_n484), .ZN(G160));
  XNOR2_X1  g060(.A(new_n482), .B(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n468), .A2(new_n469), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n466), .ZN(new_n489));
  MUX2_X1   g064(.A(G100), .B(G112), .S(G2105), .Z(new_n490));
  AOI22_X1  g065(.A1(new_n489), .A2(G124), .B1(G2104), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n487), .A2(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n481), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n481), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n466), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n470), .A2(new_n475), .A3(G138), .A4(new_n466), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G50), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n500), .A2(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT74), .Z(new_n522));
  NOR2_X1   g097(.A1(new_n501), .A2(new_n502), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n506), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n524), .A2(G51), .B1(new_n510), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n515), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(G52), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n503), .A2(new_n510), .A3(G90), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n531), .A2(KEYINPUT75), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT75), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(KEYINPUT76), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G171));
  XOR2_X1   g114(.A(KEYINPUT77), .B(G43), .Z(new_n540));
  NOR2_X1   g115(.A1(new_n504), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n515), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n523), .B1(new_n507), .B2(new_n509), .ZN(new_n544));
  AOI211_X1 g119(.A(new_n541), .B(new_n543), .C1(G81), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n552), .B(new_n553), .C1(new_n504), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n544), .A2(G91), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n554), .B1(KEYINPUT78), .B2(KEYINPUT9), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n524), .B(new_n557), .C1(KEYINPUT78), .C2(KEYINPUT9), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n515), .B1(new_n560), .B2(KEYINPUT79), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(KEYINPUT79), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n544), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n524), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n515), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n544), .A2(G86), .B1(new_n524), .B2(G48), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n544), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n515), .B2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(new_n524), .A2(G54), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n515), .ZN(new_n579));
  XOR2_X1   g154(.A(new_n579), .B(KEYINPUT80), .Z(new_n580));
  NAND2_X1  g155(.A1(new_n544), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT10), .Z(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n584), .B2(G171), .ZN(G284));
  OAI21_X1  g161(.A(new_n585), .B1(new_n584), .B2(G171), .ZN(G321));
  AND2_X1   g162(.A1(new_n559), .A2(new_n562), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT81), .B1(new_n588), .B2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  MUX2_X1   g165(.A(KEYINPUT81), .B(new_n589), .S(new_n590), .Z(G297));
  XOR2_X1   g166(.A(G297), .B(KEYINPUT82), .Z(G280));
  AND2_X1   g167(.A1(new_n580), .A2(new_n582), .ZN(new_n593));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n545), .A2(new_n584), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n584), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g174(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g175(.A1(new_n470), .A2(new_n475), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(new_n479), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT12), .Z(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT13), .Z(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(G2100), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n489), .A2(G123), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT85), .Z(new_n607));
  MUX2_X1   g182(.A(G99), .B(G111), .S(G2105), .Z(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(G2104), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n486), .A2(G135), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT84), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(KEYINPUT15), .B(G2435), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT86), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(G2427), .B(G2430), .Z(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(KEYINPUT14), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2451), .B(G2454), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT16), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n621), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT87), .Z(new_n629));
  INV_X1    g204(.A(G14), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(G401));
  XNOR2_X1  g208(.A(G2072), .B(G2078), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT17), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NOR3_X1   g213(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n638), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(new_n637), .C1(new_n634), .C2(new_n638), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n634), .A3(new_n638), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT18), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(G227));
  XOR2_X1   g222(.A(G1956), .B(G2474), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT89), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1961), .B(G1966), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT90), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT20), .Z(new_n656));
  OR2_X1    g231(.A1(new_n649), .A2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n654), .A3(new_n652), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n656), .B(new_n658), .C1(new_n654), .C2(new_n657), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G229));
  NOR2_X1   g241(.A1(G29), .A2(G35), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(G162), .B2(G29), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT29), .Z(new_n669));
  INV_X1    g244(.A(G2090), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT99), .Z(new_n672));
  INV_X1    g247(.A(G1961), .ZN(new_n673));
  NOR2_X1   g248(.A1(G5), .A2(G16), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G171), .B2(G16), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n486), .A2(G139), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n479), .A2(G103), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT25), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n601), .A2(G127), .ZN(new_n681));
  NAND2_X1  g256(.A1(G115), .A2(G2104), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n466), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n678), .B(new_n680), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(G33), .B(new_n687), .S(G29), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2072), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G1961), .B2(new_n675), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n486), .A2(G141), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n479), .A2(G105), .ZN(new_n692));
  NAND3_X1  g267(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT26), .ZN(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(G129), .C2(new_n489), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G29), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(KEYINPUT97), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G29), .B2(G32), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n699), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT27), .B(G1996), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n704), .ZN(new_n706));
  OR2_X1    g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  NAND2_X1  g282(.A1(KEYINPUT24), .A2(G34), .ZN(new_n708));
  AOI21_X1  g283(.A(G29), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G160), .B2(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G2084), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G19), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n545), .B2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1341), .Z(new_n714));
  NAND4_X1  g289(.A1(new_n705), .A2(new_n706), .A3(new_n711), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n669), .A2(new_n670), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G1966), .ZN(new_n720));
  NOR2_X1   g295(.A1(G27), .A2(G29), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G164), .B2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT98), .B(G2078), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n716), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G11), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT30), .B(G28), .Z(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G29), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n612), .B2(G29), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n729), .B1(G2084), .B2(new_n710), .C1(G1966), .C2(new_n719), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n715), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT95), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n486), .A2(G140), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G104), .B(G116), .S(G2105), .Z(new_n739));
  AOI22_X1  g314(.A1(new_n489), .A2(G128), .B1(G2104), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n735), .B1(new_n742), .B2(new_n732), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  NOR2_X1   g319(.A1(G4), .A2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n593), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n717), .A2(G20), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT23), .Z(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G299), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1956), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n744), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n677), .A2(new_n690), .A3(new_n731), .A4(new_n753), .ZN(new_n754));
  MUX2_X1   g329(.A(G6), .B(G305), .S(G16), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT32), .B(G1981), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n717), .A2(G23), .ZN(new_n759));
  INV_X1    g334(.A(G288), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n717), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT33), .B(G1976), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G22), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G166), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1971), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n758), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT34), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G25), .A2(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n489), .A2(G119), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT91), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n486), .A2(G131), .ZN(new_n773));
  MUX2_X1   g348(.A(G95), .B(G107), .S(G2105), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2104), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n770), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(G290), .A2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G24), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT92), .B1(new_n782), .B2(G16), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n782), .A2(KEYINPUT92), .A3(G16), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1986), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n769), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n767), .A2(new_n768), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n787), .A2(KEYINPUT36), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT36), .B1(new_n787), .B2(new_n788), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n754), .B1(new_n790), .B2(new_n791), .ZN(G311));
  INV_X1    g367(.A(new_n754), .ZN(new_n793));
  INV_X1    g368(.A(new_n791), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n789), .ZN(G150));
  AOI22_X1  g370(.A1(new_n544), .A2(G93), .B1(new_n524), .B2(G55), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT100), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n515), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT101), .B(G860), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT37), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n800), .B(new_n545), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n593), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n801), .B1(new_n808), .B2(KEYINPUT39), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(G145));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT102), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n687), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n738), .A2(G164), .A3(new_n740), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(G164), .B1(new_n738), .B2(new_n740), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n697), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n820), .A2(new_n696), .A3(new_n816), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n486), .A2(G142), .ZN(new_n823));
  MUX2_X1   g398(.A(G106), .B(G118), .S(G2105), .Z(new_n824));
  AOI22_X1  g399(.A1(new_n489), .A2(G130), .B1(G2104), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n603), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n776), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n687), .A2(new_n813), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n822), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n828), .B1(new_n822), .B2(new_n829), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n815), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n822), .A2(new_n829), .ZN(new_n834));
  INV_X1    g409(.A(new_n828), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n836), .A2(new_n814), .A3(new_n830), .ZN(new_n837));
  INV_X1    g412(.A(new_n612), .ZN(new_n838));
  XOR2_X1   g413(.A(G162), .B(G160), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n833), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n840), .B1(new_n833), .B2(new_n837), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n812), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(KEYINPUT40), .A3(new_n842), .A4(new_n841), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n845), .A2(new_n847), .ZN(G395));
  OR2_X1    g423(.A1(new_n800), .A2(G868), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n583), .A2(G299), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n583), .A2(G299), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n593), .A2(new_n588), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n855), .A2(KEYINPUT41), .A3(new_n851), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(new_n855), .B2(new_n851), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n805), .B(new_n597), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n854), .B(new_n858), .S(new_n859), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n760), .B(G290), .ZN(new_n861));
  XNOR2_X1  g436(.A(G305), .B(G166), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT103), .Z(new_n864));
  OR2_X1    g439(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n860), .B(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n850), .B1(new_n868), .B2(G868), .ZN(G295));
  AOI21_X1  g444(.A(new_n850), .B1(new_n868), .B2(G868), .ZN(G331));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g446(.A1(G171), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n537), .A2(KEYINPUT104), .A3(new_n538), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(G168), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(G301), .A2(KEYINPUT104), .A3(G286), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n805), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n805), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n858), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n854), .A3(new_n876), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n881), .A3(new_n866), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n842), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n866), .B1(new_n879), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n842), .A4(new_n882), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n885), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(G397));
  XNOR2_X1  g467(.A(new_n741), .B(G2067), .ZN(new_n893));
  OAI21_X1  g468(.A(G126), .B1(new_n468), .B2(new_n469), .ZN(new_n894));
  NAND2_X1  g469(.A1(G114), .A2(G2104), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n466), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT4), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n498), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(KEYINPUT4), .A2(G138), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n488), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n494), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n466), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT105), .B(G1384), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT45), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G40), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n478), .A2(new_n906), .A3(new_n484), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(G1996), .A3(new_n696), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT106), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(G1996), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n697), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n776), .B(new_n779), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n909), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G1986), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n484), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n476), .A2(new_n477), .ZN(new_n924));
  OAI211_X1 g499(.A(G40), .B(new_n923), .C1(new_n924), .C2(new_n466), .ZN(new_n925));
  OAI21_X1  g500(.A(G8), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n760), .A2(G1976), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n760), .B2(G1976), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT49), .ZN(new_n932));
  INV_X1    g507(.A(G1981), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n571), .A2(new_n933), .A3(new_n572), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n571), .B2(new_n572), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(KEYINPUT49), .A3(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n929), .A2(new_n931), .B1(new_n940), .B2(new_n926), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n929), .A2(KEYINPUT52), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n929), .A2(new_n944), .A3(KEYINPUT52), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G8), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n898), .B2(new_n902), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n907), .B1(new_n948), .B2(KEYINPUT45), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n903), .A2(KEYINPUT45), .A3(new_n904), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1971), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n955));
  AOI21_X1  g530(.A(new_n925), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n670), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n947), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(G166), .B2(new_n947), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n907), .B1(new_n948), .B2(new_n955), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n967), .A2(KEYINPUT111), .B1(new_n968), .B2(new_n948), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n907), .B(new_n970), .C1(new_n948), .C2(new_n955), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n670), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n947), .B1(new_n972), .B2(new_n954), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n946), .B(new_n966), .C1(new_n973), .C2(new_n963), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(G164), .B2(G1384), .ZN(new_n976));
  INV_X1    g551(.A(G2078), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(new_n977), .A3(new_n907), .A4(new_n951), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G1961), .B1(new_n956), .B2(new_n957), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n975), .B(G1384), .C1(new_n898), .C2(new_n902), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n979), .A2(G2078), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n949), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT121), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n903), .A2(new_n921), .A3(new_n955), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n907), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n948), .A2(new_n968), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n673), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT121), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n948), .A2(KEYINPUT45), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n976), .A2(new_n993), .A3(new_n907), .A4(new_n984), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n981), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT122), .B1(new_n996), .B2(G301), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n980), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT122), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(G171), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n951), .A2(new_n907), .A3(new_n984), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n980), .B(new_n991), .C1(new_n905), .C2(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n997), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n1004), .B2(G171), .ZN(new_n1010));
  OAI211_X1 g585(.A(G301), .B(new_n980), .C1(new_n998), .C2(new_n999), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1966), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n949), .B2(new_n983), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT112), .B(G2084), .Z(new_n1017));
  NAND4_X1  g592(.A1(new_n957), .A2(new_n907), .A3(new_n988), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(KEYINPUT118), .A3(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n1014), .C1(new_n1023), .C2(G286), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G286), .A2(G8), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(G8), .A3(G286), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1012), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n988), .B(new_n907), .C1(new_n968), .C2(new_n948), .ZN(new_n1032));
  INV_X1    g607(.A(G1348), .ZN(new_n1033));
  INV_X1    g608(.A(G2067), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n922), .A2(new_n925), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1032), .A2(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n593), .B1(new_n1036), .B2(KEYINPUT60), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n989), .B2(new_n990), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1034), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(KEYINPUT60), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT117), .B1(new_n1036), .B2(KEYINPUT60), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1996), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n976), .A2(new_n1045), .A3(new_n907), .A4(new_n951), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT58), .B(G1341), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1035), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n545), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT59), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1051), .A3(new_n545), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n583), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1036), .A2(KEYINPUT117), .A3(KEYINPUT60), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1044), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n1061));
  XNOR2_X1  g636(.A(G299), .B(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n976), .A2(new_n907), .A3(new_n951), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n950), .A2(KEYINPUT115), .A3(new_n951), .A4(new_n1063), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1956), .B1(new_n969), .B2(new_n971), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1062), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n967), .A2(KEYINPUT111), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n948), .A2(new_n968), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n971), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n751), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n588), .B(new_n1061), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1070), .A2(new_n1076), .A3(KEYINPUT61), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT61), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1060), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1036), .A2(new_n583), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1074), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1062), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1076), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1070), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT116), .B(new_n1076), .C1(new_n1086), .C2(new_n1081), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1008), .B(new_n1031), .C1(new_n1079), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1022), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1013), .B1(new_n1092), .B2(new_n1027), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1028), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1030), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1029), .A2(new_n1097), .A3(new_n1030), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n997), .A2(new_n1002), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n974), .B1(new_n1089), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1025), .A2(G286), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n974), .B2(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n959), .A2(new_n963), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n959), .B2(new_n965), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(new_n946), .A3(new_n1107), .A4(new_n1103), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(KEYINPUT113), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(KEYINPUT113), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G288), .A2(G1976), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n940), .B2(new_n926), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n934), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(KEYINPUT110), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n926), .B1(new_n1114), .B2(KEYINPUT110), .ZN(new_n1116));
  INV_X1    g691(.A(new_n966), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1117), .B2(new_n946), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1111), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n920), .B1(new_n1101), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n909), .B1(new_n893), .B2(new_n696), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n913), .A2(KEYINPUT46), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n913), .A2(KEYINPUT46), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT125), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1121), .A2(new_n1126), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n918), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT126), .B1(new_n915), .B2(new_n917), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n908), .A2(G1986), .A3(G290), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1135), .B(new_n1136), .Z(new_n1137));
  NOR3_X1   g712(.A1(new_n1133), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n777), .A2(new_n779), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT123), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n742), .A2(new_n1034), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n908), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1131), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1120), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g720(.A1(G227), .A2(new_n464), .ZN(new_n1147));
  NOR3_X1   g721(.A1(G229), .A2(new_n1147), .A3(G401), .ZN(new_n1148));
  OAI21_X1  g722(.A(new_n1148), .B1(new_n843), .B2(new_n844), .ZN(new_n1149));
  AOI21_X1  g723(.A(new_n1149), .B1(new_n885), .B2(new_n888), .ZN(G308));
  NAND2_X1  g724(.A1(new_n885), .A2(new_n888), .ZN(new_n1151));
  OAI211_X1 g725(.A(new_n1151), .B(new_n1148), .C1(new_n844), .C2(new_n843), .ZN(G225));
endmodule


