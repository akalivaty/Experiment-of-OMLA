//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT33), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g011(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n216), .B2(new_n217), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n214), .A2(new_n215), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n204), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n211), .A2(new_n204), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n213), .A3(new_n218), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G127gat), .B(G134gat), .Z(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT71), .ZN(new_n233));
  INV_X1    g032(.A(G113gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(G120gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n236));
  INV_X1    g035(.A(G120gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(G113gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(new_n238), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n231), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT27), .B(G183gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT28), .A3(new_n217), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT69), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT27), .B1(new_n216), .B2(KEYINPUT68), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n217), .B(new_n251), .C1(new_n252), .C2(KEYINPUT68), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n257), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(KEYINPUT26), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n210), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n261), .A2(new_n262), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n230), .A2(new_n247), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n224), .A2(new_n229), .B1(new_n256), .B2(new_n263), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT74), .A3(new_n247), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n230), .A2(new_n264), .ZN(new_n270));
  INV_X1    g069(.A(new_n247), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT75), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n273), .B2(new_n276), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n203), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n267), .A2(new_n272), .A3(new_n275), .A4(new_n269), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT34), .ZN(new_n281));
  XOR2_X1   g080(.A(G15gat), .B(G43gat), .Z(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n279), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n279), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT32), .B1(new_n277), .B2(new_n278), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  INV_X1    g088(.A(new_n281), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n276), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT75), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT33), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n284), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n281), .A3(new_n284), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  OAI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(KEYINPUT76), .B2(KEYINPUT22), .ZN(new_n302));
  AND2_X1   g101(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G211gat), .B(G218gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G141gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G148gat), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT79), .B(G148gat), .Z(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(new_n314), .B2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n318));
  XNOR2_X1  g117(.A(G141gat), .B(G148gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n311), .B(new_n314), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n306), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(KEYINPUT84), .B1(G228gat), .B2(G233gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(G22gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT31), .B(G50gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G22gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n324), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n317), .B1(new_n306), .B2(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n320), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n323), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G78gat), .B(G106gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n328), .A2(new_n331), .A3(new_n338), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n288), .A2(new_n298), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n334), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n245), .A2(new_n246), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT73), .B1(new_n242), .B2(new_n244), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT4), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(new_n321), .A3(new_n245), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n316), .A2(new_n242), .A3(new_n320), .A4(new_n244), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n348), .A2(new_n349), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n245), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(new_n349), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n351), .A2(new_n356), .A3(new_n349), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n352), .A2(new_n353), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n353), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G1gat), .B(G29gat), .Z(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT83), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n367), .A2(new_n376), .A3(KEYINPUT6), .A4(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT81), .B1(new_n367), .B2(new_n372), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n381));
  INV_X1    g180(.A(new_n372), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n361), .A2(new_n366), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n380), .A2(new_n383), .A3(new_n374), .A4(new_n373), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT77), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n221), .A3(new_n212), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n204), .B1(new_n228), .B2(new_n225), .ZN(new_n390));
  INV_X1    g189(.A(new_n264), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n306), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n230), .B2(new_n264), .ZN(new_n394));
  INV_X1    g193(.A(new_n386), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n390), .B2(new_n391), .ZN(new_n398));
  INV_X1    g197(.A(new_n387), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n398), .A2(new_n399), .B1(new_n270), .B2(new_n395), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n400), .B2(new_n393), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n394), .A2(new_n387), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n268), .A2(new_n386), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n306), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n396), .A3(new_n404), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n410), .A3(KEYINPUT30), .ZN(new_n411));
  OR3_X1    g210(.A1(new_n401), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n385), .A2(new_n414), .A3(KEYINPUT35), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n287), .B1(new_n285), .B2(new_n286), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n373), .A2(KEYINPUT82), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n367), .A2(new_n418), .A3(new_n372), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n380), .A2(new_n374), .A3(new_n383), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n422), .A2(new_n379), .B1(new_n412), .B2(new_n411), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n296), .A2(new_n289), .A3(new_n297), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n416), .A2(new_n423), .A3(new_n424), .A4(new_n342), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n344), .A2(new_n415), .B1(new_n425), .B2(KEYINPUT35), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n405), .B1(new_n401), .B2(KEYINPUT37), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n392), .B(new_n306), .C1(new_n394), .C2(new_n395), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(KEYINPUT37), .C1(new_n400), .C2(new_n306), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT38), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n375), .A2(new_n377), .A3(new_n410), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT37), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n409), .B2(new_n396), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT38), .B1(new_n427), .B2(new_n435), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n432), .A2(new_n433), .A3(new_n436), .A4(new_n384), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n365), .A2(new_n351), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n359), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n357), .A2(new_n349), .A3(new_n352), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT39), .A3(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n359), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n382), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT40), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n441), .A2(KEYINPUT40), .A3(new_n382), .A4(new_n443), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n373), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n342), .B1(new_n413), .B2(new_n448), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n437), .A2(new_n449), .B1(new_n423), .B2(new_n342), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n288), .B2(new_n298), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n416), .A2(KEYINPUT36), .A3(new_n424), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n202), .B1(new_n426), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n449), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n432), .A2(new_n433), .A3(new_n436), .A4(new_n384), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n420), .A2(new_n421), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n413), .B1(new_n458), .B2(new_n378), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(new_n343), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT36), .B1(new_n416), .B2(new_n424), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n425), .A2(KEYINPUT35), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n415), .A2(new_n424), .A3(new_n416), .A4(new_n342), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n466), .A3(KEYINPUT86), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G22gat), .ZN(new_n468));
  INV_X1    g267(.A(G1gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT16), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(G1gat), .B2(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G8gat), .ZN(new_n473));
  INV_X1    g272(.A(G8gat), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n471), .B(new_n474), .C1(G1gat), .C2(new_n468), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G29gat), .ZN(new_n477));
  INV_X1    g276(.A(G36gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT14), .ZN(new_n479));
  NAND2_X1  g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT15), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n479), .A2(new_n485), .A3(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n479), .A2(new_n485), .A3(KEYINPUT15), .A4(new_n480), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n486), .B(new_n487), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n489), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n491), .A3(new_n482), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n487), .B1(new_n496), .B2(new_n486), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n476), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n475), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n486), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT18), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n502), .B(KEYINPUT13), .Z(new_n506));
  INV_X1    g305(.A(new_n501), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n498), .A2(KEYINPUT18), .A3(new_n501), .A4(new_n502), .ZN(new_n510));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G197gat), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT11), .B(G169gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT12), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT88), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n510), .A2(new_n520), .A3(new_n509), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n505), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n515), .B(KEYINPUT87), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n455), .A2(new_n467), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G57gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G64gat), .ZN(new_n534));
  INV_X1    g333(.A(G64gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G57gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n531), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n532), .A2(new_n540), .A3(KEYINPUT89), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT89), .B1(new_n532), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G127gat), .ZN(new_n548));
  XOR2_X1   g347(.A(G183gat), .B(G211gat), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n548), .A2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n540), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n540), .A3(KEYINPUT89), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n499), .B1(new_n557), .B2(KEYINPUT21), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(new_n312), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n560), .B(new_n562), .Z(new_n563));
  OR3_X1    g362(.A1(new_n551), .A2(new_n552), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n551), .B2(new_n552), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT93), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT94), .B1(new_n567), .B2(KEYINPUT7), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n572), .A3(G85gat), .A4(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n574), .A3(KEYINPUT7), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n569), .A2(new_n570), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(G85gat), .ZN(new_n578));
  INV_X1    g377(.A(G92gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(KEYINPUT8), .A2(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n576), .A2(new_n582), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n586), .A2(new_n500), .B1(KEYINPUT41), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n576), .A2(new_n582), .A3(new_n580), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n582), .B1(new_n576), .B2(new_n580), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n494), .B2(new_n497), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(KEYINPUT95), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  NOR2_X1   g396(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n594), .B(KEYINPUT95), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n588), .A2(new_n592), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n599), .A2(new_n600), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n600), .A3(new_n599), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n566), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n584), .A2(new_n555), .A3(new_n556), .A4(new_n585), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n582), .A2(KEYINPUT97), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n581), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n553), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n576), .A2(new_n580), .A3(new_n613), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n557), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n553), .B1(new_n581), .B2(new_n614), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n591), .A2(new_n543), .B1(new_n624), .B2(new_n617), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n625), .A2(new_n622), .ZN(new_n626));
  XOR2_X1   g425(.A(G120gat), .B(G148gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n621), .B2(new_n622), .ZN(new_n634));
  INV_X1    g433(.A(new_n622), .ZN(new_n635));
  AOI211_X1 g434(.A(KEYINPUT99), .B(new_n635), .C1(new_n619), .C2(new_n620), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n626), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n630), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n526), .A2(new_n610), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n458), .A2(new_n378), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n469), .ZN(G1324gat));
  NOR2_X1   g443(.A1(new_n640), .A2(new_n413), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  AOI21_X1  g445(.A(KEYINPUT42), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(G8gat), .B1(new_n640), .B2(new_n413), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n650), .B2(KEYINPUT42), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT100), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n416), .A2(new_n424), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n640), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT101), .Z(new_n656));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n461), .B2(new_n462), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n452), .A2(KEYINPUT102), .A3(new_n453), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n640), .A2(new_n653), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n656), .A2(new_n663), .ZN(G1326gat));
  NOR2_X1   g463(.A1(new_n640), .A2(new_n342), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT43), .B(G22gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NAND4_X1  g466(.A1(new_n526), .A2(new_n566), .A3(new_n609), .A4(new_n639), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(G29gat), .A3(new_n642), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n658), .A2(new_n460), .A3(new_n660), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n466), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(KEYINPUT105), .A3(new_n466), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n608), .A2(KEYINPUT44), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n455), .A2(new_n467), .A3(new_n609), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n679), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT104), .B1(new_n679), .B2(KEYINPUT44), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n566), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n637), .A2(new_n638), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n631), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n683), .A2(new_n524), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(new_n641), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n671), .B1(new_n688), .B2(new_n477), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n668), .A2(G36gat), .A3(new_n413), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n687), .A2(new_n414), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n478), .ZN(G1329gat));
  NOR3_X1   g492(.A1(new_n668), .A2(G43gat), .A3(new_n654), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n662), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n697), .A3(new_n686), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G43gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n696), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n698), .A2(G43gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n695), .B1(new_n704), .B2(new_n694), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1330gat));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n682), .A2(new_n343), .A3(new_n686), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(G50gat), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n668), .A2(G50gat), .A3(new_n342), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n708), .B2(G50gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI221_X4 g512(.A(new_n710), .B1(new_n707), .B2(KEYINPUT48), .C1(new_n708), .C2(G50gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(G1331gat));
  AND2_X1   g514(.A1(new_n675), .A2(new_n676), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n566), .A2(new_n525), .A3(new_n609), .A4(new_n639), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n642), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(new_n533), .ZN(G1332gat));
  NOR2_X1   g519(.A1(new_n718), .A2(new_n413), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  AND2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n721), .B2(new_n722), .ZN(G1333gat));
  OR3_X1    g524(.A1(new_n718), .A2(G71gat), .A3(new_n654), .ZN(new_n726));
  OAI21_X1  g525(.A(G71gat), .B1(new_n718), .B2(new_n662), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1334gat));
  NOR2_X1   g529(.A1(new_n718), .A2(new_n342), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g531(.A1(new_n683), .A2(new_n525), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n609), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT51), .B1(new_n673), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n737), .B(new_n734), .C1(new_n672), .C2(new_n466), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n639), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n578), .A3(new_n641), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n683), .A2(new_n525), .A3(new_n639), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n682), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n641), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(new_n578), .ZN(G1336gat));
  NAND3_X1  g544(.A1(new_n682), .A2(new_n414), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G92gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n413), .A2(G92gat), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n685), .B(new_n748), .C1(new_n736), .C2(new_n738), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n754), .A3(KEYINPUT52), .ZN(new_n755));
  AND4_X1   g554(.A1(new_n747), .A2(new_n753), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n753), .A2(new_n755), .B1(new_n747), .B2(new_n749), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(G1337gat));
  INV_X1    g557(.A(G99gat), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n740), .A2(new_n759), .A3(new_n424), .A4(new_n416), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n743), .A2(new_n697), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n759), .ZN(G1338gat));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  INV_X1    g562(.A(G106gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n740), .A2(new_n764), .A3(new_n343), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n743), .A2(new_n343), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n763), .B(new_n765), .C1(new_n766), .C2(new_n764), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n743), .B2(new_n343), .ZN(new_n768));
  INV_X1    g567(.A(new_n765), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT53), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT10), .B1(new_n541), .B2(new_n542), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n591), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n625), .B2(new_n612), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT99), .B1(new_n775), .B2(new_n635), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n621), .A2(new_n633), .A3(new_n622), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n621), .B2(new_n622), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n619), .A2(new_n635), .A3(new_n620), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n630), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n779), .A2(new_n782), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n779), .B2(new_n782), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n524), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n787), .A2(new_n631), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n498), .A2(new_n501), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n507), .A2(new_n508), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n791), .A2(new_n502), .B1(new_n792), .B2(new_n506), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n514), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n516), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n685), .A2(new_n796), .A3(KEYINPUT112), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n639), .B2(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n608), .B1(new_n790), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n608), .A2(new_n788), .A3(new_n795), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n631), .A3(new_n787), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n683), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n566), .A2(new_n525), .A3(new_n609), .A4(new_n685), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n772), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n800), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n789), .A3(new_n631), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n609), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n803), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n566), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n805), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(KEYINPUT113), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n641), .ZN(new_n815));
  NOR4_X1   g614(.A1(new_n815), .A2(new_n654), .A3(new_n414), .A4(new_n343), .ZN(new_n816));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n525), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n642), .A2(new_n414), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n342), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n822));
  AOI211_X1 g621(.A(new_n654), .B(new_n819), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n524), .A2(new_n234), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(G1340gat));
  AOI21_X1  g624(.A(G120gat), .B1(new_n816), .B2(new_n685), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n639), .A2(new_n237), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n823), .B2(new_n827), .ZN(G1341gat));
  INV_X1    g627(.A(G127gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n816), .A2(new_n829), .A3(new_n683), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n823), .A2(new_n683), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n829), .ZN(G1342gat));
  INV_X1    g631(.A(new_n815), .ZN(new_n833));
  INV_X1    g632(.A(G134gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n414), .A2(new_n608), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n344), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT56), .Z(new_n837));
  AND2_X1   g636(.A1(new_n823), .A2(new_n609), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n834), .ZN(G1343gat));
  NOR3_X1   g638(.A1(new_n659), .A2(new_n661), .A3(new_n819), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n806), .A2(new_n343), .A3(new_n813), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n639), .A2(new_n795), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n608), .B1(new_n790), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n803), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n805), .B1(new_n847), .B2(new_n566), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n848), .A2(new_n843), .A3(new_n342), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n842), .B1(new_n841), .B2(new_n843), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n525), .B(new_n840), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n841), .A2(new_n843), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n849), .A3(new_n844), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n525), .A4(new_n840), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n858), .A3(G141gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n658), .A2(new_n343), .A3(new_n660), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n833), .A2(KEYINPUT118), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n815), .B2(new_n860), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n525), .A2(new_n307), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT116), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n413), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n859), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n852), .A2(G141gat), .ZN(new_n873));
  NOR4_X1   g672(.A1(new_n815), .A2(new_n414), .A3(new_n867), .A4(new_n860), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n876), .B2(KEYINPUT58), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n852), .B2(G141gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(KEYINPUT117), .A3(new_n870), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n871), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT120), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n871), .B(new_n882), .C1(new_n877), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(new_n309), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n856), .A2(new_n840), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n639), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n843), .B1(new_n848), .B2(new_n342), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n841), .B2(new_n843), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(new_n685), .A3(new_n840), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n865), .A2(new_n413), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n685), .A2(new_n885), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(G1345gat));
  NAND3_X1  g696(.A1(new_n865), .A2(new_n413), .A3(new_n683), .ZN(new_n898));
  INV_X1    g697(.A(new_n887), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n566), .A2(new_n312), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT121), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n898), .A2(new_n312), .B1(new_n899), .B2(new_n901), .ZN(G1346gat));
  NAND3_X1  g701(.A1(new_n865), .A2(new_n313), .A3(new_n835), .ZN(new_n903));
  OAI21_X1  g702(.A(G162gat), .B1(new_n887), .B2(new_n608), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1347gat));
  NAND2_X1  g704(.A1(new_n821), .A2(new_n822), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n641), .A2(new_n413), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n654), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(G169gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(new_n524), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n814), .A2(new_n642), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n414), .A3(new_n344), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT122), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n525), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n911), .B2(new_n916), .ZN(G1348gat));
  INV_X1    g716(.A(G176gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n910), .A2(new_n918), .A3(new_n639), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n685), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n918), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(KEYINPUT123), .A3(new_n918), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(G1349gat));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n910), .B2(new_n566), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n906), .A2(KEYINPUT125), .A3(new_n683), .A4(new_n909), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(G183gat), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n248), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n930), .A3(new_n566), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT60), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n910), .B2(new_n608), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n915), .A2(new_n217), .A3(new_n609), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n860), .A2(new_n413), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n913), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n525), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n697), .A2(new_n908), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT126), .Z(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(new_n890), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n525), .A2(G197gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n685), .A3(new_n890), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G204gat), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n944), .A2(G204gat), .A3(new_n639), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n953), .B(new_n956), .C1(new_n958), .C2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n300), .A3(new_n683), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n947), .A2(new_n683), .A3(new_n890), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n945), .B2(new_n609), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n608), .A2(new_n301), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n949), .B2(new_n967), .ZN(G1355gat));
endmodule


