

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587;

  XNOR2_X1 U321 ( .A(KEYINPUT108), .B(KEYINPUT46), .ZN(n361) );
  XNOR2_X1 U322 ( .A(n362), .B(n361), .ZN(n381) );
  XOR2_X1 U323 ( .A(G99GAT), .B(G85GAT), .Z(n385) );
  XNOR2_X1 U324 ( .A(n385), .B(n297), .ZN(n298) );
  XNOR2_X1 U325 ( .A(n368), .B(n298), .ZN(n301) );
  XNOR2_X1 U326 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U327 ( .A(n393), .B(n392), .ZN(n396) );
  NOR2_X1 U328 ( .A1(n518), .A2(n411), .ZN(n452) );
  INV_X1 U329 ( .A(KEYINPUT124), .ZN(n447) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(n585) );
  NOR2_X1 U331 ( .A1(n531), .A2(n455), .ZN(n572) );
  NOR2_X1 U332 ( .A1(n508), .A2(n516), .ZN(n513) );
  XOR2_X1 U333 ( .A(n466), .B(KEYINPUT28), .Z(n530) );
  XNOR2_X1 U334 ( .A(n449), .B(G204GAT), .ZN(n450) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(G1353GAT) );
  XOR2_X1 U336 ( .A(G92GAT), .B(G64GAT), .Z(n290) );
  XNOR2_X1 U337 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n289) );
  XNOR2_X1 U338 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U339 ( .A(G176GAT), .B(n291), .Z(n341) );
  XOR2_X1 U340 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n293) );
  XNOR2_X1 U341 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U343 ( .A(n341), .B(n294), .Z(n308) );
  XOR2_X1 U344 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n296) );
  XNOR2_X1 U345 ( .A(G71GAT), .B(G57GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n368) );
  AND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n297) );
  INV_X1 U348 ( .A(n301), .ZN(n299) );
  NAND2_X1 U349 ( .A1(n299), .A2(KEYINPUT72), .ZN(n303) );
  INV_X1 U350 ( .A(KEYINPUT72), .ZN(n300) );
  NAND2_X1 U351 ( .A1(n301), .A2(n300), .ZN(n302) );
  NAND2_X1 U352 ( .A1(n303), .A2(n302), .ZN(n306) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(G78GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n304), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U355 ( .A(n427), .B(KEYINPUT71), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n405) );
  INV_X1 U358 ( .A(n405), .ZN(n460) );
  XOR2_X1 U359 ( .A(G127GAT), .B(G134GAT), .Z(n310) );
  XNOR2_X1 U360 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U362 ( .A(G113GAT), .B(n311), .Z(n444) );
  XOR2_X1 U363 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n313) );
  NAND2_X1 U364 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT92), .B(n314), .ZN(n329) );
  XOR2_X1 U367 ( .A(KEYINPUT1), .B(G57GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G148GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U370 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n327) );
  XOR2_X1 U374 ( .A(G85GAT), .B(G155GAT), .Z(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n322) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n428) );
  XNOR2_X1 U378 ( .A(n428), .B(G162GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n325), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U383 ( .A(n444), .B(n330), .Z(n471) );
  INV_X1 U384 ( .A(n471), .ZN(n518) );
  XOR2_X1 U385 ( .A(KEYINPUT76), .B(G218GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n394) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U389 ( .A(G197GAT), .B(KEYINPUT21), .Z(n413) );
  XNOR2_X1 U390 ( .A(n333), .B(n413), .ZN(n334) );
  XOR2_X1 U391 ( .A(n394), .B(n334), .Z(n339) );
  XOR2_X1 U392 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n336) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n433) );
  XNOR2_X1 U395 ( .A(G8GAT), .B(G183GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n337), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U397 ( .A(n433), .B(n369), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n521) );
  INV_X1 U400 ( .A(n521), .ZN(n464) );
  XOR2_X1 U401 ( .A(n405), .B(KEYINPUT41), .Z(n566) );
  XOR2_X1 U402 ( .A(KEYINPUT67), .B(KEYINPUT8), .Z(n343) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(G29GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U405 ( .A(KEYINPUT7), .B(n344), .Z(n398) );
  XOR2_X1 U406 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n346) );
  XNOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT29), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G197GAT), .Z(n348) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G50GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U412 ( .A(G8GAT), .B(G113GAT), .Z(n350) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(G141GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U415 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G1GAT), .Z(n376) );
  XOR2_X1 U417 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n354) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n376), .B(n355), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U422 ( .A(n359), .B(n358), .Z(n360) );
  XOR2_X1 U423 ( .A(n398), .B(n360), .Z(n562) );
  NAND2_X1 U424 ( .A1(n566), .A2(n562), .ZN(n362) );
  XOR2_X1 U425 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n364) );
  XNOR2_X1 U426 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n380) );
  XOR2_X1 U428 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n366) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U431 ( .A(n367), .B(KEYINPUT81), .Z(n371) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U434 ( .A(KEYINPUT79), .B(G64GAT), .Z(n373) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G78GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U437 ( .A(n375), .B(n374), .Z(n378) );
  XOR2_X1 U438 ( .A(G22GAT), .B(G155GAT), .Z(n412) );
  XNOR2_X1 U439 ( .A(n376), .B(n412), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n582) );
  XOR2_X1 U442 ( .A(KEYINPUT107), .B(n582), .Z(n539) );
  NAND2_X1 U443 ( .A1(n381), .A2(n539), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n382), .B(KEYINPUT109), .ZN(n399) );
  XOR2_X1 U445 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n384) );
  XNOR2_X1 U446 ( .A(G106GAT), .B(G92GAT), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT9), .B(n385), .Z(n387) );
  XOR2_X1 U449 ( .A(G50GAT), .B(G162GAT), .Z(n416) );
  XNOR2_X1 U450 ( .A(G134GAT), .B(n416), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U452 ( .A(n389), .B(n388), .Z(n393) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  INV_X1 U454 ( .A(KEYINPUT75), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n394), .B(KEYINPUT10), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U457 ( .A(n398), .B(n397), .Z(n571) );
  INV_X1 U458 ( .A(n571), .ZN(n559) );
  NAND2_X1 U459 ( .A1(n399), .A2(n559), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT47), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT36), .B(n559), .Z(n584) );
  INV_X1 U462 ( .A(n582), .ZN(n491) );
  NAND2_X1 U463 ( .A1(n584), .A2(n491), .ZN(n402) );
  XOR2_X1 U464 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n403) );
  INV_X1 U466 ( .A(n562), .ZN(n576) );
  NAND2_X1 U467 ( .A1(n403), .A2(n576), .ZN(n404) );
  NOR2_X1 U468 ( .A1(n405), .A2(n404), .ZN(n406) );
  NOR2_X1 U469 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT48), .ZN(n528) );
  NOR2_X1 U471 ( .A1(n464), .A2(n528), .ZN(n410) );
  INV_X1 U472 ( .A(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT22), .B(G218GAT), .Z(n415) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U477 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U478 ( .A(G211GAT), .B(G204GAT), .Z(n419) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U481 ( .A(KEYINPUT23), .B(n420), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n424) );
  XNOR2_X1 U484 ( .A(KEYINPUT87), .B(KEYINPUT89), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n466) );
  XOR2_X1 U489 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U490 ( .A(G71GAT), .B(G176GAT), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n443) );
  XOR2_X1 U492 ( .A(G99GAT), .B(G190GAT), .Z(n435) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U495 ( .A(G183GAT), .B(KEYINPUT85), .Z(n437) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(KEYINPUT83), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n531) );
  INV_X1 U503 ( .A(n531), .ZN(n523) );
  NOR2_X1 U504 ( .A1(n466), .A2(n523), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n446), .B(KEYINPUT26), .ZN(n546) );
  NAND2_X1 U506 ( .A1(n452), .A2(n546), .ZN(n448) );
  INV_X1 U507 ( .A(n585), .ZN(n581) );
  NOR2_X1 U508 ( .A1(n460), .A2(n581), .ZN(n451) );
  XNOR2_X1 U509 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n449) );
  NAND2_X1 U510 ( .A1(n466), .A2(n452), .ZN(n454) );
  INV_X1 U511 ( .A(KEYINPUT55), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  INV_X1 U513 ( .A(n572), .ZN(n456) );
  NOR2_X1 U514 ( .A1(n456), .A2(n539), .ZN(n459) );
  INV_X1 U515 ( .A(G183GAT), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT122), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  NAND2_X1 U518 ( .A1(n562), .A2(n460), .ZN(n494) );
  XNOR2_X1 U519 ( .A(KEYINPUT27), .B(n521), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n463), .A2(n518), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT94), .ZN(n529) );
  NOR2_X1 U522 ( .A1(n529), .A2(n530), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n531), .A2(n462), .ZN(n474) );
  NAND2_X1 U524 ( .A1(n463), .A2(n546), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n531), .A2(n464), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT95), .B(n465), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NAND2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT96), .ZN(n489) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n477) );
  NAND2_X1 U534 ( .A1(n491), .A2(n559), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n489), .A2(n478), .ZN(n508) );
  NOR2_X1 U537 ( .A1(n494), .A2(n508), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(n479), .Z(n487) );
  NAND2_X1 U539 ( .A1(n518), .A2(n487), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n487), .A2(n521), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT98), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U546 ( .A1(n487), .A2(n523), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U548 ( .A(G15GAT), .B(n486), .Z(G1326GAT) );
  NAND2_X1 U549 ( .A1(n487), .A2(n530), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n489), .A2(n584), .ZN(n490) );
  NOR2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(KEYINPUT101), .Z(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n517) );
  NOR2_X1 U555 ( .A1(n517), .A2(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n518), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n521), .A2(n504), .ZN(n500) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U565 ( .A1(n504), .A2(n523), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n530), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT105), .ZN(n507) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(n507), .Z(n510) );
  NAND2_X1 U573 ( .A1(n576), .A2(n566), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n513), .A2(n518), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n521), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n523), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U581 ( .A1(n513), .A2(n530), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n520) );
  NOR2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n525), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n547) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n547), .A2(n532), .ZN(n533) );
  XNOR2_X1 U597 ( .A(KEYINPUT110), .B(n533), .ZN(n542) );
  NOR2_X1 U598 ( .A1(n542), .A2(n576), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT111), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XNOR2_X1 U601 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n537) );
  INV_X1 U602 ( .A(n566), .ZN(n550) );
  NOR2_X1 U603 ( .A1(n550), .A2(n542), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n542), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(n540), .Z(n541) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n542), .A2(n559), .ZN(n544) );
  XNOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT113), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n576), .A2(n558), .ZN(n548) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n548), .Z(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT114), .B(n549), .ZN(G1344GAT) );
  NOR2_X1 U617 ( .A1(n558), .A2(n550), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT52), .Z(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n582), .A2(n558), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT118), .B(n560), .Z(n561) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n572), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n565) );
  XNOR2_X1 U632 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n570) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(n575), .ZN(G1351GAT) );
  NOR2_X1 U642 ( .A1(n576), .A2(n581), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

