//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n464), .B2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(new_n460), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n477), .A2(new_n462), .A3(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n469), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT68), .Z(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n484));
  OAI211_X1 g059(.A(G2105), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n468), .A2(G136), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(new_n461), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n471), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n491), .A2(G138), .A3(new_n460), .A4(new_n463), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n460), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n473), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(G114), .B2(new_n460), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n485), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n467), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n496), .A2(new_n497), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(new_n503), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT71), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(G543), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G62), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT72), .Z(new_n533));
  AOI21_X1  g108(.A(new_n521), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G166));
  AND2_X1   g110(.A1(new_n520), .A2(new_n525), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  INV_X1    g112(.A(new_n529), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n537), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n521), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n526), .A2(new_n547), .B1(new_n548), .B2(new_n529), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n521), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n526), .A2(new_n553), .B1(new_n554), .B2(new_n529), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  AND3_X1   g137(.A1(new_n518), .A2(G65), .A3(new_n519), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT75), .Z(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n520), .A2(G91), .A3(new_n525), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT74), .B1(new_n568), .B2(KEYINPUT73), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(KEYINPUT74), .B2(new_n568), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n570), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n522), .A2(new_n524), .A3(G53), .A4(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(new_n569), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n566), .A2(new_n567), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  XNOR2_X1  g151(.A(G171), .B(new_n576), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  XNOR2_X1  g153(.A(G166), .B(KEYINPUT77), .ZN(G303));
  NAND2_X1  g154(.A1(new_n536), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n538), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n521), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n538), .A2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n536), .A2(G86), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n521), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n526), .A2(new_n592), .B1(new_n593), .B2(new_n529), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n591), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n521), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n526), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n538), .A2(G54), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT10), .B1(new_n526), .B2(new_n599), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n598), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT78), .Z(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G321));
  XOR2_X1   g180(.A(G321), .B(KEYINPUT79), .Z(G284));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(new_n556), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n604), .A2(new_n611), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n620));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  INV_X1    g196(.A(G123), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n620), .B1(new_n467), .B2(new_n621), .C1(new_n622), .C2(new_n485), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT15), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2435), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT81), .Z(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(KEYINPUT17), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n652), .C1(new_n648), .C2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n649), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n647), .A3(new_n651), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n648), .A2(new_n653), .A3(new_n651), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n673), .C2(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT84), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT21), .Z(new_n678));
  XOR2_X1   g253(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n678), .B(new_n683), .Z(G229));
  OR2_X1    g259(.A1(G6), .A2(G16), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(G305), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT32), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n686), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n686), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(G1971), .Z(new_n697));
  NAND3_X1  g272(.A1(new_n689), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT34), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n686), .A2(G24), .ZN(new_n700));
  INV_X1    g275(.A(G290), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n686), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  OR2_X1    g281(.A1(G95), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n708));
  INV_X1    g283(.A(G131), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n467), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G119), .B2(new_n486), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n706), .B1(new_n711), .B2(new_n705), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  NAND3_X1  g289(.A1(new_n699), .A2(new_n704), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT36), .ZN(new_n716));
  NAND2_X1  g291(.A1(G168), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G16), .B2(G21), .ZN(new_n718));
  INV_X1    g293(.A(G1966), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n604), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1348), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(G160), .A2(G29), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n726), .B2(new_n730), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  OR2_X1    g308(.A1(G29), .A2(G32), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n486), .A2(G129), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G141), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n737), .B(new_n738), .C1(new_n467), .C2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n705), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n733), .A2(G2084), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G33), .ZN(new_n746));
  OR3_X1    g321(.A1(new_n745), .A2(G29), .A3(G33), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n460), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT89), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n468), .A2(G139), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT88), .Z(new_n752));
  NAND3_X1  g327(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND3_X1  g329(.A1(new_n750), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n746), .B(new_n747), .C1(new_n755), .C2(new_n705), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n744), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n705), .A2(G26), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n762));
  INV_X1    g337(.A(G140), .ZN(new_n763));
  INV_X1    g338(.A(G128), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n762), .B1(new_n467), .B2(new_n763), .C1(new_n764), .C2(new_n485), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n760), .B1(new_n765), .B2(G29), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n760), .B(new_n766), .S(KEYINPUT28), .Z(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n733), .C2(G2084), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G11), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n718), .B2(new_n719), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G35), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G162), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n774), .B1(new_n742), .B2(new_n743), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n771), .B(new_n782), .C1(new_n772), .C2(G11), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n686), .A2(KEYINPUT23), .A3(G20), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n786));
  INV_X1    g361(.A(G20), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G299), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n788), .C1(new_n789), .C2(new_n686), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(G28), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(G28), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n794), .A2(new_n795), .A3(new_n705), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n796), .C1(new_n779), .C2(new_n778), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n686), .A2(G19), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n556), .B2(new_n686), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT85), .B(G1341), .Z(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT86), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n799), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G27), .A2(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G164), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2078), .ZN(new_n805));
  NOR2_X1   g380(.A1(G171), .A2(new_n686), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G5), .B2(new_n686), .ZN(new_n807));
  INV_X1    g382(.A(G1961), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n807), .A2(new_n808), .B1(new_n705), .B2(new_n625), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n797), .A2(new_n802), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  AND4_X1   g385(.A1(new_n759), .A2(new_n783), .A3(new_n784), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n716), .A2(new_n721), .A3(new_n725), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n807), .A2(new_n808), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(G311));
  OR2_X1    g389(.A1(new_n812), .A2(new_n813), .ZN(G150));
  AOI22_X1  g390(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n521), .ZN(new_n817));
  INV_X1    g392(.A(G93), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n526), .A2(new_n818), .B1(new_n819), .B2(new_n529), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n604), .A2(G559), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(new_n556), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n613), .A2(new_n821), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n827), .B(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n824), .B1(new_n832), .B2(G860), .ZN(G145));
  INV_X1    g408(.A(new_n711), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n486), .A2(G130), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n468), .A2(G142), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n460), .A2(G118), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n834), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n625), .B(G160), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G162), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(new_n741), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n755), .B(new_n765), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(new_n501), .C1(new_n485), .C2(new_n502), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n491), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n846), .B1(new_n849), .B2(new_n501), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n508), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n628), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n845), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n843), .A2(new_n741), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n844), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n844), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n841), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n844), .A2(new_n854), .ZN(new_n859));
  INV_X1    g434(.A(new_n853), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(new_n840), .A3(new_n855), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  XNOR2_X1  g441(.A(G166), .B(G288), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G290), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(G305), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(G305), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(KEYINPUT99), .A2(KEYINPUT42), .ZN(new_n872));
  NAND2_X1  g447(.A1(KEYINPUT99), .A2(KEYINPUT42), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n830), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n616), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n615), .A2(new_n830), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n603), .A2(new_n789), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n603), .A2(new_n789), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT41), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n882), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT98), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n878), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n868), .A2(G305), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n868), .A2(G305), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n873), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n876), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n886), .B(new_n889), .C1(new_n875), .C2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G868), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n821), .A2(G868), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n866), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g477(.A(KEYINPUT100), .B(new_n900), .C1(new_n898), .C2(G868), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(G295));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n901), .ZN(G331));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NAND2_X1  g481(.A1(G301), .A2(G168), .ZN(new_n907));
  NAND2_X1  g482(.A1(G286), .A2(G171), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n830), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n830), .A3(new_n908), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n910), .B(new_n911), .C1(new_n884), .C2(new_n883), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n887), .B1(new_n913), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n863), .B1(new_n915), .B2(new_n871), .ZN(new_n916));
  INV_X1    g491(.A(new_n888), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n909), .B2(new_n913), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n893), .B1(new_n918), .B2(new_n912), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n906), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n915), .A2(new_n924), .A3(new_n871), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n912), .B(new_n914), .C1(new_n893), .C2(KEYINPUT101), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n863), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n927), .A2(new_n906), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT102), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n927), .B2(KEYINPUT43), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n933), .B2(new_n930), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(G397));
  NOR2_X1   g512(.A1(new_n834), .A2(new_n713), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n741), .B(G1996), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n765), .B(new_n768), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G160), .A2(G40), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n851), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n942), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G2067), .B2(new_n765), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  INV_X1    g526(.A(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT127), .Z(new_n954));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n955));
  OR3_X1    g530(.A1(new_n948), .A2(new_n955), .A3(G1996), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n741), .B2(new_n941), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n948), .B2(G1996), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n701), .A2(new_n703), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n948), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT48), .ZN(new_n963));
  INV_X1    g538(.A(new_n938), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n834), .A2(new_n713), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n942), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n952), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n954), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n503), .A2(KEYINPUT97), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n847), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n971), .B2(new_n508), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n973));
  AND4_X1   g548(.A1(new_n969), .A2(new_n851), .A3(KEYINPUT45), .A4(new_n946), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n504), .A2(new_n511), .A3(new_n946), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n943), .B1(new_n976), .B2(new_n945), .ZN(new_n977));
  AOI21_X1  g552(.A(G1971), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n944), .C1(KEYINPUT50), .C2(new_n976), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G2090), .ZN(new_n981));
  OAI21_X1  g556(.A(G8), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G303), .A2(G8), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT106), .B(KEYINPUT55), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(G303), .A2(G8), .A3(new_n984), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n943), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n972), .A2(KEYINPUT105), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT105), .B1(new_n972), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G2090), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n988), .B(G8), .C1(new_n978), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G305), .A2(KEYINPUT49), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n585), .A2(new_n999), .A3(new_n586), .A4(new_n587), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n585), .A2(KEYINPUT107), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G1981), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n947), .A2(new_n943), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n998), .A2(G1981), .A3(new_n1002), .A4(new_n1000), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G288), .A2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1005), .A2(new_n1011), .A3(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1012), .B(new_n1013), .C1(G1976), .C2(new_n691), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n990), .A2(new_n997), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n504), .A2(new_n511), .A3(KEYINPUT45), .A4(new_n946), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n943), .B1(new_n947), .B2(new_n945), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n719), .ZN(new_n1025));
  INV_X1    g600(.A(G2084), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n991), .C1(new_n993), .C2(new_n994), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(G168), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT51), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1006), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G286), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1028), .A2(KEYINPUT122), .A3(new_n1033), .A4(G8), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1018), .B1(new_n1035), .B2(KEYINPUT62), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  INV_X1    g612(.A(G2078), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n977), .B(new_n1038), .C1(new_n973), .C2(new_n974), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1037), .A2(new_n1039), .B1(new_n995), .B2(new_n808), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1022), .A2(KEYINPUT53), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1041), .A2(new_n1038), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G301), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1030), .A2(new_n1045), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1036), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1009), .A2(new_n1010), .A3(new_n691), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G1981), .B2(G305), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1007), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n997), .B2(new_n1016), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1031), .A2(G168), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1018), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n978), .B2(new_n996), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n989), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1053), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n997), .A4(new_n1017), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1051), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1047), .A2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT114), .B(G1996), .Z(new_n1061));
  OAI211_X1 g636(.A(new_n977), .B(new_n1061), .C1(new_n973), .C2(new_n974), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n947), .B2(new_n943), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n556), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1065), .B2(new_n556), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT115), .B(new_n613), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n1071), .B2(KEYINPUT59), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  NOR4_X1   g649(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1067), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1067), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n980), .A2(new_n791), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT112), .B(KEYINPUT56), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(G2072), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n977), .B(new_n1083), .C1(new_n973), .C2(new_n974), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n574), .A2(KEYINPUT110), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n571), .A2(new_n1087), .A3(new_n573), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n566), .A3(new_n567), .A4(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT109), .B(KEYINPUT57), .Z(new_n1090));
  AND3_X1   g665(.A1(new_n1089), .A2(KEYINPUT111), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT111), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(G299), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g671(.A(KEYINPUT113), .B1(new_n1093), .B2(G299), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1085), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1081), .A2(new_n1084), .A3(new_n1094), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT61), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1080), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1099), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n995), .A2(new_n724), .B1(new_n768), .B2(new_n1005), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT121), .B(new_n603), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n603), .A2(KEYINPUT121), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n603), .A2(KEYINPUT121), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1094), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1085), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1099), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1085), .B2(new_n1115), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1104), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1077), .A2(new_n1079), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1105), .A2(new_n603), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1098), .B1(new_n1099), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n975), .A2(KEYINPUT53), .A3(new_n1038), .A4(new_n1022), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1040), .A2(G301), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(KEYINPUT54), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT123), .B(new_n1127), .C1(new_n1043), .C2(G301), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1018), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1040), .A2(new_n1126), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  INV_X1    g710(.A(G171), .ZN(new_n1136));
  AOI211_X1 g711(.A(KEYINPUT124), .B(new_n1136), .C1(new_n1040), .C2(new_n1126), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1039), .A2(new_n1037), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n995), .A2(new_n808), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1042), .A2(new_n1139), .A3(new_n1140), .A4(G301), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT54), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1132), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1135), .A2(new_n1137), .A3(KEYINPUT125), .A4(new_n1142), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1131), .B(new_n1035), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1060), .B1(new_n1125), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n966), .B1(G1986), .B2(G290), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n948), .B1(new_n1149), .B2(new_n961), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n968), .B1(new_n1148), .B2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g726(.A1(new_n864), .A2(new_n645), .A3(new_n662), .ZN(new_n1153));
  INV_X1    g727(.A(G229), .ZN(new_n1154));
  AND4_X1   g728(.A1(G319), .A2(new_n934), .A3(new_n1153), .A4(new_n1154), .ZN(G308));
  NAND4_X1  g729(.A1(new_n934), .A2(new_n1153), .A3(G319), .A4(new_n1154), .ZN(G225));
endmodule


