//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G77), .B2(G244), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(G50), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n224), .B(new_n228), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n210), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT69), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n230), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G238), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G97), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G226), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G232), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G1698), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n258), .B(new_n261), .C1(new_n268), .C2(new_n255), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n216), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n265), .A2(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n262), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n255), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(new_n258), .A4(new_n261), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n270), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G200), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n253), .A2(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n286), .A2(G77), .B1(new_n287), .B2(G50), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n217), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n229), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n292), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n256), .A2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G68), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT11), .B1(new_n290), .B2(new_n292), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n289), .A2(G1), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n297), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n270), .A2(G190), .A3(new_n283), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n285), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n284), .A2(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n270), .A2(G179), .A3(new_n283), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n284), .A2(new_n308), .A3(G169), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n302), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT17), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n316));
  OAI211_X1 g0116(.A(G223), .B(new_n271), .C1(new_n316), .C2(new_n253), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT76), .B1(new_n317), .B2(G1698), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n253), .A2(new_n207), .ZN(new_n319));
  INV_X1    g0119(.A(new_n271), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n272), .A2(KEYINPUT74), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n320), .B1(new_n324), .B2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n216), .A2(new_n275), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n325), .A2(new_n328), .A3(G223), .A4(new_n275), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n318), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n280), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n255), .A2(new_n257), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n261), .B1(new_n332), .B2(new_n265), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(G200), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(G190), .B(new_n333), .C1(new_n330), .C2(new_n280), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n321), .A2(new_n323), .A3(new_n253), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n273), .ZN(new_n340));
  INV_X1    g0140(.A(G20), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(G20), .B2(new_n267), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n217), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G58), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n217), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(new_n202), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n338), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n253), .B1(new_n321), .B2(new_n323), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n344), .B(new_n341), .C1(new_n353), .C2(new_n320), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n272), .A2(KEYINPUT74), .ZN(new_n356));
  OAI21_X1  g0156(.A(G33), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(G20), .B1(new_n357), .B2(new_n271), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT7), .ZN(new_n359));
  OAI211_X1 g0159(.A(G68), .B(new_n354), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT16), .A3(new_n350), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n352), .A2(new_n361), .A3(new_n292), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n292), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(KEYINPUT70), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n295), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT8), .B(G58), .Z(new_n369));
  MUX2_X1   g0169(.A(new_n363), .B(new_n368), .S(new_n369), .Z(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n315), .B1(new_n337), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n331), .A2(new_n373), .A3(new_n334), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n333), .B1(new_n330), .B2(new_n280), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(G200), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n376), .A2(KEYINPUT17), .A3(new_n362), .A4(new_n370), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n331), .A2(G179), .A3(new_n334), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n375), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT18), .B1(new_n382), .B2(new_n371), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n382), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n379), .B1(new_n383), .B2(new_n384), .C1(KEYINPUT73), .C2(new_n313), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G223), .A2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n275), .A2(G222), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n267), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n280), .C1(G77), .C2(new_n267), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(new_n261), .C1(new_n216), .C2(new_n332), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n366), .A2(new_n367), .A3(G50), .A4(new_n295), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n364), .A2(new_n215), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n369), .A2(new_n286), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n395));
  INV_X1    g0195(.A(G150), .ZN(new_n396));
  INV_X1    g0196(.A(new_n287), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n394), .B(new_n395), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n292), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n393), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n390), .A2(new_n381), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n391), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n392), .A2(new_n399), .A3(KEYINPUT9), .A4(new_n393), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT71), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n390), .A2(new_n373), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT9), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n400), .A2(new_n406), .B1(G200), .B2(new_n390), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT10), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT10), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n404), .A2(new_n410), .A3(new_n405), .A4(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n402), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n274), .B1(G232), .B2(new_n275), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n218), .B2(new_n275), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n280), .C1(G107), .C2(new_n267), .ZN(new_n415));
  INV_X1    g0215(.A(new_n332), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G244), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n261), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n381), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT15), .B(G87), .Z(new_n420));
  AOI22_X1  g0220(.A1(new_n287), .A2(new_n369), .B1(new_n420), .B2(new_n286), .ZN(new_n421));
  INV_X1    g0221(.A(G77), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n341), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n292), .B1(new_n422), .B2(new_n364), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n294), .A2(G77), .A3(new_n295), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n419), .B(new_n426), .C1(G179), .C2(new_n418), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(G200), .B2(new_n418), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n373), .B2(new_n418), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n412), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT72), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n412), .A2(KEYINPUT72), .A3(new_n427), .A4(new_n429), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n314), .B(new_n385), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT5), .B(G41), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n256), .A2(G45), .A3(G274), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n256), .A3(G45), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n255), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n442), .B2(G264), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G294), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n208), .A2(new_n275), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n271), .B(new_n445), .C1(new_n316), .C2(new_n253), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n275), .A2(G257), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n280), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n443), .A2(new_n449), .A3(G179), .ZN(new_n450));
  INV_X1    g0250(.A(new_n439), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n441), .B2(new_n210), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT84), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(new_n454), .A3(new_n280), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n450), .B1(new_n456), .B2(new_n381), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n341), .B(new_n271), .C1(new_n316), .C2(new_n253), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT22), .B1(new_n458), .B2(new_n207), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n274), .A2(new_n460), .A3(G20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n286), .A2(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n209), .A2(G20), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT23), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT24), .ZN(new_n469));
  INV_X1    g0269(.A(new_n464), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n459), .B2(new_n462), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n467), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n294), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n256), .A2(G33), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n365), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n209), .ZN(new_n477));
  XOR2_X1   g0277(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n478));
  NOR2_X1   g0278(.A1(new_n363), .A2(G107), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n457), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n472), .B1(new_n471), .B2(new_n467), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n357), .A2(new_n341), .A3(G87), .A4(new_n271), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(KEYINPUT22), .B1(new_n461), .B2(G87), .ZN(new_n486));
  NOR4_X1   g0286(.A1(new_n486), .A2(KEYINPUT24), .A3(new_n470), .A4(new_n466), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n292), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n448), .A2(new_n454), .A3(new_n280), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n454), .B1(new_n448), .B2(new_n280), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n373), .B(new_n443), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n443), .A2(new_n449), .ZN(new_n492));
  INV_X1    g0292(.A(G200), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n488), .A2(new_n495), .A3(new_n481), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n483), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n210), .A2(G1698), .ZN(new_n498));
  OR2_X1    g0298(.A1(G257), .A2(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n357), .A2(new_n271), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n274), .A2(G303), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n280), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n440), .A2(G270), .A3(new_n255), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n451), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G179), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n364), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n294), .A2(G116), .A3(new_n363), .A4(new_n475), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n291), .A2(new_n229), .B1(G20), .B2(new_n508), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  INV_X1    g0312(.A(G97), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n341), .C1(G33), .C2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n511), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n509), .B(new_n510), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n506), .A2(new_n507), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n506), .A2(G169), .A3(new_n517), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT21), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n504), .B1(new_n502), .B2(new_n280), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n381), .B1(new_n522), .B2(new_n451), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT21), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n517), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n519), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n503), .A2(G190), .A3(new_n451), .A4(new_n505), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n518), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n493), .B1(new_n522), .B2(new_n451), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n506), .A2(G200), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(KEYINPUT81), .A3(new_n518), .A4(new_n528), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n267), .B2(G250), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n512), .C1(new_n538), .C2(new_n275), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT4), .B1(new_n325), .B2(G244), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n280), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n442), .A2(G257), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n541), .A2(new_n373), .A3(new_n451), .A4(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n541), .A2(new_n451), .A3(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(G200), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n364), .A2(new_n513), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n476), .B2(new_n513), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT77), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n343), .B1(new_n341), .B2(new_n274), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(new_n339), .B2(new_n273), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(KEYINPUT7), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n209), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  XOR2_X1   g0353(.A(G97), .B(G107), .Z(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(KEYINPUT6), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G20), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n359), .B(G20), .C1(new_n339), .C2(new_n273), .ZN(new_n557));
  OAI211_X1 g0357(.A(KEYINPUT77), .B(G107), .C1(new_n557), .C2(new_n549), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n287), .A2(G77), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n552), .A2(new_n556), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n547), .B1(new_n560), .B2(new_n292), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n545), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n541), .A2(new_n451), .A3(new_n542), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n381), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n541), .A2(new_n507), .A3(new_n451), .A4(new_n542), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n561), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n365), .A2(new_n420), .A3(new_n475), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n458), .A2(new_n217), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n262), .A2(KEYINPUT19), .A3(G20), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G87), .A2(G97), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n209), .B1(new_n262), .B2(new_n341), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n292), .B1(new_n570), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n420), .A2(new_n363), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT79), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n325), .A2(new_n341), .A3(G68), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n294), .B1(new_n582), .B2(new_n576), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n583), .A2(new_n584), .A3(new_n579), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n569), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n275), .A2(G244), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G238), .A2(G1698), .ZN(new_n588));
  NOR4_X1   g0388(.A1(new_n353), .A2(new_n320), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n253), .A2(new_n508), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n280), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n438), .B(KEYINPUT78), .ZN(new_n592));
  INV_X1    g0392(.A(G45), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n255), .B(G250), .C1(G1), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n381), .ZN(new_n596));
  INV_X1    g0396(.A(new_n594), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n357), .B(new_n271), .C1(G238), .C2(G1698), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n598), .A2(new_n587), .B1(new_n253), .B2(new_n508), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n599), .B2(new_n280), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n507), .A3(new_n592), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n586), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n476), .A2(new_n207), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n580), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n584), .B1(new_n583), .B2(new_n579), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n595), .A2(G200), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n600), .A2(KEYINPUT80), .A3(G190), .A4(new_n592), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n591), .A2(G190), .A3(new_n592), .A4(new_n594), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT80), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n497), .A2(new_n535), .A3(new_n568), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n435), .A2(new_n615), .ZN(G372));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n384), .B2(new_n383), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT18), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n362), .A2(new_n370), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n381), .B1(new_n331), .B2(new_n334), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n507), .B(new_n333), .C1(new_n330), .C2(new_n280), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n619), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n382), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(KEYINPUT87), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n308), .B1(new_n284), .B2(G169), .ZN(new_n628));
  AOI211_X1 g0428(.A(KEYINPUT14), .B(new_n381), .C1(new_n270), .C2(new_n283), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n302), .B1(new_n630), .B2(new_n307), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n427), .A2(new_n304), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n379), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n409), .A2(new_n411), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n402), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n602), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n483), .A2(new_n526), .A3(KEYINPUT85), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n568), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n604), .A2(new_n605), .ZN(new_n640));
  INV_X1    g0440(.A(new_n603), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n607), .A3(new_n641), .A4(new_n609), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n496), .A2(new_n602), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n483), .A2(new_n526), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n637), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n560), .A2(new_n292), .ZN(new_n648));
  INV_X1    g0448(.A(new_n547), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n564), .A2(new_n565), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n602), .A2(new_n650), .A3(new_n651), .A4(new_n642), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n614), .A2(KEYINPUT26), .A3(new_n567), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n652), .A2(KEYINPUT86), .A3(new_n653), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n647), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n636), .B1(new_n435), .B2(new_n661), .ZN(G369));
  XNOR2_X1  g0462(.A(KEYINPUT91), .B(G330), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n299), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n256), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n517), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n535), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT89), .B1(new_n526), .B2(new_n673), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n526), .A2(KEYINPUT89), .A3(new_n673), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT90), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n674), .A2(KEYINPUT90), .A3(new_n675), .A4(new_n676), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n664), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n671), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n488), .B2(new_n481), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT92), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT92), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n497), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n443), .B1(new_n489), .B2(new_n490), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G169), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n488), .A2(new_n481), .B1(new_n688), .B2(new_n450), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n671), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n681), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n526), .A2(new_n671), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n684), .A2(new_n497), .A3(new_n685), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n682), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n225), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G1), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n573), .A2(new_n209), .A3(new_n508), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n702), .A2(new_n703), .B1(new_n232), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n450), .A2(new_n595), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n544), .A3(new_n522), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n506), .A2(new_n595), .A3(new_n507), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n563), .A2(new_n492), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n671), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n714), .B(KEYINPUT31), .C1(new_n615), .C2(new_n671), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n671), .C1(new_n709), .C2(new_n713), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n664), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n660), .A2(new_n682), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n496), .A2(new_n602), .A3(new_n642), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n568), .A3(new_n644), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n614), .A2(new_n653), .A3(new_n567), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n637), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .A3(new_n682), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n719), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n705), .B1(new_n729), .B2(G1), .ZN(G364));
  AOI21_X1  g0530(.A(new_n702), .B1(G45), .B2(new_n665), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n373), .A2(G20), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G159), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT32), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(G190), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n513), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n341), .A2(new_n373), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n507), .A2(new_n493), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n493), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n746), .A2(new_n215), .B1(new_n748), .B2(new_n207), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n507), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n733), .A2(new_n745), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n267), .B1(new_n751), .B2(new_n347), .C1(new_n752), .C2(new_n217), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n733), .A2(new_n747), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n749), .B(new_n753), .C1(G107), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n733), .A2(new_n750), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n743), .B(new_n756), .C1(new_n422), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n746), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n748), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  INV_X1    g0563(.A(G329), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n754), .A2(new_n763), .B1(new_n735), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n757), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n762), .B(new_n765), .C1(G311), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n274), .B1(new_n751), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n752), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n767), .B(new_n772), .C1(new_n773), .C2(new_n741), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n758), .B1(new_n760), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n229), .B1(G20), .B2(new_n381), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n299), .A2(new_n253), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT95), .Z(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n776), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n267), .A2(G355), .A3(new_n225), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n325), .A2(new_n699), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n248), .B2(new_n593), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n233), .A2(G45), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n782), .B1(G116), .B2(new_n225), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n775), .A2(new_n776), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n679), .A2(new_n680), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n780), .B(KEYINPUT96), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n731), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n681), .A2(new_n731), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n788), .B2(new_n663), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n426), .A2(new_n671), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n429), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n427), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n427), .A2(new_n671), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n652), .A2(KEYINPUT86), .A3(new_n653), .ZN(new_n801));
  AOI21_X1  g0601(.A(KEYINPUT86), .B1(new_n652), .B2(new_n653), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n651), .A2(new_n650), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n613), .A2(new_n803), .A3(new_n653), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n519), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n524), .B1(new_n523), .B2(new_n517), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n255), .B1(new_n500), .B2(new_n501), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(new_n439), .A3(new_n504), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n809), .A2(KEYINPUT21), .A3(new_n518), .A4(new_n381), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n806), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n645), .B1(new_n689), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n812), .A2(new_n723), .A3(new_n568), .A4(new_n638), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n602), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n682), .B(new_n800), .C1(new_n805), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OR3_X1    g0616(.A1(new_n719), .A2(new_n816), .A3(KEYINPUT99), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n719), .B1(new_n816), .B2(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(new_n720), .A3(new_n799), .ZN(new_n820));
  INV_X1    g0620(.A(new_n731), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n671), .B1(new_n647), .B2(new_n659), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n817), .B(new_n818), .C1(new_n822), .C2(new_n800), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n754), .A2(new_n207), .ZN(new_n825));
  INV_X1    g0625(.A(new_n751), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G294), .B2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n209), .B2(new_n748), .C1(new_n761), .C2(new_n746), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n274), .B1(new_n757), .B2(new_n508), .C1(new_n763), .C2(new_n752), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n828), .A2(new_n742), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n735), .ZN(new_n832));
  INV_X1    g0632(.A(new_n325), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G58), .B2(new_n740), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n754), .A2(new_n217), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G132), .B2(new_n736), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n215), .C2(new_n748), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT98), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n770), .A2(G150), .B1(new_n826), .B2(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G159), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n746), .C1(new_n843), .C2(new_n757), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n839), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n832), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n776), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n777), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n849), .A2(new_n776), .B1(new_n422), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n731), .B(new_n853), .C1(new_n800), .C2(new_n779), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n824), .A2(new_n854), .ZN(G384));
  INV_X1    g0655(.A(new_n669), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n371), .B1(new_n382), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n362), .B(new_n370), .C1(new_n335), .C2(new_n336), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n361), .A2(new_n292), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n360), .B2(new_n350), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n370), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n382), .B2(new_n856), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n859), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n860), .B1(new_n865), .B2(new_n858), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n863), .A2(new_n856), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n384), .A2(new_n383), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n378), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n717), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n545), .A2(new_n561), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n803), .A2(new_n483), .A3(new_n496), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n526), .A2(new_n534), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n876), .A2(new_n613), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n716), .B1(new_n878), .B2(new_n682), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(new_n714), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  INV_X1    g0681(.A(new_n304), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n311), .A2(new_n671), .ZN(new_n883));
  INV_X1    g0683(.A(new_n307), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n628), .A2(new_n629), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n882), .B(new_n883), .C1(new_n885), .C2(new_n302), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n310), .A2(new_n311), .A3(new_n671), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n881), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT102), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT102), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n312), .A2(new_n883), .B1(new_n631), .B2(new_n671), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n892), .B(new_n889), .C1(new_n893), .C2(new_n881), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n891), .A2(new_n894), .A3(new_n800), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n873), .A2(new_n880), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n860), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n858), .B1(new_n857), .B2(new_n859), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n859), .A2(new_n315), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT17), .B1(new_n620), .B2(new_n376), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT103), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT103), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n372), .A2(new_n377), .A3(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n905), .A2(new_n618), .A3(new_n626), .A4(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n620), .A2(new_n669), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n872), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(new_n880), .A3(KEYINPUT40), .A4(new_n895), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n435), .A2(new_n718), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n663), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n722), .A2(new_n434), .A3(new_n728), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n917), .A2(new_n636), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n911), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n631), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n671), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n870), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n920), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n891), .A2(new_n894), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n815), .B2(new_n798), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n873), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n627), .A2(new_n856), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n918), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n916), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n256), .B2(new_n665), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n232), .A2(new_n422), .A3(new_n348), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n201), .A2(new_n217), .ZN(new_n936));
  OAI211_X1 g0736(.A(G1), .B(new_n299), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(G20), .B(new_n230), .C1(new_n555), .C2(KEYINPUT35), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n508), .B(new_n938), .C1(KEYINPUT35), .C2(new_n555), .ZN(new_n939));
  XNOR2_X1  g0739(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n937), .A3(new_n941), .ZN(G367));
  AOI21_X1  g0742(.A(new_n274), .B1(new_n826), .B2(G150), .ZN(new_n943));
  INV_X1    g0743(.A(new_n201), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(new_n217), .B2(new_n741), .C1(new_n944), .C2(new_n757), .ZN(new_n945));
  INV_X1    g0745(.A(new_n746), .ZN(new_n946));
  INV_X1    g0746(.A(new_n748), .ZN(new_n947));
  AOI22_X1  g0747(.A1(G143), .A2(new_n946), .B1(new_n947), .B2(G58), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(new_n422), .B2(new_n754), .C1(new_n842), .C2(new_n735), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n945), .B(new_n949), .C1(G159), .C2(new_n770), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n770), .A2(G294), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n754), .A2(new_n513), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G317), .B2(new_n736), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n763), .B2(new_n757), .C1(new_n761), .C2(new_n751), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n947), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n748), .B2(new_n508), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n209), .C2(new_n741), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n833), .B1(new_n831), .B2(new_n746), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n950), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  AOI21_X1  g0762(.A(new_n821), .B1(new_n962), .B2(new_n776), .ZN(new_n963));
  INV_X1    g0763(.A(new_n420), .ZN(new_n964));
  INV_X1    g0764(.A(new_n783), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n781), .B1(new_n225), .B2(new_n964), .C1(new_n244), .C2(new_n965), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n602), .A2(new_n606), .A3(new_n682), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n602), .B(new_n642), .C1(new_n606), .C2(new_n682), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n963), .B(new_n966), .C1(new_n789), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n256), .B1(new_n665), .B2(G45), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n650), .A2(new_n671), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n568), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n567), .A2(new_n671), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n694), .A3(new_n695), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT45), .Z(new_n978));
  INV_X1    g0778(.A(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n696), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n692), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT107), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n982), .A3(new_n692), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n681), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n681), .B2(KEYINPUT108), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n729), .C1(new_n983), .C2(KEYINPUT107), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n729), .B1(new_n986), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n700), .B(KEYINPUT41), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n972), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n568), .A2(new_n689), .A3(new_n973), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n803), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT105), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(KEYINPUT105), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n682), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT42), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n694), .A2(new_n1003), .A3(new_n974), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n694), .B2(new_n974), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n969), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT106), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1008), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(KEYINPUT106), .B(new_n969), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1011));
  OAI211_X1 g0811(.A(KEYINPUT43), .B(new_n1007), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n969), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1007), .A2(new_n1009), .A3(new_n1008), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1012), .B1(KEYINPUT43), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n692), .A2(new_n979), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1012), .B(new_n1018), .C1(KEYINPUT43), .C2(new_n1016), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n970), .B1(new_n997), .B2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n369), .A2(new_n215), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n703), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(G68), .A2(G77), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n593), .A4(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n783), .B(new_n1028), .C1(new_n240), .C2(new_n593), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n267), .A2(new_n703), .A3(new_n225), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G107), .C2(new_n225), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n781), .B1(new_n1031), .B2(KEYINPUT109), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT109), .B2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n766), .A2(G303), .B1(new_n826), .B2(G317), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(KEYINPUT110), .B1(G311), .B2(new_n770), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(KEYINPUT110), .B2(new_n1034), .C1(new_n768), .C2(new_n746), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n763), .B2(new_n741), .C1(new_n773), .C2(new_n748), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT49), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n325), .B1(G116), .B2(new_n755), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n759), .C2(new_n735), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n757), .A2(new_n217), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n748), .A2(new_n422), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1043), .B(new_n952), .C1(new_n369), .C2(new_n770), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n735), .A2(new_n396), .B1(new_n751), .B2(new_n215), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G159), .B2(new_n946), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n741), .A2(new_n964), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n833), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1041), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1033), .B1(new_n1050), .B2(new_n776), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n731), .C1(new_n691), .C2(new_n789), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n990), .A2(new_n992), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n729), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n1053), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n700), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1053), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1052), .B1(new_n971), .B2(new_n1053), .C1(new_n1056), .C2(new_n1057), .ZN(G393));
  NAND2_X1  g0858(.A1(new_n978), .A2(new_n982), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n692), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT107), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1063), .A2(new_n1057), .A3(new_n985), .A4(new_n984), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT111), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1065), .A3(new_n985), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n978), .A2(new_n982), .A3(KEYINPUT111), .A4(new_n692), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1064), .B(new_n700), .C1(new_n1068), .C2(new_n1057), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n781), .B1(new_n513), .B2(new_n225), .C1(new_n251), .C2(new_n965), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n976), .A2(G20), .A3(new_n779), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n267), .B1(new_n755), .B2(G107), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n763), .B2(new_n748), .C1(new_n768), .C2(new_n735), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT112), .Z(new_n1074));
  NAND2_X1  g0874(.A1(new_n766), .A2(G294), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n946), .A2(G317), .B1(new_n826), .B2(G311), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n770), .A2(G303), .B1(G116), .B2(new_n740), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n741), .A2(new_n422), .ZN(new_n1080));
  INV_X1    g0880(.A(G143), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n752), .A2(new_n944), .B1(new_n735), .B2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(G68), .C2(new_n947), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n825), .B(new_n833), .C1(new_n369), .C2(new_n766), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n746), .A2(new_n396), .B1(new_n751), .B2(new_n843), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n850), .B1(new_n1079), .B2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1071), .A2(new_n821), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1068), .A2(new_n972), .B1(new_n1070), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1069), .A2(new_n1090), .ZN(G390));
  NAND3_X1  g0891(.A1(new_n434), .A2(G330), .A3(new_n880), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n917), .A2(new_n1092), .A3(new_n636), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n927), .ZN(new_n1094));
  INV_X1    g0894(.A(G330), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n718), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(new_n800), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n727), .A2(new_n682), .A3(new_n797), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n798), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n715), .A2(new_n663), .A3(new_n717), .A4(new_n800), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n927), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n798), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n822), .B2(new_n800), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n718), .A2(new_n1095), .A3(new_n799), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1094), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n927), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1093), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT38), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n909), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n372), .A2(new_n906), .A3(new_n377), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n906), .B1(new_n372), .B2(new_n377), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1111), .B1(new_n627), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1110), .B1(new_n1115), .B2(new_n902), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT39), .B1(new_n1116), .B2(new_n872), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n873), .A2(new_n919), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1117), .A2(new_n1118), .B1(new_n928), .B2(new_n922), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT113), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n922), .B1(new_n1116), .B2(new_n872), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n927), .B1(new_n798), .B2(new_n1098), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n922), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n911), .A2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1126), .A2(KEYINPUT113), .A3(new_n1122), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1106), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1119), .B(new_n1101), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1109), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(new_n701), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1129), .A2(new_n1109), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n971), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT114), .ZN(new_n1136));
  INV_X1    g0936(.A(G132), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n751), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n267), .B1(new_n746), .B2(new_n1139), .C1(new_n842), .C2(new_n752), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G159), .C2(new_n740), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n748), .A2(new_n396), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT53), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  AOI22_X1  g0944(.A1(new_n755), .A2(new_n201), .B1(new_n766), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G125), .B2(new_n736), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n766), .A2(G97), .B1(new_n826), .B2(G116), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n209), .B2(new_n752), .C1(new_n763), .C2(new_n746), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n274), .B1(new_n748), .B2(new_n207), .C1(new_n735), .C2(new_n773), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1149), .A2(new_n835), .A3(new_n1080), .A4(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n776), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n369), .B2(new_n851), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n920), .A2(new_n925), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n821), .B(new_n1153), .C1(new_n1154), .C2(new_n778), .ZN(new_n1155));
  OR3_X1    g0955(.A1(new_n1135), .A2(new_n1136), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1136), .B1(new_n1135), .B2(new_n1155), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1134), .A2(new_n1156), .A3(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1093), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1121), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT113), .B1(new_n1126), .B2(new_n1122), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1125), .B1(new_n1104), .B2(new_n927), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1161), .A2(new_n1162), .B1(new_n1163), .B2(new_n1154), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1106), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1130), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1102), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1108), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1160), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n891), .A2(new_n894), .A3(new_n800), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n924), .A2(new_n718), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n912), .B(G330), .C1(new_n1172), .C2(new_n897), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n400), .A2(new_n856), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT56), .Z(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT55), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n412), .A2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(KEYINPUT55), .B(new_n402), .C1(new_n409), .C2(new_n411), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1176), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1173), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT118), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n1180), .A3(KEYINPUT118), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n899), .A2(new_n1189), .A3(G330), .A4(new_n912), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n931), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1184), .A2(new_n931), .A3(new_n1190), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1159), .B1(new_n1170), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1184), .A2(new_n931), .A3(new_n1190), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n931), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(KEYINPUT57), .C1(new_n1131), .C2(new_n1160), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1200), .A3(new_n700), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1186), .A2(new_n1188), .A3(new_n778), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n741), .A2(new_n396), .B1(new_n751), .B2(new_n1139), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n766), .A2(G137), .B1(new_n947), .B2(new_n1144), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1137), .B2(new_n752), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G125), .C2(new_n946), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G41), .B1(new_n736), .B2(G124), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G33), .B1(new_n755), .B2(G159), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n833), .B(new_n254), .C1(new_n422), .C2(new_n748), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT115), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n754), .A2(new_n347), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n752), .A2(new_n513), .B1(new_n735), .B2(new_n763), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n420), .C2(new_n766), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n741), .A2(new_n217), .B1(new_n746), .B2(new_n508), .ZN(new_n1216));
  OR3_X1    g1016(.A1(new_n751), .A2(KEYINPUT116), .A3(new_n209), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT116), .B1(new_n751), .B2(new_n209), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1212), .A2(new_n1215), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1220), .B(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G41), .B1(new_n316), .B2(G33), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1210), .B(new_n1222), .C1(G50), .C2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1224), .A2(new_n776), .B1(new_n944), .B2(new_n852), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1202), .A2(new_n731), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1199), .B2(new_n972), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1201), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT119), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1201), .A2(KEYINPUT119), .A3(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(G375));
  NAND3_X1  g1032(.A1(new_n1160), .A2(new_n1168), .A3(new_n1167), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n996), .A3(new_n1109), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1094), .A2(new_n777), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n766), .A2(G107), .B1(new_n826), .B2(G283), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n513), .B2(new_n748), .C1(new_n773), .C2(new_n746), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n752), .A2(new_n508), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n274), .B1(new_n735), .B2(new_n761), .C1(new_n422), .C2(new_n754), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1237), .A2(new_n1047), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1213), .B1(G159), .B2(new_n947), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n842), .B2(new_n751), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n770), .A2(new_n1144), .B1(new_n946), .B2(G132), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n396), .B2(new_n757), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n735), .A2(new_n1139), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n325), .B1(new_n741), .B2(new_n215), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n776), .B1(new_n1240), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(G68), .B2(new_n851), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1235), .A2(new_n821), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1169), .B2(new_n972), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1234), .A2(new_n1251), .ZN(G381));
  AND3_X1   g1052(.A1(new_n1201), .A2(KEYINPUT119), .A3(new_n1227), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT119), .B1(new_n1201), .B2(new_n1227), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT121), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT121), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1230), .A2(new_n1256), .A3(new_n1231), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT120), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n996), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1064), .B2(new_n729), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1020), .B(new_n1021), .C1(new_n1260), .C2(new_n972), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1069), .A2(new_n1090), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n970), .A4(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G381), .A2(G384), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1258), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(G387), .A2(G390), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(KEYINPUT120), .A3(new_n1265), .A4(new_n1263), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1134), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1255), .A2(new_n1257), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT122), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1272), .B(new_n1273), .ZN(G407));
  NAND4_X1  g1074(.A1(new_n1255), .A2(new_n1257), .A3(new_n670), .A4(new_n1271), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1275), .A2(G213), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT123), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(KEYINPUT123), .A3(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G409));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(G393), .A2(G396), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(new_n1263), .ZN(new_n1287));
  OR3_X1    g1087(.A1(new_n1285), .A2(new_n1268), .A3(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1285), .B2(new_n1268), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n670), .A2(G213), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1199), .B1(new_n1131), .B2(new_n1160), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1227), .B1(new_n1292), .B2(new_n1259), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1271), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G378), .A2(new_n1227), .A3(new_n1201), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1291), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1233), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1160), .A2(new_n1167), .A3(KEYINPUT60), .A4(new_n1168), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n700), .A3(new_n1109), .A4(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G384), .B1(new_n1300), .B2(new_n1251), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(G384), .A3(new_n1251), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1296), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(KEYINPUT125), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1296), .B2(new_n1305), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1307), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1291), .B(new_n1304), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1291), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1304), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1302), .A2(new_n1303), .A3(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1319), .A2(new_n1296), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1313), .A2(new_n1314), .A3(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1290), .B1(new_n1311), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT63), .B1(new_n1319), .B2(new_n1296), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1306), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1290), .B1(new_n1312), .B2(KEYINPUT63), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1324), .A2(KEYINPUT124), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT124), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1322), .B1(new_n1326), .B2(new_n1327), .ZN(G405));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1329), .B(new_n1271), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G378), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1295), .A2(KEYINPUT126), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1305), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1290), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1330), .B(new_n1304), .C1(new_n1331), .C2(new_n1332), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1290), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1334), .A2(KEYINPUT127), .A3(new_n1335), .A4(new_n1336), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1339), .A2(new_n1341), .A3(new_n1342), .ZN(G402));
endmodule


