//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n203), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n220), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NOR2_X1   g0043(.A1(G20), .A2(G33), .ZN(new_n244));
  AOI22_X1  g0044(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n202), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n208), .A2(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n245), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n216), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n201), .ZN(new_n258));
  INV_X1    g0058(.A(new_n254), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G1), .B2(new_n208), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n255), .B(new_n258), .C1(new_n201), .C2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT9), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G222), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G223), .A2(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n267), .B(new_n268), .C1(G77), .C2(new_n263), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT64), .B(G45), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n207), .B(G274), .C1(new_n270), .C2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n269), .A2(new_n271), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G200), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT10), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n279), .A2(new_n280), .B1(KEYINPUT69), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(G190), .B2(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n262), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n261), .B(new_n288), .C1(G169), .C2(new_n279), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT66), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT15), .B(G87), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT67), .B1(new_n291), .B2(new_n251), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n208), .A2(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n292), .B1(new_n208), .B2(new_n293), .C1(new_n295), .C2(new_n246), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n291), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n254), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n257), .A2(new_n293), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n259), .A2(new_n300), .A3(new_n256), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT68), .B1(new_n257), .B2(new_n254), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G1), .B2(new_n208), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n298), .B(new_n299), .C1(new_n293), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G238), .A2(G1698), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n263), .B(new_n306), .C1(new_n220), .C2(G1698), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n268), .C1(G107), .C2(new_n263), .ZN(new_n308));
  INV_X1    g0108(.A(G244), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(new_n271), .C1(new_n309), .C2(new_n275), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(G179), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(G200), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n310), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(new_n305), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n290), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n203), .A2(G20), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n320), .B1(new_n251), .B2(new_n293), .C1(new_n201), .C2(new_n295), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n254), .ZN(new_n322));
  XOR2_X1   g0122(.A(new_n322), .B(KEYINPUT71), .Z(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n304), .A2(KEYINPUT12), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT12), .ZN(new_n328));
  INV_X1    g0128(.A(G13), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n328), .A2(new_n329), .A3(G1), .ZN(new_n330));
  INV_X1    g0130(.A(new_n320), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(new_n328), .B2(new_n256), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n221), .B1(new_n275), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n334), .B2(new_n275), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n220), .A2(G1698), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G226), .B2(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT3), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n337), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n268), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n336), .A2(new_n271), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT13), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(KEYINPUT13), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n287), .B2(new_n349), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n349), .B2(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n333), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n280), .B1(new_n347), .B2(new_n348), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n349), .A2(new_n316), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n333), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n286), .A2(new_n319), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(G223), .A2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G226), .B2(new_n264), .ZN(new_n360));
  INV_X1    g0160(.A(G87), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n360), .A2(new_n343), .B1(new_n294), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n362), .A2(new_n268), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n271), .B1(new_n220), .B2(new_n275), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n312), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n207), .A2(G274), .ZN(new_n367));
  INV_X1    g0167(.A(new_n270), .ZN(new_n368));
  INV_X1    g0168(.A(G41), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n275), .A2(new_n220), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(G179), .B1(new_n362), .B2(new_n268), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n271), .B(KEYINPUT75), .C1(new_n220), .C2(new_n275), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n295), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n244), .A2(KEYINPUT73), .A3(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n202), .A2(new_n203), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n263), .B2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT72), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(KEYINPUT72), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n294), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n342), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT74), .B1(new_n294), .B2(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT7), .B(new_n208), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n203), .B1(new_n397), .B2(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(new_n385), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n399), .A3(new_n254), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n250), .A2(new_n260), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n250), .B2(new_n257), .ZN(new_n402));
  AOI211_X1 g0202(.A(KEYINPUT18), .B(new_n376), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n402), .ZN(new_n405));
  INV_X1    g0205(.A(new_n376), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  INV_X1    g0209(.A(new_n402), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n343), .B2(new_n208), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n203), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT72), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n385), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n259), .B1(new_n415), .B2(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n410), .B1(new_n416), .B2(new_n399), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n362), .A2(new_n268), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n372), .A2(new_n374), .A3(new_n316), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n280), .B1(new_n363), .B2(new_n364), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n409), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  AND4_X1   g0222(.A1(new_n409), .A2(new_n400), .A3(new_n421), .A4(new_n402), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n408), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n358), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n340), .A2(new_n342), .A3(G244), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT4), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(G1698), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n263), .A2(G244), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G283), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n263), .A2(G250), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n264), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n268), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n207), .A2(G45), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(G41), .ZN(new_n438));
  INV_X1    g0238(.A(G274), .ZN(new_n439));
  INV_X1    g0239(.A(new_n216), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n272), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n369), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n437), .B2(G41), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n437), .A2(G41), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n442), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G257), .A3(new_n273), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n435), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n435), .A2(new_n454), .A3(new_n451), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(G200), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n435), .A2(KEYINPUT78), .A3(new_n451), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(G190), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n397), .B2(new_n388), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n244), .A2(G77), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n464), .A2(new_n465), .A3(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(G97), .B(G107), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n463), .B1(new_n468), .B2(new_n208), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n254), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n256), .A2(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n207), .A2(G33), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n259), .A2(new_n256), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n456), .A2(new_n460), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n435), .A2(KEYINPUT78), .A3(new_n451), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT78), .B1(new_n435), .B2(new_n451), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n312), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n435), .A2(new_n451), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n287), .B1(new_n470), .B2(new_n475), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n309), .A2(G1698), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G238), .B2(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n487), .A2(new_n343), .B1(new_n294), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n268), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT79), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n436), .A2(G250), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n268), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n273), .A2(KEYINPUT79), .A3(G250), .A4(new_n436), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n441), .A2(new_n447), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n490), .A2(new_n495), .A3(G190), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n489), .A2(new_n268), .B1(new_n441), .B2(new_n447), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(KEYINPUT82), .A3(G190), .A4(new_n495), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n291), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n256), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n340), .A2(new_n342), .A3(new_n208), .A4(G68), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT81), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n208), .B1(new_n337), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n361), .A2(new_n465), .A3(new_n461), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(KEYINPUT80), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n511), .A2(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n504), .B1(new_n515), .B2(new_n254), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n500), .A2(new_n495), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(G200), .B1(G87), .B2(new_n474), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n502), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n312), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n500), .A2(new_n287), .A3(new_n495), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT81), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n505), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n511), .A2(new_n512), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n513), .A2(new_n507), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n510), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n254), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n504), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n473), .A2(new_n291), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n520), .B(new_n521), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n519), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n264), .A2(G257), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G264), .A2(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n340), .A2(new_n342), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n268), .C1(G303), .C2(new_n263), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n449), .A2(G270), .A3(new_n273), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n445), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n257), .A2(new_n488), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n253), .A2(new_n216), .B1(G20), .B2(new_n488), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n431), .B(new_n208), .C1(G33), .C2(new_n465), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n540), .A2(KEYINPUT20), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT20), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n488), .B1(new_n207), .B2(G33), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n301), .A2(new_n302), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G169), .B(new_n538), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT21), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n536), .A2(new_n445), .A3(new_n537), .A4(G179), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n301), .A2(new_n302), .A3(new_n545), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n539), .C1(new_n543), .C2(new_n542), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n547), .A2(new_n548), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n538), .A2(G200), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n316), .C2(new_n538), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n549), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n532), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n257), .A2(new_n461), .ZN(new_n560));
  NOR2_X1   g0360(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n560), .B2(new_n561), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n562), .A2(new_n564), .B1(new_n474), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n567), .A2(new_n208), .A3(G107), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT23), .B1(new_n461), .B2(G20), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n340), .A2(new_n342), .A3(new_n208), .A4(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n263), .A2(new_n573), .A3(new_n208), .A4(G87), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n254), .B1(new_n575), .B2(KEYINPUT24), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n577), .B(new_n570), .C1(new_n572), .C2(new_n574), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n565), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n263), .A2(G250), .A3(new_n264), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n263), .A2(G257), .A3(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n268), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n449), .A2(G264), .A3(new_n273), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n445), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n587), .A2(new_n316), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(G200), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n580), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n585), .A2(new_n287), .A3(new_n445), .A4(new_n586), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n312), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n579), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT84), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n559), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n425), .A2(new_n485), .A3(new_n598), .ZN(G372));
  INV_X1    g0399(.A(new_n290), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n352), .A2(new_n353), .ZN(new_n601));
  INV_X1    g0401(.A(new_n314), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n333), .B1(new_n357), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n422), .A2(new_n423), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n408), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n600), .B1(new_n605), .B2(new_n286), .ZN(new_n606));
  INV_X1    g0406(.A(new_n425), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G238), .A2(G1698), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n309), .B2(G1698), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n263), .B1(G33), .B2(G116), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n496), .B1(new_n610), .B2(new_n273), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n493), .A2(new_n494), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n474), .A2(G87), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT85), .B1(new_n615), .B2(new_n529), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n518), .A2(new_n516), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n618), .A3(new_n502), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n435), .A2(new_n287), .A3(new_n451), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n476), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n458), .A2(new_n459), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n312), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n619), .A2(new_n623), .A3(new_n624), .A4(new_n531), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT26), .B1(new_n532), .B2(new_n484), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n531), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT86), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT86), .A4(new_n531), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n594), .A2(new_n549), .A3(new_n554), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n478), .A2(new_n631), .A3(new_n484), .A4(new_n590), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n619), .A2(new_n531), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n606), .B1(new_n607), .B2(new_n637), .ZN(G369));
  NAND2_X1  g0438(.A1(new_n597), .A2(new_n595), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n329), .A2(G1), .A3(G20), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT87), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT27), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G213), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n579), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT88), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n549), .A2(new_n554), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n594), .B2(new_n647), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n594), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n647), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n647), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n555), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n558), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n662), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n652), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n656), .A2(new_n668), .ZN(G399));
  OR2_X1    g0469(.A1(new_n509), .A2(G116), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT89), .Z(new_n671));
  INV_X1    g0471(.A(new_n211), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n671), .A2(new_n207), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n215), .B2(new_n673), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT90), .Z(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n585), .A2(new_n586), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n679), .A2(new_n517), .A3(new_n550), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n458), .A3(new_n459), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n680), .A2(new_n458), .A3(KEYINPUT30), .A4(new_n459), .ZN(new_n684));
  AOI21_X1  g0484(.A(G179), .B1(new_n500), .B2(new_n495), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n452), .A2(new_n685), .A3(new_n587), .A4(new_n538), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n687), .A2(KEYINPUT91), .A3(KEYINPUT31), .A4(new_n647), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n647), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n692), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n532), .A2(new_n558), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n639), .A2(new_n485), .A3(new_n700), .A4(new_n661), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT93), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n598), .A2(new_n703), .A3(new_n485), .A4(new_n661), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n678), .B1(new_n699), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n634), .B1(new_n628), .B2(new_n627), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n647), .B1(new_n707), .B2(new_n630), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n619), .A2(new_n623), .A3(KEYINPUT26), .A4(new_n531), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n624), .B1(new_n532), .B2(new_n484), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n531), .B1(new_n632), .B2(new_n633), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n661), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n706), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n677), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR2_X1   g0516(.A1(new_n208), .A2(new_n287), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n316), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G322), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n208), .A2(G179), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n316), .A3(G200), .ZN(new_n726));
  INV_X1    g0526(.A(G283), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n343), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n718), .A2(new_n287), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(G294), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n717), .A2(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n316), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(G190), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT33), .B(G317), .ZN(new_n735));
  AOI22_X1  g0535(.A1(G326), .A2(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G303), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n725), .A2(G190), .A3(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G190), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n717), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n737), .A2(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n725), .A2(new_n739), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(G329), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n724), .A2(new_n731), .A3(new_n736), .A4(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n722), .B(KEYINPUT96), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n202), .ZN(new_n748));
  INV_X1    g0548(.A(new_n734), .ZN(new_n749));
  INV_X1    g0549(.A(new_n730), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n749), .A2(new_n203), .B1(new_n750), .B2(new_n465), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(G50), .B2(new_n733), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n743), .A2(new_n378), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n726), .A2(new_n461), .B1(new_n738), .B2(new_n361), .ZN(new_n755));
  INV_X1    g0555(.A(new_n740), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n343), .B(new_n755), .C1(G77), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n752), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n746), .B1(new_n748), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n216), .B1(G20), .B2(new_n312), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n329), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n207), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n673), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n211), .A2(G355), .A3(new_n263), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n672), .A2(new_n263), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n214), .B2(new_n270), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n239), .A2(new_n446), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n767), .B1(G116), .B2(new_n211), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n760), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n766), .B1(new_n771), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n761), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT97), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n665), .B2(new_n775), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n665), .A2(G330), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n666), .A2(new_n766), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(G396));
  NOR2_X1   g0585(.A1(new_n760), .A2(new_n772), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n766), .B1(new_n293), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n305), .A2(new_n311), .A3(new_n313), .A4(new_n647), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n305), .A2(new_n647), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n318), .A2(new_n314), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n722), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n726), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n461), .B2(new_n738), .C1(new_n741), .C2(new_n743), .ZN(new_n797));
  INV_X1    g0597(.A(new_n733), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n749), .A2(new_n727), .B1(new_n798), .B2(new_n737), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n343), .B1(new_n740), .B2(new_n488), .C1(new_n750), .C2(new_n465), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n794), .A2(new_n797), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT98), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n750), .A2(new_n202), .ZN(new_n803));
  INV_X1    g0603(.A(new_n738), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n804), .A2(G50), .B1(new_n744), .B2(G132), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n805), .B(new_n263), .C1(new_n203), .C2(new_n726), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n734), .A2(G150), .B1(new_n756), .B2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n798), .ZN(new_n809));
  INV_X1    g0609(.A(new_n747), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(G143), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n803), .B(new_n806), .C1(new_n811), .C2(KEYINPUT34), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n787), .B1(new_n792), .B2(new_n773), .C1(new_n814), .C2(new_n776), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n708), .B(new_n792), .ZN(new_n816));
  INV_X1    g0616(.A(new_n706), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT100), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n766), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n815), .B1(new_n819), .B2(new_n821), .ZN(G384));
  INV_X1    g0622(.A(new_n468), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT35), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(KEYINPUT35), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n824), .A2(G116), .A3(new_n217), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT36), .Z(new_n827));
  NAND2_X1  g0627(.A1(new_n201), .A2(G68), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT101), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n215), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n207), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n601), .A2(new_n333), .A3(new_n647), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n333), .A2(new_n647), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n354), .A2(new_n357), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n636), .A2(new_n661), .A3(new_n792), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n314), .A2(new_n647), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n417), .B1(new_n376), .B2(new_n645), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n400), .A2(new_n421), .A3(new_n402), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n416), .B1(KEYINPUT16), .B2(new_n415), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n402), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n406), .ZN(new_n849));
  INV_X1    g0649(.A(new_n645), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n851), .A3(new_n843), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n852), .B2(KEYINPUT37), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n417), .A2(new_n409), .A3(new_n421), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n843), .A2(KEYINPUT17), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n851), .B1(new_n408), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n853), .B2(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n841), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n408), .B2(new_n850), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n601), .A2(new_n333), .A3(new_n661), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n860), .B2(new_n861), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT105), .B1(new_n422), .B2(new_n423), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n854), .A2(new_n855), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n408), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n417), .A2(new_n645), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n417), .A2(KEYINPUT103), .A3(new_n421), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n405), .B1(new_n406), .B2(new_n850), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n843), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n842), .B2(new_n845), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n844), .A4(new_n843), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n872), .A2(KEYINPUT106), .A3(new_n873), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n876), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n889));
  AOI21_X1  g0689(.A(new_n859), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n868), .B1(new_n890), .B2(new_n867), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n864), .B1(new_n866), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n709), .A2(new_n425), .A3(new_n714), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n606), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n893), .B(new_n895), .Z(new_n896));
  NAND2_X1  g0696(.A1(new_n697), .A2(new_n688), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n702), .B2(new_n704), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n792), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n837), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n901), .A3(new_n862), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n872), .A2(KEYINPUT106), .A3(new_n873), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT106), .B1(new_n872), .B2(new_n873), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n889), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n860), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n899), .A4(new_n901), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n607), .B2(new_n898), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n904), .A2(new_n911), .A3(new_n425), .A4(new_n899), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(G330), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n896), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n207), .B2(new_n762), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n896), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n832), .B1(new_n917), .B2(new_n918), .ZN(G367));
  NAND2_X1  g0719(.A1(new_n516), .A2(new_n614), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n647), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n619), .A2(new_n531), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n531), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n478), .B(new_n484), .C1(new_n477), .C2(new_n661), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT107), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n925), .A2(new_n926), .B1(new_n623), .B2(new_n647), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n657), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n647), .B1(new_n931), .B2(new_n484), .ZN(new_n932));
  INV_X1    g0732(.A(new_n654), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n929), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n924), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(KEYINPUT109), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(KEYINPUT43), .B2(new_n923), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n930), .A2(new_n667), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n940), .A2(new_n667), .A3(new_n930), .A4(new_n942), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n655), .B1(new_n927), .B2(new_n928), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT44), .B1(new_n656), .B2(new_n929), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n656), .A2(KEYINPUT44), .A3(new_n929), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n667), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n668), .A3(new_n949), .A4(new_n950), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n933), .A2(KEYINPUT110), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT110), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n654), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n659), .C2(new_n653), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(new_n666), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n715), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n715), .B1(new_n954), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n673), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n945), .B(new_n946), .C1(new_n964), .C2(new_n764), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n778), .B1(new_n211), .B2(new_n291), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n768), .A2(new_n235), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n765), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n723), .A2(G150), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n750), .A2(new_n203), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G159), .B2(new_n734), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n263), .B1(new_n726), .B2(new_n293), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G143), .B2(new_n733), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n740), .A2(new_n201), .B1(new_n743), .B2(new_n808), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G58), .B2(new_n804), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n969), .A2(new_n971), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n810), .A2(G303), .B1(G311), .B2(new_n733), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT111), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n738), .A2(new_n488), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n979), .A2(KEYINPUT46), .B1(new_n730), .B2(G107), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(KEYINPUT46), .B2(new_n979), .C1(new_n793), .C2(new_n749), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT112), .B(G317), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n343), .B1(new_n982), .B2(new_n743), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n465), .A2(new_n726), .B1(new_n740), .B2(new_n727), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n978), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n977), .A2(KEYINPUT111), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n976), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n968), .B1(new_n989), .B2(new_n760), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n775), .B2(new_n923), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT113), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n965), .A2(new_n992), .ZN(G387));
  NOR2_X1   g0793(.A1(new_n959), .A2(new_n715), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n960), .A2(new_n673), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(KEYINPUT117), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(KEYINPUT117), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n959), .A2(new_n764), .ZN(new_n998));
  INV_X1    g0798(.A(new_n768), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n232), .B2(new_n270), .ZN(new_n1000));
  AOI211_X1 g0800(.A(G45), .B(new_n671), .C1(G68), .C2(G77), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT114), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n246), .A2(G50), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT114), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1000), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n671), .A2(new_n211), .A3(new_n263), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G107), .C2(new_n211), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n766), .B1(new_n1010), .B2(new_n778), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n733), .A2(G159), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT115), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n201), .B2(new_n722), .C1(new_n250), .C2(new_n749), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n804), .A2(G77), .ZN(new_n1015));
  INV_X1    g0815(.A(G150), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n203), .B2(new_n740), .C1(new_n1016), .C2(new_n743), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n750), .A2(new_n291), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n263), .B1(new_n726), .B2(new_n465), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n733), .A2(G322), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n734), .A2(G311), .B1(new_n756), .B2(G303), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n747), .C2(new_n982), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n804), .A2(G294), .B1(new_n730), .B2(G283), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT49), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n726), .A2(new_n488), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n263), .B(new_n1030), .C1(G326), .C2(new_n744), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1020), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1011), .B1(new_n1032), .B2(new_n776), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT116), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n660), .B2(new_n774), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n997), .A2(new_n998), .A3(new_n1037), .ZN(G393));
  NAND3_X1  g0838(.A1(new_n952), .A2(new_n764), .A3(new_n953), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n778), .B1(new_n465), .B2(new_n211), .C1(new_n242), .C2(new_n999), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT118), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n766), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n723), .A2(G311), .B1(G317), .B2(new_n733), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  AOI22_X1  g0845(.A1(G294), .A2(new_n756), .B1(new_n744), .B2(G322), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n727), .B2(new_n738), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n343), .B1(new_n461), .B2(new_n726), .C1(new_n749), .C2(new_n737), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G116), .C2(new_n730), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n722), .A2(new_n378), .B1(new_n1016), .B2(new_n798), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  INV_X1    g0852(.A(G143), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n740), .A2(new_n246), .B1(new_n743), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n804), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n750), .A2(new_n293), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n796), .A2(new_n263), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(G50), .C2(new_n734), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1052), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1050), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1043), .B1(new_n1060), .B2(new_n760), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n930), .B2(new_n775), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1039), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n954), .A2(new_n960), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n673), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n954), .A2(new_n960), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  OAI211_X1 g0869(.A(new_n867), .B(new_n860), .C1(new_n908), .C2(new_n909), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n868), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n866), .C2(new_n841), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n699), .A2(new_n705), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1073), .A2(G330), .A3(new_n792), .A4(new_n836), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n661), .B(new_n792), .C1(new_n712), .C2(new_n713), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n840), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n836), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n865), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1078), .A2(new_n890), .A3(KEYINPUT119), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT119), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n866), .B1(new_n1076), .B2(new_n836), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n910), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1072), .B(new_n1074), .C1(new_n1079), .C2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT119), .B1(new_n1078), .B2(new_n890), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n910), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n839), .B1(new_n708), .B2(new_n792), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n865), .B1(new_n1086), .B2(new_n837), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1084), .A2(new_n1085), .B1(new_n891), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n898), .A2(new_n678), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n901), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n425), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n894), .A2(new_n606), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1076), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1074), .A2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n898), .A2(new_n678), .A3(new_n900), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n836), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n702), .A2(new_n704), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n692), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n698), .A2(new_n696), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(G330), .B(new_n792), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n837), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1086), .B1(new_n1105), .B2(new_n1090), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1094), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(KEYINPUT120), .B1(new_n1091), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1086), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1089), .A2(new_n901), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n836), .B1(new_n706), .B2(new_n792), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1074), .B(new_n1095), .C1(new_n836), .C2(new_n1097), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1093), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1072), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1110), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT120), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1083), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1065), .B1(new_n1091), .B2(new_n1107), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1091), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n891), .A2(new_n772), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n250), .A2(new_n786), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n263), .B(new_n1056), .C1(G87), .C2(new_n804), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G107), .A2(new_n734), .B1(new_n733), .B2(G283), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n723), .A2(G116), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n726), .A2(new_n203), .B1(new_n743), .B2(new_n793), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G97), .B2(new_n756), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n733), .A2(G128), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n804), .A2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1131), .B1(new_n750), .B2(new_n378), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n723), .A2(G132), .ZN(new_n1136));
  INV_X1    g0936(.A(G125), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n263), .B1(new_n743), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G50), .B2(new_n795), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1132), .A2(new_n1134), .B1(new_n734), .B2(G137), .ZN(new_n1140));
  XOR2_X1   g0940(.A(KEYINPUT54), .B(G143), .Z(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n756), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1130), .B1(new_n1135), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT123), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n776), .B1(new_n1145), .B2(KEYINPUT123), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n766), .B(new_n1124), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1122), .A2(new_n764), .B1(new_n1123), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1121), .A2(new_n1149), .ZN(G378));
  AOI21_X1  g0950(.A(new_n766), .B1(new_n201), .B2(new_n786), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n503), .A2(new_n756), .B1(new_n744), .B2(G283), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n202), .B2(new_n726), .C1(new_n722), .C2(new_n461), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1015), .A2(new_n369), .A3(new_n343), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n749), .A2(new_n465), .B1(new_n798), .B2(new_n488), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1153), .A2(new_n970), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G50), .B1(new_n294), .B2(new_n369), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n263), .B2(G41), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1142), .A2(new_n804), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT124), .Z(new_n1163));
  OAI22_X1  g0963(.A1(new_n750), .A2(new_n1016), .B1(new_n740), .B2(new_n808), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n798), .A2(new_n1137), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G132), .C2(new_n734), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1163), .B(new_n1166), .C1(new_n1167), .C2(new_n722), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n744), .C2(G124), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n378), .B2(new_n726), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1168), .B2(KEYINPUT59), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1161), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n286), .A2(new_n289), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n261), .A2(new_n850), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1151), .B1(new_n776), .B2(new_n1173), .C1(new_n1178), .C2(new_n773), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n912), .B2(new_n678), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n904), .A3(new_n911), .A4(G330), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1181), .A2(new_n893), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n893), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1179), .B1(new_n1185), .B2(new_n763), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1119), .A2(new_n1094), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1185), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1093), .B1(new_n1108), .B2(new_n1118), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n673), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1187), .B1(new_n1190), .B2(new_n1193), .ZN(G375));
  AOI21_X1  g0994(.A(new_n763), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n837), .A2(new_n772), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n766), .B1(new_n203), .B2(new_n786), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT125), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n263), .B(new_n1018), .C1(G77), .C2(new_n795), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G116), .A2(new_n734), .B1(new_n733), .B2(G294), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n723), .A2(G283), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n740), .A2(new_n461), .B1(new_n743), .B2(new_n737), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G97), .B2(new_n804), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n747), .A2(new_n808), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1142), .A2(new_n734), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n740), .A2(new_n1016), .B1(new_n743), .B2(new_n1167), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G159), .B2(new_n804), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n733), .A2(G132), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n263), .B1(new_n726), .B2(new_n202), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G50), .B2(new_n730), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1205), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1198), .B1(new_n760), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1195), .B1(new_n1196), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1112), .A2(new_n1113), .A3(new_n1093), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1107), .A2(new_n963), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(G381));
  NAND3_X1  g1018(.A1(new_n965), .A2(new_n992), .A3(new_n1068), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1121), .A2(new_n1149), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(G375), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n646), .A2(G213), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1221), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G375), .C2(new_n1227), .ZN(G409));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G378), .B(new_n1187), .C1(new_n1190), .C2(new_n1193), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1191), .A2(new_n962), .A3(new_n1185), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1221), .B1(new_n1186), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1225), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1216), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1216), .A2(new_n1235), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n673), .A3(new_n1107), .A4(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G384), .B1(new_n1238), .B2(new_n1215), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(G384), .A3(new_n1215), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1234), .A2(new_n1242), .A3(KEYINPUT126), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1226), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1242), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1229), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(G393), .B(G396), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1068), .B1(new_n965), .B2(new_n992), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1220), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1219), .A3(new_n1249), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(KEYINPUT61), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1233), .B2(new_n1225), .ZN(new_n1258));
  AOI211_X1 g1058(.A(KEYINPUT127), .B(new_n1226), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1246), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1226), .A2(G2897), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1242), .B(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1234), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1248), .A2(new_n1256), .A3(new_n1261), .A4(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1260), .A2(KEYINPUT62), .A3(new_n1246), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1268), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1255), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1265), .B1(new_n1272), .B2(new_n1273), .ZN(G405));
  XNOR2_X1  g1074(.A(G375), .B(G378), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(new_n1242), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(new_n1255), .ZN(G402));
endmodule


