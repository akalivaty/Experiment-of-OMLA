//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1293, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(new_n219), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G169), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n206), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n251), .A2(G238), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n249), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(new_n254), .A3(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G226), .A2(G1698), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n219), .B2(G1698), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n260), .A2(new_n261), .B1(G33), .B2(G97), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n256), .B(new_n258), .C1(new_n262), .C2(new_n254), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n219), .A2(G1698), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G226), .B2(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n265), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n256), .A4(new_n258), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n248), .B1(new_n264), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT14), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n264), .A2(new_n276), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n278), .A3(G169), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n213), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  XOR2_X1   g0090(.A(new_n290), .B(KEYINPUT70), .Z(new_n291));
  NAND2_X1  g0091(.A1(new_n207), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n292), .A2(new_n293), .B1(new_n207), .B2(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n288), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT11), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n300), .A2(G20), .A3(new_n242), .A4(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n302), .B(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n288), .B1(new_n206), .B2(G20), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(G68), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n297), .A2(new_n298), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n286), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n279), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n279), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n311), .A2(new_n307), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(G50), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n305), .B2(G50), .ZN(new_n318));
  OAI21_X1  g0118(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  INV_X1    g0120(.A(new_n289), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n218), .A2(KEYINPUT8), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT67), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT8), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(G58), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT66), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT66), .B1(new_n325), .B2(G58), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n292), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n322), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n288), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n318), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n336), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n251), .A2(new_n255), .A3(new_n254), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G226), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n271), .A2(new_n293), .ZN(new_n341));
  MUX2_X1   g0141(.A(G222), .B(G223), .S(G1698), .Z(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n273), .C1(new_n271), .C2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n343), .A3(new_n258), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n312), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G200), .B2(new_n344), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(new_n338), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n337), .A2(new_n346), .A3(new_n349), .A4(new_n338), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n344), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n280), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT68), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n335), .B1(G169), .B2(new_n353), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT17), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n324), .A2(new_n330), .A3(new_n316), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n305), .B1(new_n324), .B2(new_n330), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n218), .A2(new_n242), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n364), .B2(new_n201), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n289), .A2(G159), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n269), .A2(G33), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n207), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n371), .A2(new_n372), .B1(new_n271), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n368), .B(KEYINPUT16), .C1(new_n374), .C2(new_n242), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n288), .ZN(new_n376));
  INV_X1    g0176(.A(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT73), .B1(new_n269), .B2(G33), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n369), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n269), .A2(KEYINPUT73), .A3(G33), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(G20), .B1(new_n268), .B2(new_n270), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(KEYINPUT7), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT16), .B1(new_n384), .B2(new_n368), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n363), .B1(new_n376), .B2(new_n385), .ZN(new_n386));
  MUX2_X1   g0186(.A(G223), .B(G226), .S(G1698), .Z(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n261), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n273), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n251), .A2(G232), .A3(new_n254), .A4(new_n255), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(G190), .A3(new_n258), .A4(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n387), .A2(new_n261), .B1(G33), .B2(G87), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n258), .B(new_n392), .C1(new_n394), .C2(new_n254), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n360), .B1(new_n386), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n361), .A2(new_n362), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n382), .A2(KEYINPUT7), .B1(new_n261), .B2(new_n377), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n367), .B1(new_n400), .B2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n334), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n371), .A2(new_n372), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(new_n268), .A3(new_n380), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n373), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n242), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n403), .B1(new_n409), .B2(new_n367), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n399), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n391), .A2(G179), .A3(new_n258), .A4(new_n392), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n395), .A2(G169), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT18), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n386), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n393), .A2(new_n396), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n411), .A2(new_n419), .A3(KEYINPUT17), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n398), .A2(new_n415), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n261), .A2(G238), .A3(G1698), .ZN(new_n423));
  INV_X1    g0223(.A(G1698), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n261), .A2(G232), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G107), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n423), .B(new_n425), .C1(new_n426), .C2(new_n261), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n273), .ZN(new_n428));
  INV_X1    g0228(.A(G274), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n273), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n339), .A2(G244), .B1(new_n257), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT69), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(new_n431), .A3(KEYINPUT69), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G190), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G20), .A2(G77), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n323), .A2(new_n326), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n438), .B1(new_n439), .B2(new_n292), .C1(new_n440), .C2(new_n321), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(new_n288), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n305), .A2(G77), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G77), .B2(new_n316), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G200), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n437), .B(new_n445), .C1(new_n436), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n436), .B2(new_n280), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n434), .A2(new_n248), .A3(new_n435), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  AND4_X1   g0251(.A1(new_n315), .A2(new_n359), .A3(new_n422), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT88), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT78), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n253), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G264), .A3(new_n254), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n430), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G250), .A2(G1698), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n221), .B2(G1698), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(new_n261), .B1(G33), .B2(G294), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n273), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n464), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n221), .A2(G1698), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n261), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G294), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n471), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n461), .B(new_n463), .C1(new_n468), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n248), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n466), .A2(new_n467), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n273), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(new_n280), .A3(new_n461), .A4(new_n463), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n268), .A2(new_n270), .A3(new_n207), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n261), .A2(new_n207), .A3(G87), .A4(new_n483), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n207), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n426), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(KEYINPUT86), .A3(KEYINPUT24), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT86), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n485), .B2(new_n486), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n498), .A2(KEYINPUT85), .A3(new_n499), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT85), .B1(new_n498), .B2(new_n499), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n334), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n316), .B1(G1), .B2(new_n252), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n288), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n316), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT25), .A3(new_n426), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT25), .B1(new_n509), .B2(new_n426), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n508), .A2(new_n426), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n453), .B(new_n481), .C1(new_n505), .C2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n495), .B2(KEYINPUT24), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n498), .A2(KEYINPUT85), .A3(new_n499), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n496), .A3(new_n517), .A4(new_n500), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n513), .B1(new_n518), .B2(new_n288), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n475), .A2(new_n480), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT88), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n288), .ZN(new_n522));
  INV_X1    g0322(.A(new_n513), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n474), .A2(new_n446), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n479), .A2(new_n312), .A3(new_n461), .A4(new_n463), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n514), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n508), .A2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n316), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n220), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G97), .ZN(new_n535));
  AOI21_X1  g0335(.A(G33), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n207), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT82), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n538), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT74), .B(G97), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(G33), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n288), .B1(new_n207), .B2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT20), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT20), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n548), .B(new_n545), .C1(new_n539), .C2(new_n543), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n532), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n261), .A2(G257), .A3(new_n424), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n261), .A2(G264), .A3(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(G303), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n261), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n273), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n460), .A2(G270), .A3(new_n254), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(G179), .A3(new_n463), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n463), .A2(new_n556), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n273), .B2(new_n554), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n248), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n563), .B2(new_n550), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n562), .A2(new_n446), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n544), .A2(new_n546), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n548), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n544), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(new_n570), .B1(new_n529), .B2(new_n531), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n562), .A2(G190), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n560), .B(KEYINPUT21), .C1(new_n563), .C2(new_n550), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n566), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n439), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n316), .ZN(new_n578));
  INV_X1    g0378(.A(G87), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n506), .A2(new_n579), .A3(new_n288), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n207), .B1(new_n265), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n533), .A2(new_n535), .A3(new_n426), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n582), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n261), .A2(new_n207), .A3(G68), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n581), .B1(new_n542), .B2(new_n292), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n578), .B(new_n580), .C1(new_n591), .C2(new_n288), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G116), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n268), .A2(new_n270), .A3(G238), .A4(new_n424), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n268), .A2(new_n270), .A3(G244), .A4(G1698), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(KEYINPUT79), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n273), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n430), .A2(new_n458), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n254), .B(G250), .C1(G1), .C2(new_n457), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n601), .A3(G190), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT79), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n261), .A2(new_n605), .A3(G244), .A4(G1698), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n606), .A3(new_n593), .A4(new_n594), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n607), .B2(new_n273), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n592), .B(new_n602), .C1(new_n446), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n591), .A2(new_n288), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n507), .A2(new_n577), .ZN(new_n611));
  INV_X1    g0411(.A(new_n578), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n598), .A2(new_n601), .A3(new_n280), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n613), .B(new_n614), .C1(new_n608), .C2(G169), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n609), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n609), .B2(new_n615), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n460), .A2(G257), .A3(new_n254), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n463), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n268), .A2(new_n270), .A3(G244), .A4(new_n424), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT4), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n424), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n537), .A4(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n628), .A2(KEYINPUT77), .A3(new_n273), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT77), .B1(new_n628), .B2(new_n273), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n280), .B(new_n622), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n621), .B1(new_n273), .B2(new_n628), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(G169), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT76), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n372), .A2(new_n371), .B1(new_n407), .B2(new_n373), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n426), .ZN(new_n637));
  OAI211_X1 g0437(.A(KEYINPUT76), .B(G107), .C1(new_n381), .C2(new_n383), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT6), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n220), .A2(KEYINPUT6), .A3(G107), .ZN(new_n640));
  OAI21_X1  g0440(.A(G107), .B1(new_n220), .B2(KEYINPUT6), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(G20), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n289), .A2(G77), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT75), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(KEYINPUT75), .A3(new_n643), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n637), .A2(new_n638), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n288), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n316), .A2(G97), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n507), .B2(G97), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n631), .B(new_n634), .C1(new_n649), .C2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G200), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n652), .B1(new_n648), .B2(new_n288), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n632), .A2(G190), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n619), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n452), .A2(new_n528), .A3(new_n576), .A4(new_n660), .ZN(G372));
  AND2_X1   g0461(.A1(new_n415), .A2(new_n418), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n450), .A2(new_n314), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n309), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n398), .A2(new_n420), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT90), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n352), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n358), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n609), .A2(new_n615), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n653), .A2(new_n527), .A3(new_n658), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n519), .A2(new_n520), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n566), .A2(new_n575), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n631), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n677), .A2(new_n656), .A3(new_n633), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n671), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n615), .B(KEYINPUT89), .Z(new_n681));
  NAND2_X1  g0481(.A1(new_n609), .A2(new_n615), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT81), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n609), .A2(new_n615), .A3(new_n616), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n653), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n680), .B(new_n681), .C1(new_n685), .C2(new_n679), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n452), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n670), .A2(new_n687), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n300), .A2(new_n207), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(G343), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(G343), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n673), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n505), .B2(new_n513), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n514), .A2(new_n521), .A3(new_n701), .A4(new_n527), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT94), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n571), .A2(new_n698), .ZN(new_n707));
  NOR4_X1   g0507(.A1(new_n566), .A2(new_n575), .A3(new_n574), .A4(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n707), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n675), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT92), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n576), .A2(new_n709), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT92), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n563), .A2(new_n550), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT83), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT21), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n564), .A2(new_n565), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n559), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n707), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n712), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT93), .B1(new_n721), .B2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n723), .B(new_n724), .C1(new_n711), .C2(new_n720), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n706), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n698), .B(KEYINPUT95), .Z(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n673), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n528), .A2(KEYINPUT94), .A3(new_n701), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n702), .A2(new_n703), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n718), .A3(new_n698), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n726), .A2(new_n729), .A3(new_n732), .ZN(G399));
  INV_X1    g0533(.A(new_n210), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G41), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G1), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n583), .A2(new_n587), .A3(G116), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(new_n216), .B2(new_n736), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n678), .B(new_n679), .C1(new_n617), .C2(new_n618), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT26), .B1(new_n653), .B2(new_n682), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n681), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n659), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n682), .B1(new_n519), .B2(new_n526), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n514), .A2(new_n521), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n718), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n699), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n728), .B1(new_n686), .B2(new_n676), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n528), .A2(new_n660), .A3(new_n576), .A4(new_n728), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT97), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n562), .A2(G179), .A3(new_n461), .A4(new_n479), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n632), .A2(new_n608), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n628), .A2(new_n273), .ZN(new_n759));
  AND4_X1   g0559(.A1(new_n622), .A2(new_n759), .A3(new_n598), .A4(new_n601), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n479), .A2(new_n461), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n760), .A2(new_n558), .A3(KEYINPUT30), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n562), .A2(G179), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT96), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n608), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n598), .A2(new_n601), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n763), .A2(new_n474), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n654), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n758), .B(new_n762), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n727), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n758), .A2(new_n762), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n763), .A2(new_n474), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n773), .A2(new_n654), .A3(new_n765), .A4(new_n767), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n698), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n754), .B(new_n771), .C1(new_n775), .C2(KEYINPUT31), .ZN(new_n776));
  AOI21_X1  g0576(.A(KEYINPUT31), .B1(new_n770), .B2(new_n699), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n772), .B2(new_n774), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT97), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n753), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n749), .A2(new_n752), .B1(G330), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n740), .B1(new_n782), .B2(G1), .ZN(G364));
  NOR3_X1   g0583(.A1(new_n312), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n207), .ZN(new_n785));
  INV_X1    g0585(.A(G294), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n207), .A2(new_n280), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n785), .A2(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(KEYINPUT99), .B1(G311), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(KEYINPUT99), .B2(new_n791), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT100), .Z(new_n797));
  NOR2_X1   g0597(.A1(new_n207), .A2(G179), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n792), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(G190), .A3(new_n446), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n271), .B1(new_n799), .B2(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n787), .A2(new_n312), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n798), .A2(new_n312), .A3(G200), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n809), .B1(new_n810), .B2(new_n811), .C1(new_n553), .C2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n797), .A2(new_n803), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n785), .ZN(new_n815));
  INV_X1    g0615(.A(new_n812), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(G97), .B1(new_n816), .B2(new_n587), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n240), .B2(new_n788), .C1(new_n426), .C2(new_n811), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n799), .A2(KEYINPUT32), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT32), .B1(new_n799), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n242), .B2(new_n804), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n261), .B1(new_n793), .B2(new_n293), .C1(new_n218), .C2(new_n801), .ZN(new_n823));
  NOR4_X1   g0623(.A1(new_n818), .A2(new_n820), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  OR3_X1    g0624(.A1(new_n814), .A2(KEYINPUT101), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT101), .B1(new_n814), .B2(new_n824), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n213), .B1(G20), .B2(new_n248), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n299), .A2(G20), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n206), .B1(new_n832), .B2(G45), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n735), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n734), .A2(new_n271), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G355), .B1(new_n530), .B2(new_n734), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n734), .A2(new_n261), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(G45), .B2(new_n216), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n246), .A2(new_n457), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(G13), .A2(G33), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(G20), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n830), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n836), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n831), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT102), .Z(new_n849));
  INV_X1    g0649(.A(new_n721), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n845), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n721), .A2(G330), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n722), .A2(new_n725), .A3(new_n852), .A4(new_n835), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NOR2_X1   g0655(.A1(new_n450), .A2(new_n699), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n447), .B1(new_n445), .B2(new_n698), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n450), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n728), .B(new_n858), .C1(new_n686), .C2(new_n676), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n861));
  INV_X1    g0661(.A(new_n858), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n750), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n861), .B(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n781), .A2(G330), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n836), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n830), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n844), .ZN(new_n870));
  INV_X1    g0670(.A(new_n799), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n261), .B1(new_n871), .B2(G311), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n872), .B1(new_n530), .B2(new_n793), .C1(new_n786), .C2(new_n801), .ZN(new_n873));
  INV_X1    g0673(.A(new_n788), .ZN(new_n874));
  INV_X1    g0674(.A(new_n811), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G303), .A2(new_n874), .B1(new_n875), .B2(G87), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n426), .B2(new_n812), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n785), .A2(new_n220), .B1(new_n804), .B2(new_n810), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n261), .B1(new_n799), .B2(new_n880), .C1(new_n240), .C2(new_n812), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n785), .A2(new_n218), .B1(new_n811), .B2(new_n242), .ZN(new_n882));
  INV_X1    g0682(.A(new_n801), .ZN(new_n883));
  XNOR2_X1  g0683(.A(KEYINPUT103), .B(G143), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n883), .A2(new_n884), .B1(new_n794), .B2(G159), .ZN(new_n885));
  INV_X1    g0685(.A(G137), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n885), .B1(new_n886), .B2(new_n788), .C1(new_n320), .C2(new_n804), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT104), .Z(new_n888));
  INV_X1    g0688(.A(KEYINPUT34), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n881), .B(new_n882), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n879), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n835), .B1(G77), .B2(new_n870), .C1(new_n892), .C2(new_n869), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT105), .Z(new_n894));
  NOR2_X1   g0694(.A1(new_n858), .A2(new_n844), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n868), .A2(new_n896), .ZN(G384));
  NAND3_X1  g0697(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT35), .ZN(new_n899));
  OAI211_X1 g0699(.A(G116), .B(new_n214), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  OR3_X1    g0702(.A1(new_n216), .A2(new_n293), .A3(new_n364), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n206), .B(G13), .C1(new_n903), .C2(new_n241), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n279), .A2(G169), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n264), .A2(new_n276), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n906), .A2(KEYINPUT14), .B1(new_n907), .B2(G179), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n282), .A2(new_n283), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT72), .B1(new_n277), .B2(new_n278), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n307), .B(new_n699), .C1(new_n911), .C2(new_n314), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n308), .B(new_n310), .C1(new_n312), .C2(new_n279), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n307), .A2(new_n699), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n913), .B(new_n914), .C1(new_n286), .C2(new_n308), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n856), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n859), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n271), .A2(new_n373), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n242), .B1(new_n404), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n403), .B1(new_n921), .B2(new_n367), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n399), .B1(new_n402), .B2(new_n922), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n386), .A2(new_n397), .B1(new_n923), .B2(new_n692), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n414), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n386), .A2(new_n417), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n386), .A2(new_n693), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT37), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n411), .A2(new_n419), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n923), .A2(new_n692), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n421), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n662), .A2(new_n693), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n919), .B2(new_n938), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT107), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n931), .ZN(new_n949));
  INV_X1    g0749(.A(new_n928), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n421), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT38), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT39), .B1(new_n954), .B2(new_n937), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n932), .A2(KEYINPUT38), .A3(new_n934), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n956), .A2(new_n935), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n309), .A2(new_n698), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n943), .A2(new_n946), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n749), .A2(new_n452), .A3(new_n752), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n670), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n963), .B(new_n965), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n777), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n753), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n916), .A2(new_n858), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n948), .A2(new_n931), .B1(new_n421), .B2(new_n950), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n937), .B1(KEYINPUT38), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT40), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n916), .A2(new_n858), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n753), .B2(new_n968), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT40), .B1(new_n936), .B2(new_n937), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n452), .A3(new_n969), .ZN(new_n980));
  AOI22_X1  g0780(.A1(KEYINPUT40), .A2(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n981));
  INV_X1    g0781(.A(new_n452), .ZN(new_n982));
  INV_X1    g0782(.A(new_n969), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n984), .A3(G330), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n966), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n206), .B2(new_n832), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n966), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n905), .B1(new_n987), .B2(new_n988), .ZN(G367));
  OAI21_X1  g0789(.A(new_n744), .B1(new_n656), .B2(new_n728), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n678), .A2(new_n727), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n718), .A2(new_n698), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n992), .A2(new_n730), .A3(new_n731), .A4(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n746), .A2(new_n658), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n727), .B1(new_n997), .B2(new_n653), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n995), .B2(KEYINPUT42), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n592), .A2(new_n698), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n671), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(KEYINPUT108), .B(new_n1001), .C1(new_n681), .C2(new_n1000), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n996), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT43), .B2(new_n1005), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT43), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n996), .A2(new_n999), .A3(new_n1008), .A4(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n992), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n726), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1010), .B(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n735), .B(new_n1014), .Z(new_n1015));
  OAI211_X1 g0815(.A(new_n700), .B(new_n993), .C1(new_n704), .C2(new_n705), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n732), .B(new_n1016), .C1(new_n722), .C2(new_n725), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n708), .A2(new_n710), .A3(KEYINPUT92), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n713), .B1(new_n712), .B2(new_n719), .ZN(new_n1019));
  OAI21_X1  g0819(.A(G330), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n723), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n721), .A2(KEYINPUT93), .A3(G330), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1016), .A2(new_n732), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1017), .A2(new_n782), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT110), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n732), .A2(new_n729), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(new_n1011), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n732), .A2(KEYINPUT45), .A3(new_n729), .A4(new_n992), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT44), .B1(new_n1028), .B2(new_n1011), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n1011), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n726), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT110), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1017), .A2(new_n1037), .A3(new_n1024), .A4(new_n782), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1031), .B(new_n726), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1026), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1015), .B1(new_n1040), .B2(new_n782), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1013), .B1(new_n1041), .B2(new_n834), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n845), .B(new_n830), .C1(new_n734), .C2(new_n577), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n839), .A2(new_n235), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n836), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n801), .A2(new_n320), .B1(new_n799), .B2(new_n886), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n271), .B(new_n1046), .C1(G50), .C2(new_n794), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n804), .A2(new_n819), .B1(new_n811), .B2(new_n293), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G58), .B2(new_n816), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n874), .A2(new_n884), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n815), .A2(G68), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G107), .A2(new_n815), .B1(new_n805), .B2(G294), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n542), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G311), .A2(new_n874), .B1(new_n875), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n261), .B1(new_n883), .B2(G303), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G283), .A2(new_n794), .B1(new_n871), .B2(G317), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n812), .A2(new_n530), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT46), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT47), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n830), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n845), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1045), .B1(new_n1063), .B2(new_n1064), .C1(new_n1005), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1042), .A2(new_n1066), .ZN(G387));
  NAND2_X1  g0867(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(new_n833), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n706), .A2(new_n1065), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n883), .A2(G317), .B1(new_n794), .B2(G303), .ZN(new_n1071));
  INV_X1    g0871(.A(G311), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n804), .C1(new_n802), .C2(new_n788), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n810), .B2(new_n785), .C1(new_n786), .C2(new_n812), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(KEYINPUT49), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n271), .B1(new_n799), .B2(new_n789), .C1(new_n530), .C2(new_n811), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(KEYINPUT49), .B2(new_n1078), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n816), .A2(G77), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n320), .B2(new_n799), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT112), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n788), .A2(new_n819), .B1(new_n811), .B2(new_n220), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n577), .B2(new_n815), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n261), .B1(new_n793), .B2(new_n242), .C1(new_n240), .C2(new_n801), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n331), .B2(new_n805), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n869), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(G45), .B(new_n738), .C1(G68), .C2(G77), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n440), .A2(G50), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT50), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n839), .C1(new_n457), .C2(new_n232), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n837), .A2(new_n738), .B1(new_n426), .B2(new_n734), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT111), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n836), .B(new_n1091), .C1(new_n846), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1069), .B1(new_n1070), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT114), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n782), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1068), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(KEYINPUT114), .B(new_n782), .C1(new_n1017), .C2(new_n1024), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n736), .B1(new_n1026), .B2(new_n1038), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(KEYINPUT113), .B(new_n736), .C1(new_n1026), .C2(new_n1038), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1101), .B1(new_n1109), .B2(new_n1110), .ZN(G393));
  NAND3_X1  g0911(.A1(new_n1036), .A2(new_n834), .A3(new_n1039), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n846), .B1(new_n210), .B2(new_n542), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n239), .A2(new_n734), .A3(new_n261), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n835), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n785), .A2(new_n293), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n804), .A2(new_n240), .B1(new_n811), .B2(new_n579), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G68), .C2(new_n816), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n320), .A2(new_n788), .B1(new_n801), .B2(new_n819), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n440), .A2(new_n793), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n271), .B(new_n1121), .C1(new_n871), .C2(new_n884), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1072), .A2(new_n801), .B1(new_n788), .B2(new_n806), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT52), .Z(new_n1125));
  OAI221_X1 g0925(.A(new_n271), .B1(new_n799), .B2(new_n802), .C1(new_n786), .C2(new_n793), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n426), .A2(new_n811), .B1(new_n812), .B2(new_n810), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n785), .A2(new_n530), .B1(new_n804), .B2(new_n553), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1123), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1115), .B1(new_n1130), .B2(new_n830), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n992), .B2(new_n1065), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1040), .A2(new_n735), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1026), .A2(new_n1038), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1112), .B(new_n1132), .C1(new_n1133), .C2(new_n1134), .ZN(G390));
  AOI21_X1  g0935(.A(new_n724), .B1(new_n753), .B2(new_n968), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(new_n970), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n859), .A2(new_n918), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n916), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n959), .B1(new_n1139), .B2(new_n960), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n972), .A2(new_n960), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n743), .A2(new_n747), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n857), .A2(new_n450), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n698), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n918), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1141), .B1(new_n1145), .B2(new_n916), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1137), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n972), .A2(new_n957), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n938), .B2(new_n957), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n919), .B2(new_n961), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n781), .A2(G330), .A3(new_n858), .A4(new_n916), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n856), .B1(new_n748), .B2(new_n1143), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(new_n917), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n1151), .C1(new_n1153), .C2(new_n1141), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n833), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G137), .A2(new_n805), .B1(new_n875), .B2(G50), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n788), .C1(new_n819), .C2(new_n785), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n816), .A2(G150), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n261), .B1(new_n799), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n801), .A2(new_n880), .B1(new_n793), .B2(new_n1164), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1159), .A2(new_n1161), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G107), .A2(new_n805), .B1(new_n874), .B2(G283), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n579), .B2(new_n812), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n261), .B1(new_n871), .B2(G294), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n530), .B2(new_n801), .C1(new_n542), .C2(new_n793), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n811), .A2(new_n242), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1116), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n830), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n835), .C1(new_n331), .C2(new_n870), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1149), .B2(new_n843), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT115), .Z(new_n1176));
  NOR2_X1   g0976(.A1(new_n1156), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n781), .A2(G330), .A3(new_n858), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1178), .A2(new_n917), .B1(new_n970), .B2(new_n1136), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1138), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n916), .B1(new_n1136), .B2(new_n858), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1179), .A2(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n452), .A2(new_n1136), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n670), .A2(new_n964), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1155), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1147), .A2(new_n1154), .A3(new_n1185), .A4(new_n1183), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n735), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1177), .A2(new_n1189), .ZN(G378));
  NAND2_X1  g0990(.A1(new_n335), .A2(new_n693), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT55), .Z(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n352), .B2(new_n358), .ZN(new_n1193));
  XOR2_X1   g0993(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1194));
  INV_X1    g0994(.A(new_n1192), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n351), .A2(new_n1195), .A3(new_n357), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1194), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n351), .A2(new_n1195), .A3(new_n357), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n351), .B2(new_n357), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n843), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n835), .B1(new_n870), .B2(G50), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n271), .A2(new_n253), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n240), .C1(G33), .C2(G41), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n801), .A2(new_n426), .B1(new_n799), .B2(new_n810), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n577), .C2(new_n794), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n788), .A2(new_n530), .B1(new_n811), .B2(new_n218), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G97), .B2(new_n805), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n1051), .A3(new_n1083), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n801), .A2(new_n1158), .B1(new_n812), .B2(new_n1164), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT116), .Z(new_n1216));
  AOI22_X1  g1016(.A1(new_n874), .A2(G125), .B1(new_n794), .B2(G137), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G132), .A2(new_n805), .B1(new_n815), .B2(G150), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT117), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n875), .A2(G159), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n871), .C2(G124), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1214), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1204), .B1(new_n1227), .B2(new_n830), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1203), .A2(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT119), .Z(new_n1230));
  NOR3_X1   g1030(.A1(new_n981), .A2(new_n724), .A3(new_n1202), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1202), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n979), .B2(G330), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT120), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n962), .B1(new_n944), .B2(new_n945), .ZN(new_n1235));
  AOI211_X1 g1035(.A(KEYINPUT107), .B(new_n940), .C1(new_n919), .C2(new_n938), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1235), .A2(KEYINPUT121), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1202), .B1(new_n981), .B2(new_n724), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n979), .A2(G330), .A3(new_n1232), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(KEYINPUT121), .B1(new_n963), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1149), .A2(new_n960), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n942), .B2(KEYINPUT107), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT121), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n946), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT120), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1238), .A2(new_n1242), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1230), .B1(new_n1250), .B2(new_n834), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1188), .A2(new_n1185), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1188), .A2(KEYINPUT122), .A3(new_n1185), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1256), .B2(new_n1250), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT57), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n963), .A2(new_n1241), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1244), .A2(new_n946), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1188), .A2(KEYINPUT122), .A3(new_n1185), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT122), .B1(new_n1188), .B2(new_n1185), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n735), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1251), .B1(new_n1257), .B2(new_n1265), .ZN(G375));
  OR2_X1    g1066(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1015), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1186), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n917), .A2(new_n843), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n835), .B1(new_n870), .B2(G68), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n785), .A2(new_n240), .B1(new_n812), .B2(new_n819), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G132), .B2(new_n874), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n271), .B1(new_n871), .B2(G128), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n883), .A2(G137), .B1(new_n794), .B2(G150), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1164), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n805), .A2(new_n1276), .B1(new_n875), .B2(G58), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n271), .B1(new_n811), .B2(new_n293), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT123), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n793), .A2(new_n426), .B1(new_n799), .B2(new_n553), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G283), .B2(new_n883), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n577), .A2(new_n815), .B1(new_n805), .B2(G116), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(G294), .A2(new_n874), .B1(new_n816), .B2(G97), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1278), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1271), .B1(new_n1286), .B2(new_n830), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1183), .A2(new_n834), .B1(new_n1270), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1269), .A2(new_n1288), .ZN(G381));
  OR4_X1    g1089(.A1(G384), .A2(G390), .A3(G378), .A4(G381), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n854), .B(new_n1101), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1291));
  OR4_X1    g1091(.A1(G387), .A2(new_n1290), .A3(G375), .A4(new_n1291), .ZN(G407));
  INV_X1    g1092(.A(G378), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n695), .A2(new_n696), .A3(G213), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G407), .B(G213), .C1(G375), .C2(new_n1296), .ZN(G409));
  OAI211_X1 g1097(.A(G378), .B(new_n1251), .C1(new_n1257), .C2(new_n1265), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1250), .B(new_n1268), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n833), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1229), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n834), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(KEYINPUT124), .A3(new_n1229), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1299), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1293), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1295), .B1(new_n1298), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1186), .A2(KEYINPUT60), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1312), .A2(new_n1267), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n735), .B1(new_n1312), .B2(new_n1267), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1288), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G384), .B(new_n1288), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1309), .A2(new_n1310), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1295), .A2(G2897), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1316), .A2(new_n1317), .A3(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1321), .B1(new_n1309), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1310), .B1(new_n1309), .B2(new_n1319), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1320), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G393), .A2(G396), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1291), .ZN(new_n1331));
  INV_X1    g1131(.A(G390), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G387), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1042), .A2(new_n1066), .A3(G390), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT125), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1331), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1042), .A2(new_n1066), .A3(G390), .ZN(new_n1338));
  AOI21_X1  g1138(.A(G390), .B1(new_n1042), .B2(new_n1066), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1331), .B(new_n1336), .C1(new_n1338), .C2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1298), .A2(new_n1308), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1294), .ZN(new_n1344));
  AND2_X1   g1144(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1343), .A2(new_n1294), .A3(new_n1319), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1346), .A2(new_n1342), .A3(new_n1349), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1343), .A2(KEYINPUT63), .A3(new_n1294), .A4(new_n1319), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT126), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1309), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1319), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  OAI22_X1  g1155(.A1(new_n1329), .A2(new_n1342), .B1(new_n1350), .B2(new_n1355), .ZN(G405));
  INV_X1    g1156(.A(KEYINPUT127), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1357), .B1(new_n1337), .B2(new_n1341), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1336), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1359), .A2(new_n1291), .A3(new_n1330), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1360), .A2(KEYINPUT127), .A3(new_n1340), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(G375), .A2(new_n1293), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n1298), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1364), .A2(new_n1319), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1363), .A2(new_n1298), .A3(new_n1318), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1362), .A2(new_n1367), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1358), .A2(new_n1361), .A3(new_n1365), .A4(new_n1366), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1368), .A2(new_n1369), .ZN(G402));
endmodule


