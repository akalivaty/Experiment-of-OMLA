//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  AOI22_X1  g031(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g048(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n474));
  OAI221_X1 g049(.A(G2104), .B1(G112), .B2(new_n463), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n476), .A2(new_n477), .B1(G136), .B2(new_n462), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n461), .B2(new_n463), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n478), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n459), .B2(new_n460), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n497), .C1(new_n460), .C2(new_n459), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n502), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(G88), .B1(G50), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(G50), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n517), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n508), .B1(new_n516), .B2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(new_n511), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n505), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n503), .A2(new_n504), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n532), .B1(new_n510), .B2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n525), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n541), .B1(new_n537), .B2(new_n538), .C1(new_n536), .C2(new_n525), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n505), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n534), .B1(new_n546), .B2(KEYINPUT73), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(KEYINPUT73), .B2(new_n546), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT74), .B(G43), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n512), .A2(G81), .B1(new_n513), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n513), .A2(G53), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n532), .A2(G65), .ZN(new_n562));
  INV_X1    g137(.A(G78), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT76), .B1(new_n563), .B2(new_n502), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n563), .A2(new_n502), .A3(KEYINPUT76), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n512), .A2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  OAI21_X1  g148(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n512), .A2(G87), .B1(G49), .B2(new_n513), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n512), .A2(G86), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n503), .B2(new_n504), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g158(.A(G48), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n578), .A2(new_n583), .A3(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n512), .A2(G85), .B1(G47), .B2(new_n513), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n534), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT78), .ZN(G290));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n590));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(G171), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n513), .A2(G54), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n532), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT80), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n534), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n595), .B1(new_n594), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n512), .A2(G92), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT10), .Z(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI211_X1 g180(.A(new_n590), .B(new_n592), .C1(new_n591), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n590), .B2(new_n592), .ZN(G284));
  AOI21_X1  g182(.A(new_n606), .B1(new_n590), .B2(new_n592), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n570), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n570), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(new_n605), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n482), .A2(new_n464), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n623), .A2(KEYINPUT82), .A3(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT82), .B1(new_n623), .B2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n462), .A2(G135), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n484), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n622), .A2(G2100), .B1(G2096), .B2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n631), .B(new_n632), .C1(G2100), .C2(new_n622), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT84), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n658), .B2(new_n654), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT86), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n654), .A3(new_n652), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n653), .A3(new_n652), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT88), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT91), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(new_n677), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n681), .C1(new_n675), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT90), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G1986), .ZN(new_n686));
  INV_X1    g261(.A(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n672), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n690), .A3(new_n672), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n693), .ZN(new_n696));
  INV_X1    g271(.A(new_n694), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT29), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G2090), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G20), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT23), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n570), .B2(new_n707), .ZN(new_n710));
  INV_X1    g285(.A(G1956), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n706), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n716));
  NOR2_X1   g291(.A1(G4), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n612), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT99), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT100), .B(G1348), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n719), .A2(new_n721), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G19), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n552), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT101), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1341), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n722), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n701), .A2(G33), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(new_n463), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT102), .B(KEYINPUT25), .Z(new_n732));
  NAND3_X1  g307(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  AOI211_X1 g309(.A(new_n731), .B(new_n734), .C1(G139), .C2(new_n462), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n729), .B1(new_n735), .B2(new_n701), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G2072), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(G164), .A2(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G27), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NOR4_X1   g318(.A1(new_n737), .A2(new_n738), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n484), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G129), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n464), .A2(G105), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n747), .B(new_n749), .C1(G141), .C2(new_n462), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(new_n701), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n701), .B2(G32), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n707), .A2(G21), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G168), .B2(new_n707), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT106), .B(G1966), .Z(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  OR2_X1    g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  NAND2_X1  g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n762), .A2(new_n701), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT103), .B(KEYINPUT24), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G34), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(new_n701), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n470), .B2(new_n701), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n765), .B1(new_n701), .B2(new_n630), .C1(new_n770), .C2(G2084), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n756), .A2(new_n761), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(G2084), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT104), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n744), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n701), .A2(G26), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT28), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n745), .A2(G128), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n779));
  INV_X1    g354(.A(G116), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G2105), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n462), .B2(G140), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n777), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n707), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n707), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1961), .Z(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n788), .C1(new_n704), .C2(G2090), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n754), .A2(new_n755), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT105), .Z(new_n791));
  NOR3_X1   g366(.A1(new_n775), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n728), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n715), .A2(new_n716), .A3(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT32), .B(G1981), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n707), .A2(G22), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT97), .Z(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n707), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(G16), .A2(G23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G288), .B2(new_n707), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n805), .B(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n796), .B2(new_n797), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n798), .A2(new_n803), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n462), .A2(G131), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n463), .A2(G107), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(G119), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n814), .B1(new_n815), .B2(new_n816), .C1(new_n484), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT92), .ZN(new_n819));
  MUX2_X1   g394(.A(G25), .B(new_n819), .S(G29), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G24), .B(G290), .S(G16), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(G1986), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n811), .A2(new_n812), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n813), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT98), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n826), .A3(new_n830), .A4(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(KEYINPUT36), .A3(new_n831), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n794), .A2(new_n834), .A3(new_n835), .ZN(G311));
  NAND3_X1  g411(.A1(new_n794), .A2(new_n834), .A3(new_n835), .ZN(G150));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n525), .A2(new_n838), .B1(new_n537), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n534), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n613), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n548), .A2(new_n843), .A3(new_n550), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n843), .B1(new_n548), .B2(new_n550), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n848), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT109), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n844), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n846), .B1(new_n856), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(G160), .B(new_n630), .ZN(new_n859));
  XNOR2_X1  g434(.A(G162), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n462), .A2(G142), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n463), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G130), .B2(new_n745), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n620), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n818), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n751), .B(new_n783), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n496), .A2(new_n498), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n487), .A2(new_n491), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n868), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(new_n735), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n735), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT110), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n867), .A3(new_n874), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g453(.A(KEYINPUT110), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n860), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n860), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n875), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g461(.A(new_n591), .B1(new_n840), .B2(new_n842), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n615), .B(new_n852), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n602), .A2(new_n570), .A3(new_n604), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n570), .B1(new_n602), .B2(new_n604), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n605), .A2(G299), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n602), .A2(new_n570), .A3(new_n604), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n891), .A2(new_n892), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n888), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT42), .ZN(new_n903));
  XNOR2_X1  g478(.A(G290), .B(G166), .ZN(new_n904));
  XOR2_X1   g479(.A(G288), .B(G305), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n903), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n887), .B1(new_n908), .B2(new_n591), .ZN(G295));
  OAI21_X1  g484(.A(new_n887), .B1(new_n908), .B2(new_n591), .ZN(G331));
  INV_X1    g485(.A(new_n851), .ZN(new_n911));
  AOI21_X1  g486(.A(G301), .B1(new_n911), .B2(new_n849), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n850), .A2(G171), .A3(new_n851), .ZN(new_n913));
  OAI21_X1  g488(.A(G286), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(G171), .B1(new_n850), .B2(new_n851), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(G301), .A3(new_n849), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(G168), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n901), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n898), .A2(new_n914), .A3(new_n920), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n915), .A2(new_n916), .A3(G168), .ZN(new_n923));
  AOI21_X1  g498(.A(G168), .B1(new_n915), .B2(new_n916), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n925), .B2(new_n898), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n907), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT112), .B1(new_n918), .B2(new_n899), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n906), .A3(new_n919), .A4(new_n921), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(new_n928), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n901), .A2(new_n890), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(KEYINPUT41), .B2(new_n901), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n919), .B1(new_n918), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G37), .B1(new_n935), .B2(new_n907), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n930), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n932), .C1(new_n937), .C2(new_n928), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n927), .A2(new_n931), .A3(new_n930), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n928), .A3(new_n930), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT113), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n945), .B(KEYINPUT44), .C1(new_n940), .C2(new_n941), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n944), .B2(new_n946), .ZN(G397));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n871), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT45), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n465), .A2(new_n469), .A3(G40), .ZN(new_n952));
  NOR2_X1   g527(.A1(G164), .A2(G1384), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT114), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n783), .A2(G2067), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n783), .A2(G2067), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(G1996), .B2(new_n751), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n955), .A2(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n752), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n962), .A2(KEYINPUT115), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(KEYINPUT115), .ZN(new_n964));
  OAI22_X1  g539(.A1(new_n960), .A2(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n965), .A2(new_n819), .A3(new_n821), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n955), .B1(new_n966), .B2(new_n956), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n961), .B(KEYINPUT46), .Z(new_n968));
  INV_X1    g543(.A(new_n955), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n959), .B2(new_n751), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n818), .B(new_n821), .Z(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(new_n955), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(G290), .A2(new_n955), .A3(G1986), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT48), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n967), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT126), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT116), .B1(G164), .B2(G1384), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  INV_X1    g560(.A(new_n498), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n497), .B1(new_n482), .B2(new_n494), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n985), .B(new_n948), .C1(new_n988), .C2(new_n492), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n983), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n983), .A2(new_n989), .A3(new_n991), .A4(new_n984), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n465), .A2(new_n469), .A3(G40), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G2084), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n985), .B1(new_n871), .B2(new_n948), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT116), .B(G1384), .C1(new_n869), .C2(new_n870), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n953), .B2(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n995), .A2(new_n997), .B1(new_n1003), .B2(new_n759), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n982), .B1(new_n1004), .B2(G168), .ZN(new_n1005));
  INV_X1    g580(.A(new_n997), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n993), .B2(new_n994), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n760), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1008));
  OAI21_X1  g583(.A(G286), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n981), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT51), .B(new_n982), .C1(new_n1004), .C2(G168), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT62), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1013));
  AND3_X1   g588(.A1(G303), .A2(G8), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(G303), .B2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g591(.A(G2090), .B(new_n996), .C1(new_n993), .C2(new_n994), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n949), .A2(new_n998), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1002), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n802), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(G8), .B(new_n1016), .C1(new_n1017), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G86), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n584), .B1(new_n537), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n583), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n578), .A2(new_n687), .A3(new_n583), .A4(new_n584), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G305), .A2(KEYINPUT119), .A3(G1981), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n983), .A2(new_n952), .A3(new_n989), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(new_n1034), .A3(new_n1030), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(G8), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G288), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT52), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(G8), .A4(new_n1033), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1036), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1022), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n984), .B1(new_n983), .B2(new_n989), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n996), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT50), .B1(new_n999), .B2(new_n1000), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT120), .A3(new_n952), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n953), .A2(new_n984), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1020), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1016), .B1(new_n1054), .B2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1019), .B2(G2078), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1001), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n1002), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n996), .B1(new_n993), .B2(new_n994), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(G1961), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G171), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1045), .A2(new_n1055), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n995), .A2(new_n997), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1008), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(G168), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(G8), .A3(new_n1009), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT51), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1005), .A2(new_n981), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1012), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n982), .B1(new_n1053), .B2(new_n1020), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1022), .B(new_n1044), .C1(new_n1073), .C2(new_n1016), .ZN(new_n1074));
  NOR2_X1   g649(.A1(G286), .A2(new_n982), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(new_n1022), .A3(new_n1081), .A4(new_n1044), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1036), .A2(new_n1038), .A3(new_n575), .A4(new_n576), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1037), .B1(new_n1084), .B2(new_n1027), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1022), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(new_n1044), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1071), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  NAND2_X1  g664(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1090), .B(new_n1093), .C1(new_n561), .C2(new_n569), .ZN(new_n1094));
  INV_X1    g669(.A(new_n569), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n559), .B(KEYINPUT9), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n711), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(G2072), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1002), .A2(new_n1018), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1099), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1104), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1106), .B(new_n1098), .C1(new_n1100), .C2(new_n711), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1089), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1098), .B(KEYINPUT123), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n983), .A2(new_n989), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n996), .B1(new_n1110), .B2(KEYINPUT50), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1111), .A2(KEYINPUT120), .B1(new_n984), .B2(new_n953), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1956), .B1(new_n1112), .B2(new_n1048), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1113), .B2(new_n1106), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1106), .B1(new_n1100), .B2(new_n711), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1099), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n953), .A2(KEYINPUT45), .ZN(new_n1118));
  INV_X1    g693(.A(G1996), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1018), .A3(new_n1119), .A4(new_n952), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1033), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n551), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1033), .A2(G2067), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT60), .B(new_n1126), .C1(new_n1059), .C2(new_n721), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(new_n605), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1059), .B2(new_n721), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n612), .A3(new_n1127), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1108), .A2(new_n1117), .A3(new_n1129), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n612), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1098), .B(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1115), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1139), .B2(new_n1116), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1135), .A3(new_n1116), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1134), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1045), .A2(new_n1055), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1060), .A2(G171), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n951), .A2(new_n954), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n1002), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1149), .B(new_n1057), .C1(new_n1059), .C2(G1961), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(G171), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1146), .B1(new_n1150), .B2(G171), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(G171), .B2(new_n1060), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1144), .A2(new_n1145), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1088), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(G290), .B(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n975), .B1(new_n969), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n980), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1139), .A2(new_n1135), .A3(new_n1116), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n1140), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1155), .B1(new_n1163), .B2(new_n1134), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1071), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n980), .B(new_n1160), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n979), .B1(new_n1161), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g743(.A1(new_n650), .A2(new_n457), .ZN(new_n1170));
  NOR2_X1   g744(.A1(G227), .A2(new_n1170), .ZN(new_n1171));
  AND4_X1   g745(.A1(new_n699), .A2(new_n942), .A3(new_n885), .A4(new_n1171), .ZN(G308));
  NAND4_X1  g746(.A1(new_n699), .A2(new_n885), .A3(new_n942), .A4(new_n1171), .ZN(G225));
endmodule


