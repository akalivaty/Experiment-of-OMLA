

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829;

  NOR2_X1 U375 ( .A1(G902), .A2(n787), .ZN(n614) );
  XNOR2_X1 U376 ( .A(n377), .B(n511), .ZN(n787) );
  NOR2_X1 U377 ( .A1(n674), .A2(n653), .ZN(n654) );
  INV_X1 U378 ( .A(G953), .ZN(n817) );
  XOR2_X1 U379 ( .A(n602), .B(n601), .Z(n353) );
  AND2_X1 U380 ( .A1(n658), .A2(n532), .ZN(n354) );
  XOR2_X1 U381 ( .A(n709), .B(KEYINPUT90), .Z(n355) );
  AND2_X1 U382 ( .A1(n766), .A2(n779), .ZN(n356) );
  AND2_X1 U383 ( .A1(n412), .A2(n404), .ZN(n357) );
  AND2_X1 U384 ( .A1(n416), .A2(n415), .ZN(n358) );
  AND2_X1 U385 ( .A1(n407), .A2(n406), .ZN(n359) );
  AND2_X1 U386 ( .A1(n515), .A2(n423), .ZN(n360) );
  XNOR2_X1 U387 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n361) );
  XOR2_X1 U388 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n362) );
  OR2_X1 U389 ( .A1(n516), .A2(KEYINPUT121), .ZN(n519) );
  AND2_X1 U390 ( .A1(n558), .A2(G475), .ZN(n542) );
  XNOR2_X2 U391 ( .A(n644), .B(KEYINPUT35), .ZN(n825) );
  NAND2_X2 U392 ( .A1(n359), .A2(n378), .ZN(n644) );
  NAND2_X2 U393 ( .A1(n566), .A2(n565), .ZN(n568) );
  INV_X1 U394 ( .A(n674), .ZN(n363) );
  XNOR2_X2 U395 ( .A(n553), .B(n541), .ZN(n453) );
  NOR2_X2 U396 ( .A1(n708), .A2(n709), .ZN(n649) );
  XNOR2_X2 U397 ( .A(n671), .B(KEYINPUT1), .ZN(n709) );
  INV_X1 U398 ( .A(n777), .ZN(n450) );
  NAND2_X1 U399 ( .A1(n645), .A2(n647), .ZN(n728) );
  XNOR2_X1 U400 ( .A(n485), .B(KEYINPUT48), .ZN(n392) );
  AND2_X1 U401 ( .A1(n400), .A2(n675), .ZN(n498) );
  NOR2_X1 U402 ( .A1(n674), .A2(n401), .ZN(n400) );
  NOR2_X1 U403 ( .A1(n731), .A2(n728), .ZN(n394) );
  NAND2_X1 U404 ( .A1(n499), .A2(n364), .ZN(n401) );
  AND2_X1 U405 ( .A1(n439), .A2(n677), .ZN(n499) );
  NAND2_X1 U406 ( .A1(n355), .A2(n636), .ZN(n370) );
  XNOR2_X1 U407 ( .A(n697), .B(KEYINPUT38), .ZN(n725) );
  INV_X1 U408 ( .A(n638), .ZN(n680) );
  XNOR2_X1 U409 ( .A(n660), .B(n528), .ZN(n675) );
  AND2_X1 U410 ( .A1(n402), .A2(n456), .ZN(n405) );
  XNOR2_X1 U411 ( .A(n377), .B(n634), .ZN(n761) );
  XNOR2_X1 U412 ( .A(n381), .B(n380), .ZN(n647) );
  OR2_X1 U413 ( .A1(n793), .A2(G902), .ZN(n381) );
  XNOR2_X1 U414 ( .A(n383), .B(n382), .ZN(n645) );
  OR2_X1 U415 ( .A1(n704), .A2(G902), .ZN(n383) );
  INV_X1 U416 ( .A(KEYINPUT89), .ZN(n533) );
  INV_X1 U417 ( .A(G478), .ZN(n380) );
  XNOR2_X1 U418 ( .A(n365), .B(n362), .ZN(G60) );
  NAND2_X1 U419 ( .A1(n465), .A2(n464), .ZN(n365) );
  AND2_X1 U420 ( .A1(n515), .A2(n420), .ZN(n397) );
  NAND2_X1 U421 ( .A1(n480), .A2(n542), .ZN(n707) );
  NOR2_X1 U422 ( .A1(n816), .A2(n432), .ZN(n468) );
  NAND2_X1 U423 ( .A1(n388), .A2(n434), .ZN(n387) );
  AND2_X1 U424 ( .A1(n411), .A2(n404), .ZN(n403) );
  NAND2_X1 U425 ( .A1(n414), .A2(n413), .ZN(n404) );
  NOR2_X1 U426 ( .A1(n495), .A2(n492), .ZN(n491) );
  NAND2_X1 U427 ( .A1(n824), .A2(n533), .ZN(n415) );
  AND2_X1 U428 ( .A1(n536), .A2(n418), .ZN(n535) );
  NAND2_X1 U429 ( .A1(n540), .A2(n538), .ZN(n534) );
  NAND2_X1 U430 ( .A1(n410), .A2(n379), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n551), .B(n550), .ZN(n824) );
  XNOR2_X1 U432 ( .A(n498), .B(KEYINPUT111), .ZN(n826) );
  NOR2_X1 U433 ( .A1(n650), .A2(n718), .ZN(n651) );
  XNOR2_X1 U434 ( .A(n394), .B(n510), .ZN(n722) );
  OR2_X1 U435 ( .A1(n774), .A2(n691), .ZN(n692) );
  INV_X1 U436 ( .A(n655), .ZN(n369) );
  NOR2_X1 U437 ( .A1(n730), .A2(n689), .ZN(n366) );
  AND2_X1 U438 ( .A1(n649), .A2(n638), .ZN(n639) );
  NAND2_X1 U439 ( .A1(n724), .A2(n715), .ZN(n660) );
  XNOR2_X1 U440 ( .A(n715), .B(n361), .ZN(n638) );
  XNOR2_X1 U441 ( .A(n648), .B(KEYINPUT104), .ZN(n688) );
  NAND2_X2 U442 ( .A1(n457), .A2(n405), .ZN(n715) );
  XNOR2_X1 U443 ( .A(n761), .B(KEYINPUT62), .ZN(n762) );
  NOR2_X1 U444 ( .A1(n647), .A2(n646), .ZN(n770) );
  OR2_X1 U445 ( .A1(n761), .A2(n454), .ZN(n402) );
  INV_X1 U446 ( .A(n676), .ZN(n364) );
  XNOR2_X1 U447 ( .A(n608), .B(n353), .ZN(n793) );
  XNOR2_X1 U448 ( .A(n598), .B(n597), .ZN(n704) );
  XNOR2_X1 U449 ( .A(n577), .B(KEYINPUT94), .ZN(n578) );
  XNOR2_X1 U450 ( .A(n615), .B(n502), .ZN(n813) );
  XNOR2_X1 U451 ( .A(n376), .B(n531), .ZN(n612) );
  NAND2_X1 U452 ( .A1(G214), .A2(n579), .ZN(n724) );
  INV_X1 U453 ( .A(n562), .ZN(n382) );
  XNOR2_X1 U454 ( .A(n603), .B(n385), .ZN(n384) );
  INV_X1 U455 ( .A(n659), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n575), .B(KEYINPUT92), .ZN(n699) );
  XNOR2_X1 U457 ( .A(n569), .B(G107), .ZN(n805) );
  XNOR2_X1 U458 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n367) );
  XNOR2_X1 U459 ( .A(G146), .B(G125), .ZN(n570) );
  XNOR2_X1 U460 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n385) );
  INV_X1 U461 ( .A(G113), .ZN(n564) );
  XNOR2_X1 U462 ( .A(G143), .B(G113), .ZN(n588) );
  XNOR2_X1 U463 ( .A(G110), .B(G104), .ZN(n569) );
  INV_X1 U464 ( .A(KEYINPUT69), .ZN(n549) );
  NAND2_X1 U465 ( .A1(n522), .A2(n431), .ZN(n494) );
  NAND2_X1 U466 ( .A1(n523), .A2(n363), .ZN(n522) );
  NOR2_X1 U467 ( .A1(n690), .A2(n366), .ZN(n691) );
  XNOR2_X1 U468 ( .A(n615), .B(n367), .ZN(n598) );
  NOR2_X2 U469 ( .A1(n764), .A2(n368), .ZN(n658) );
  NOR2_X1 U470 ( .A1(n356), .A2(n369), .ZN(n368) );
  NAND2_X1 U471 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X2 U472 ( .A1(n358), .A2(n658), .ZN(n375) );
  NOR2_X1 U473 ( .A1(n637), .A2(n370), .ZN(n551) );
  NAND2_X1 U474 ( .A1(n371), .A2(n354), .ZN(n374) );
  NAND2_X1 U475 ( .A1(n403), .A2(n358), .ZN(n371) );
  XNOR2_X2 U476 ( .A(n372), .B(n395), .ZN(n745) );
  NAND2_X1 U477 ( .A1(n375), .A2(n357), .ZN(n373) );
  XNOR2_X1 U478 ( .A(n703), .B(KEYINPUT75), .ZN(n750) );
  NOR2_X1 U479 ( .A1(n745), .A2(n746), .ZN(n561) );
  XNOR2_X1 U480 ( .A(n376), .B(n384), .ZN(n607) );
  XNOR2_X2 U481 ( .A(n386), .B(G143), .ZN(n376) );
  XNOR2_X2 U482 ( .A(n814), .B(G146), .ZN(n377) );
  INV_X1 U483 ( .A(n735), .ZN(n379) );
  XNOR2_X2 U484 ( .A(G128), .B(KEYINPUT79), .ZN(n386) );
  NAND2_X2 U485 ( .A1(n389), .A2(n387), .ZN(n816) );
  INV_X1 U486 ( .A(n392), .ZN(n388) );
  AND2_X2 U487 ( .A1(n390), .A2(n430), .ZN(n389) );
  NAND2_X1 U488 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U489 ( .A(KEYINPUT85), .ZN(n391) );
  XNOR2_X2 U490 ( .A(n393), .B(KEYINPUT42), .ZN(n827) );
  NAND2_X1 U491 ( .A1(n428), .A2(n722), .ZN(n393) );
  XNOR2_X1 U492 ( .A(n651), .B(KEYINPUT31), .ZN(n779) );
  XNOR2_X1 U493 ( .A(n654), .B(KEYINPUT97), .ZN(n766) );
  NAND2_X1 U494 ( .A1(n396), .A2(n521), .ZN(n399) );
  NAND2_X1 U495 ( .A1(n397), .A2(n519), .ZN(n396) );
  NAND2_X1 U496 ( .A1(n399), .A2(n398), .ZN(G75) );
  NAND2_X1 U497 ( .A1(n360), .A2(n519), .ZN(n398) );
  NAND2_X1 U498 ( .A1(n735), .A2(n642), .ZN(n406) );
  INV_X1 U499 ( .A(n408), .ZN(n407) );
  NAND2_X1 U500 ( .A1(n409), .A2(n643), .ZN(n408) );
  NAND2_X1 U501 ( .A1(n650), .A2(n642), .ZN(n409) );
  NOR2_X1 U502 ( .A1(n650), .A2(n642), .ZN(n410) );
  XNOR2_X2 U503 ( .A(n639), .B(KEYINPUT33), .ZN(n735) );
  INV_X1 U504 ( .A(n825), .ZN(n411) );
  NOR2_X1 U505 ( .A1(n825), .A2(n532), .ZN(n412) );
  INV_X1 U506 ( .A(n829), .ZN(n413) );
  NOR2_X1 U507 ( .A1(n824), .A2(n533), .ZN(n414) );
  NAND2_X1 U508 ( .A1(n829), .A2(n533), .ZN(n416) );
  NAND2_X1 U509 ( .A1(n678), .A2(n584), .ZN(n586) );
  XNOR2_X2 U510 ( .A(n417), .B(KEYINPUT19), .ZN(n678) );
  NAND2_X2 U511 ( .A1(n661), .A2(n724), .ZN(n417) );
  XNOR2_X2 U512 ( .A(n451), .B(n578), .ZN(n661) );
  AND2_X1 U513 ( .A1(n478), .A2(n468), .ZN(n467) );
  INV_X1 U514 ( .A(n750), .ZN(n558) );
  AND2_X1 U515 ( .A1(n480), .A2(n558), .ZN(n794) );
  INV_X1 U516 ( .A(KEYINPUT44), .ZN(n532) );
  NOR2_X1 U517 ( .A1(G902), .A2(G237), .ZN(n576) );
  XOR2_X1 U518 ( .A(G134), .B(G131), .Z(n560) );
  XNOR2_X1 U519 ( .A(n570), .B(KEYINPUT10), .ZN(n615) );
  XOR2_X1 U520 ( .A(G137), .B(G140), .Z(n616) );
  XNOR2_X1 U521 ( .A(G902), .B(KEYINPUT15), .ZN(n575) );
  AND2_X1 U522 ( .A1(n682), .A2(n545), .ZN(n544) );
  NOR2_X1 U523 ( .A1(n681), .A2(n546), .ZN(n545) );
  INV_X1 U524 ( .A(n724), .ZN(n546) );
  INV_X1 U525 ( .A(KEYINPUT36), .ZN(n449) );
  AND2_X1 U526 ( .A1(n544), .A2(n450), .ZN(n438) );
  XNOR2_X1 U527 ( .A(n624), .B(KEYINPUT25), .ZN(n625) );
  NOR2_X1 U528 ( .A1(n796), .A2(G902), .ZN(n626) );
  XNOR2_X1 U529 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n484) );
  XNOR2_X1 U530 ( .A(n782), .B(n486), .ZN(n683) );
  INV_X1 U531 ( .A(KEYINPUT87), .ZN(n486) );
  XNOR2_X1 U532 ( .A(G131), .B(G140), .ZN(n590) );
  INV_X1 U533 ( .A(KEYINPUT83), .ZN(n479) );
  NOR2_X1 U534 ( .A1(n436), .A2(n435), .ZN(n434) );
  INV_X1 U535 ( .A(KEYINPUT85), .ZN(n435) );
  XOR2_X1 U536 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n659) );
  XNOR2_X1 U537 ( .A(n738), .B(n483), .ZN(n739) );
  XNOR2_X1 U538 ( .A(KEYINPUT120), .B(KEYINPUT52), .ZN(n483) );
  AND2_X1 U539 ( .A1(n675), .A2(n527), .ZN(n523) );
  INV_X1 U540 ( .A(n529), .ZN(n527) );
  INV_X1 U541 ( .A(KEYINPUT107), .ZN(n539) );
  NOR2_X1 U542 ( .A1(n728), .A2(n681), .ZN(n609) );
  XNOR2_X1 U543 ( .A(n629), .B(n547), .ZN(n633) );
  XOR2_X1 U544 ( .A(KEYINPUT9), .B(G107), .Z(n602) );
  XNOR2_X1 U545 ( .A(n613), .B(n482), .ZN(n511) );
  XNOR2_X1 U546 ( .A(n616), .B(n427), .ZN(n482) );
  INV_X1 U547 ( .A(KEYINPUT84), .ZN(n466) );
  NAND2_X1 U548 ( .A1(n447), .A2(KEYINPUT40), .ZN(n493) );
  AND2_X1 U549 ( .A1(n524), .A2(n490), .ZN(n489) );
  AND2_X1 U550 ( .A1(n450), .A2(n669), .ZN(n490) );
  NOR2_X1 U551 ( .A1(n524), .A2(n669), .ZN(n495) );
  NOR2_X1 U552 ( .A1(n447), .A2(n449), .ZN(n441) );
  AND2_X1 U553 ( .A1(n445), .A2(n444), .ZN(n443) );
  NAND2_X1 U554 ( .A1(n680), .A2(n449), .ZN(n444) );
  NOR2_X1 U555 ( .A1(n694), .A2(n539), .ZN(n538) );
  XNOR2_X1 U556 ( .A(n813), .B(n513), .ZN(n622) );
  XNOR2_X1 U557 ( .A(n710), .B(n484), .ZN(n717) );
  XNOR2_X1 U558 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U559 ( .A(KEYINPUT76), .B(KEYINPUT93), .ZN(n572) );
  XOR2_X1 U560 ( .A(KEYINPUT77), .B(KEYINPUT17), .Z(n573) );
  XNOR2_X1 U561 ( .A(n549), .B(G101), .ZN(n627) );
  NAND2_X1 U562 ( .A1(n497), .A2(n455), .ZN(n454) );
  INV_X1 U563 ( .A(G902), .ZN(n455) );
  NAND2_X1 U564 ( .A1(n761), .A2(n635), .ZN(n457) );
  XNOR2_X1 U565 ( .A(n473), .B(KEYINPUT21), .ZN(n681) );
  NAND2_X1 U566 ( .A1(n623), .A2(G221), .ZN(n473) );
  XNOR2_X1 U567 ( .A(n627), .B(n548), .ZN(n547) );
  XNOR2_X1 U568 ( .A(KEYINPUT5), .B(KEYINPUT96), .ZN(n548) );
  NAND2_X1 U569 ( .A1(n477), .A2(n476), .ZN(n475) );
  NOR2_X1 U570 ( .A1(n699), .A2(n479), .ZN(n476) );
  INV_X1 U571 ( .A(KEYINPUT4), .ZN(n531) );
  XNOR2_X1 U572 ( .A(n587), .B(KEYINPUT18), .ZN(n555) );
  XNOR2_X1 U573 ( .A(n556), .B(n805), .ZN(n613) );
  XNOR2_X1 U574 ( .A(n627), .B(KEYINPUT70), .ZN(n556) );
  NAND2_X1 U575 ( .A1(n725), .A2(n364), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n474), .B(KEYINPUT20), .ZN(n623) );
  NAND2_X1 U577 ( .A1(n699), .A2(G234), .ZN(n474) );
  INV_X1 U578 ( .A(KEYINPUT30), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G234), .A2(G237), .ZN(n581) );
  XNOR2_X1 U580 ( .A(KEYINPUT16), .B(G122), .ZN(n554) );
  INV_X1 U581 ( .A(n616), .ZN(n502) );
  XNOR2_X1 U582 ( .A(n617), .B(n514), .ZN(n513) );
  INV_X1 U583 ( .A(KEYINPUT24), .ZN(n514) );
  XNOR2_X1 U584 ( .A(G128), .B(G110), .ZN(n617) );
  XNOR2_X1 U585 ( .A(n453), .B(n452), .ZN(n755) );
  XNOR2_X1 U586 ( .A(n613), .B(n612), .ZN(n452) );
  XNOR2_X1 U587 ( .A(n555), .B(n571), .ZN(n541) );
  INV_X1 U588 ( .A(KEYINPUT41), .ZN(n510) );
  XNOR2_X1 U589 ( .A(n641), .B(KEYINPUT34), .ZN(n642) );
  INV_X1 U590 ( .A(n671), .ZN(n469) );
  XNOR2_X1 U591 ( .A(n471), .B(n670), .ZN(n470) );
  XNOR2_X1 U592 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U593 ( .A(G116), .B(G122), .ZN(n601) );
  AND2_X1 U594 ( .A1(n558), .A2(G210), .ZN(n503) );
  INV_X1 U595 ( .A(n752), .ZN(n517) );
  NAND2_X1 U596 ( .A1(n446), .A2(n438), .ZN(n693) );
  NAND2_X1 U597 ( .A1(n421), .A2(n489), .ZN(n488) );
  AND2_X1 U598 ( .A1(n504), .A2(n355), .ZN(n782) );
  NAND2_X1 U599 ( .A1(n442), .A2(n441), .ZN(n440) );
  XNOR2_X1 U600 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n550) );
  INV_X1 U601 ( .A(n774), .ZN(n771) );
  INV_X1 U602 ( .A(KEYINPUT108), .ZN(n552) );
  NAND2_X1 U603 ( .A1(n652), .A2(n496), .ZN(n653) );
  INV_X1 U604 ( .A(KEYINPUT63), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n795), .B(n796), .ZN(n512) );
  XNOR2_X1 U606 ( .A(n790), .B(n791), .ZN(n507) );
  AND2_X1 U607 ( .A1(n537), .A2(n429), .ZN(n418) );
  XOR2_X1 U608 ( .A(KEYINPUT88), .B(KEYINPUT39), .Z(n419) );
  AND2_X1 U609 ( .A1(n518), .A2(n817), .ZN(n420) );
  NAND2_X1 U610 ( .A1(n647), .A2(n646), .ZN(n777) );
  NAND2_X1 U611 ( .A1(n522), .A2(n419), .ZN(n421) );
  AND2_X1 U612 ( .A1(n540), .A2(n709), .ZN(n422) );
  AND2_X1 U613 ( .A1(n420), .A2(n753), .ZN(n423) );
  AND2_X1 U614 ( .A1(n558), .A2(G472), .ZN(n424) );
  AND2_X1 U615 ( .A1(n517), .A2(KEYINPUT121), .ZN(n425) );
  OR2_X1 U616 ( .A1(n786), .A2(KEYINPUT85), .ZN(n426) );
  INV_X1 U617 ( .A(n697), .ZN(n439) );
  AND2_X1 U618 ( .A1(G227), .A2(n817), .ZN(n427) );
  AND2_X1 U619 ( .A1(n470), .A2(n469), .ZN(n428) );
  AND2_X1 U620 ( .A1(n496), .A2(n657), .ZN(n429) );
  AND2_X1 U621 ( .A1(n426), .A2(n785), .ZN(n430) );
  AND2_X1 U622 ( .A1(n419), .A2(KEYINPUT40), .ZN(n431) );
  AND2_X1 U623 ( .A1(n699), .A2(n479), .ZN(n432) );
  XOR2_X1 U624 ( .A(n706), .B(n705), .Z(n433) );
  NOR2_X1 U625 ( .A1(G952), .A2(n817), .ZN(n797) );
  INV_X1 U626 ( .A(n797), .ZN(n464) );
  INV_X1 U627 ( .A(n786), .ZN(n436) );
  NAND2_X1 U628 ( .A1(n437), .A2(n449), .ZN(n445) );
  NAND2_X1 U629 ( .A1(n438), .A2(n439), .ZN(n437) );
  INV_X1 U630 ( .A(n450), .ZN(n447) );
  NAND2_X1 U631 ( .A1(n439), .A2(n544), .ZN(n448) );
  INV_X1 U632 ( .A(n680), .ZN(n446) );
  NAND2_X1 U633 ( .A1(n443), .A2(n440), .ZN(n504) );
  NOR2_X1 U634 ( .A1(n680), .A2(n448), .ZN(n442) );
  NAND2_X1 U635 ( .A1(n755), .A2(n699), .ZN(n451) );
  NAND2_X1 U636 ( .A1(n635), .A2(G902), .ZN(n456) );
  XNOR2_X1 U637 ( .A(n792), .B(n793), .ZN(n505) );
  AND2_X1 U638 ( .A1(n682), .A2(n715), .ZN(n472) );
  BUF_X1 U639 ( .A(n804), .Z(n458) );
  NOR2_X1 U640 ( .A1(n708), .A2(n671), .ZN(n530) );
  BUF_X1 U641 ( .A(n755), .Z(n459) );
  NAND2_X1 U642 ( .A1(n804), .A2(n574), .ZN(n462) );
  NAND2_X1 U643 ( .A1(n460), .A2(n461), .ZN(n463) );
  NAND2_X1 U644 ( .A1(n462), .A2(n463), .ZN(n553) );
  INV_X1 U645 ( .A(n804), .ZN(n460) );
  INV_X1 U646 ( .A(n574), .ZN(n461) );
  INV_X1 U647 ( .A(n661), .ZN(n697) );
  INV_X1 U648 ( .A(n753), .ZN(n521) );
  XNOR2_X1 U649 ( .A(n707), .B(n433), .ZN(n465) );
  NAND2_X1 U650 ( .A1(n745), .A2(n479), .ZN(n478) );
  NAND2_X1 U651 ( .A1(n701), .A2(n700), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n751), .B(n466), .ZN(n516) );
  INV_X1 U653 ( .A(n816), .ZN(n702) );
  NAND2_X1 U654 ( .A1(n467), .A2(n475), .ZN(n701) );
  NAND2_X1 U655 ( .A1(n712), .A2(n472), .ZN(n471) );
  INV_X1 U656 ( .A(n745), .ZN(n477) );
  NAND2_X1 U657 ( .A1(n480), .A2(n424), .ZN(n557) );
  NAND2_X1 U658 ( .A1(n480), .A2(n503), .ZN(n757) );
  XNOR2_X2 U659 ( .A(n543), .B(n559), .ZN(n480) );
  NAND2_X1 U660 ( .A1(n481), .A2(n722), .ZN(n723) );
  XNOR2_X1 U661 ( .A(n721), .B(n720), .ZN(n481) );
  NAND2_X1 U662 ( .A1(n752), .A2(n520), .ZN(n518) );
  NAND2_X1 U663 ( .A1(n487), .A2(n686), .ZN(n485) );
  AND2_X1 U664 ( .A1(n685), .A2(n692), .ZN(n487) );
  NAND2_X1 U665 ( .A1(n491), .A2(n488), .ZN(n828) );
  NAND2_X1 U666 ( .A1(n494), .A2(n493), .ZN(n492) );
  NAND2_X1 U667 ( .A1(n421), .A2(n524), .ZN(n698) );
  INV_X1 U668 ( .A(n715), .ZN(n496) );
  INV_X1 U669 ( .A(n635), .ZN(n497) );
  NAND2_X1 U670 ( .A1(n500), .A2(n826), .ZN(n684) );
  NAND2_X1 U671 ( .A1(n501), .A2(KEYINPUT47), .ZN(n500) );
  NAND2_X1 U672 ( .A1(n771), .A2(n688), .ZN(n501) );
  INV_X1 U673 ( .A(n570), .ZN(n587) );
  NOR2_X1 U674 ( .A1(n711), .A2(n676), .ZN(n682) );
  XNOR2_X2 U675 ( .A(n626), .B(n625), .ZN(n711) );
  XNOR2_X1 U676 ( .A(n586), .B(n585), .ZN(n640) );
  NAND2_X2 U677 ( .A1(n535), .A2(n534), .ZN(n506) );
  NOR2_X1 U678 ( .A1(n505), .A2(n797), .ZN(G63) );
  XNOR2_X2 U679 ( .A(n506), .B(n552), .ZN(n829) );
  XNOR2_X2 U680 ( .A(n614), .B(G469), .ZN(n671) );
  NOR2_X1 U681 ( .A1(n507), .A2(n797), .ZN(G54) );
  NAND2_X1 U682 ( .A1(n828), .A2(n827), .ZN(n673) );
  XNOR2_X1 U683 ( .A(n509), .B(n508), .ZN(G57) );
  NOR2_X2 U684 ( .A1(n763), .A2(n797), .ZN(n509) );
  NOR2_X1 U685 ( .A1(n512), .A2(n797), .ZN(G66) );
  XNOR2_X1 U686 ( .A(n557), .B(n762), .ZN(n763) );
  AND2_X1 U687 ( .A1(n675), .A2(n526), .ZN(n525) );
  XNOR2_X1 U688 ( .A(n530), .B(KEYINPUT95), .ZN(n674) );
  NAND2_X1 U689 ( .A1(n516), .A2(n425), .ZN(n515) );
  INV_X1 U690 ( .A(KEYINPUT121), .ZN(n520) );
  NAND2_X1 U691 ( .A1(n525), .A2(n363), .ZN(n524) );
  NOR2_X1 U692 ( .A1(n529), .A2(n419), .ZN(n526) );
  XNOR2_X2 U693 ( .A(n612), .B(n560), .ZN(n814) );
  INV_X1 U694 ( .A(n637), .ZN(n540) );
  NAND2_X1 U695 ( .A1(n637), .A2(n539), .ZN(n536) );
  NAND2_X1 U696 ( .A1(n694), .A2(n539), .ZN(n537) );
  XNOR2_X2 U697 ( .A(n611), .B(KEYINPUT22), .ZN(n637) );
  NAND2_X1 U698 ( .A1(n561), .A2(n702), .ZN(n703) );
  XNOR2_X2 U699 ( .A(n630), .B(n554), .ZN(n804) );
  INV_X1 U700 ( .A(KEYINPUT65), .ZN(n559) );
  BUF_X1 U701 ( .A(n630), .Z(n631) );
  XOR2_X1 U702 ( .A(n600), .B(n599), .Z(n562) );
  XNOR2_X1 U703 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U704 ( .A(n620), .B(n619), .ZN(n621) );
  INV_X1 U705 ( .A(G116), .ZN(n563) );
  NAND2_X1 U706 ( .A1(n563), .A2(G113), .ZN(n566) );
  NAND2_X1 U707 ( .A1(n564), .A2(G116), .ZN(n565) );
  XNOR2_X2 U708 ( .A(G119), .B(KEYINPUT3), .ZN(n567) );
  XNOR2_X2 U709 ( .A(n568), .B(n567), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G224), .A2(n817), .ZN(n571) );
  XNOR2_X1 U711 ( .A(n576), .B(KEYINPUT73), .ZN(n579) );
  AND2_X1 U712 ( .A1(G210), .A2(n579), .ZN(n577) );
  NAND2_X1 U713 ( .A1(G952), .A2(n817), .ZN(n666) );
  NOR2_X1 U714 ( .A1(G898), .A2(n817), .ZN(n809) );
  NAND2_X1 U715 ( .A1(G902), .A2(n809), .ZN(n580) );
  NAND2_X1 U716 ( .A1(n666), .A2(n580), .ZN(n583) );
  XOR2_X1 U717 ( .A(KEYINPUT14), .B(n581), .Z(n740) );
  INV_X1 U718 ( .A(n740), .ZN(n582) );
  AND2_X1 U719 ( .A1(n583), .A2(n582), .ZN(n584) );
  INV_X1 U720 ( .A(KEYINPUT0), .ZN(n585) );
  XOR2_X1 U721 ( .A(G104), .B(G122), .Z(n589) );
  XNOR2_X1 U722 ( .A(n589), .B(n588), .ZN(n593) );
  XOR2_X1 U723 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n591) );
  XNOR2_X1 U724 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U725 ( .A(n593), .B(n592), .ZN(n596) );
  NOR2_X1 U726 ( .A1(G237), .A2(G953), .ZN(n594) );
  XNOR2_X1 U727 ( .A(n594), .B(KEYINPUT74), .ZN(n628) );
  NAND2_X1 U728 ( .A1(n628), .A2(G214), .ZN(n595) );
  XOR2_X1 U729 ( .A(KEYINPUT13), .B(KEYINPUT100), .Z(n600) );
  XNOR2_X1 U730 ( .A(KEYINPUT101), .B(G475), .ZN(n599) );
  XNOR2_X1 U731 ( .A(G134), .B(KEYINPUT7), .ZN(n603) );
  NAND2_X1 U732 ( .A1(n817), .A2(G234), .ZN(n605) );
  XNOR2_X1 U733 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n604) );
  XNOR2_X1 U734 ( .A(n605), .B(n604), .ZN(n618) );
  NAND2_X1 U735 ( .A1(G217), .A2(n618), .ZN(n606) );
  XNOR2_X1 U736 ( .A(n609), .B(KEYINPUT106), .ZN(n610) );
  NAND2_X1 U737 ( .A1(n640), .A2(n610), .ZN(n611) );
  NAND2_X1 U738 ( .A1(G221), .A2(n618), .ZN(n620) );
  XOR2_X1 U739 ( .A(G119), .B(KEYINPUT23), .Z(n619) );
  XNOR2_X1 U740 ( .A(n622), .B(n621), .ZN(n796) );
  NAND2_X1 U741 ( .A1(n623), .A2(G217), .ZN(n624) );
  NAND2_X1 U742 ( .A1(G210), .A2(n628), .ZN(n629) );
  XNOR2_X1 U743 ( .A(n631), .B(G137), .ZN(n632) );
  XNOR2_X1 U744 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U745 ( .A(G472), .B(KEYINPUT72), .ZN(n635) );
  NOR2_X1 U746 ( .A1(n711), .A2(n638), .ZN(n636) );
  INV_X1 U747 ( .A(n711), .ZN(n657) );
  INV_X1 U748 ( .A(n709), .ZN(n694) );
  INV_X1 U749 ( .A(n681), .ZN(n712) );
  NAND2_X1 U750 ( .A1(n712), .A2(n711), .ZN(n708) );
  BUF_X1 U751 ( .A(n640), .Z(n652) );
  INV_X1 U752 ( .A(n652), .ZN(n650) );
  INV_X1 U753 ( .A(KEYINPUT71), .ZN(n641) );
  NOR2_X1 U754 ( .A1(n645), .A2(n647), .ZN(n677) );
  XNOR2_X1 U755 ( .A(n677), .B(KEYINPUT78), .ZN(n643) );
  INV_X1 U756 ( .A(n645), .ZN(n646) );
  INV_X1 U757 ( .A(n770), .ZN(n780) );
  NAND2_X1 U758 ( .A1(n777), .A2(n780), .ZN(n648) );
  XNOR2_X1 U759 ( .A(KEYINPUT80), .B(n688), .ZN(n655) );
  NAND2_X1 U760 ( .A1(n649), .A2(n715), .ZN(n718) );
  NAND2_X1 U761 ( .A1(n680), .A2(n422), .ZN(n656) );
  NOR2_X1 U762 ( .A1(n657), .A2(n656), .ZN(n764) );
  NAND2_X1 U763 ( .A1(G953), .A2(G902), .ZN(n662) );
  NOR2_X1 U764 ( .A1(n740), .A2(n662), .ZN(n663) );
  XNOR2_X1 U765 ( .A(n663), .B(KEYINPUT109), .ZN(n664) );
  NOR2_X1 U766 ( .A1(G900), .A2(n664), .ZN(n665) );
  XNOR2_X1 U767 ( .A(n665), .B(KEYINPUT110), .ZN(n668) );
  NOR2_X1 U768 ( .A1(n666), .A2(n740), .ZN(n667) );
  NOR2_X1 U769 ( .A1(n668), .A2(n667), .ZN(n676) );
  INV_X1 U770 ( .A(KEYINPUT40), .ZN(n669) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(n731) );
  XOR2_X1 U772 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n670) );
  XOR2_X1 U773 ( .A(KEYINPUT46), .B(KEYINPUT86), .Z(n672) );
  XNOR2_X1 U774 ( .A(n673), .B(n672), .ZN(n686) );
  BUF_X1 U775 ( .A(n678), .Z(n679) );
  NAND2_X1 U776 ( .A1(n428), .A2(n679), .ZN(n774) );
  NOR2_X1 U777 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U778 ( .A1(KEYINPUT80), .A2(n688), .ZN(n690) );
  INV_X1 U779 ( .A(KEYINPUT47), .ZN(n687) );
  NAND2_X1 U780 ( .A1(KEYINPUT80), .A2(n687), .ZN(n689) );
  INV_X1 U781 ( .A(n688), .ZN(n730) );
  NOR2_X1 U782 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U783 ( .A(KEYINPUT43), .B(n695), .Z(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n786) );
  OR2_X1 U785 ( .A1(n780), .A2(n698), .ZN(n785) );
  INV_X1 U786 ( .A(KEYINPUT2), .ZN(n746) );
  OR2_X1 U787 ( .A1(n746), .A2(n699), .ZN(n700) );
  XOR2_X1 U788 ( .A(KEYINPUT91), .B(KEYINPUT67), .Z(n706) );
  XNOR2_X1 U789 ( .A(n704), .B(KEYINPUT59), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n379), .A2(n722), .ZN(n743) );
  AND2_X1 U791 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U792 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U793 ( .A(KEYINPUT49), .B(n713), .Z(n714) );
  NOR2_X1 U794 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U795 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U796 ( .A1(n719), .A2(n718), .ZN(n721) );
  XOR2_X1 U797 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n720) );
  XNOR2_X1 U798 ( .A(n723), .B(KEYINPUT117), .ZN(n737) );
  NOR2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U800 ( .A(n726), .B(KEYINPUT118), .ZN(n727) );
  NOR2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U802 ( .A(KEYINPUT119), .B(n729), .Z(n733) );
  NOR2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U807 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U808 ( .A1(n741), .A2(G952), .ZN(n742) );
  NAND2_X1 U809 ( .A1(n743), .A2(n742), .ZN(n752) );
  NAND2_X1 U810 ( .A1(n816), .A2(n746), .ZN(n744) );
  XNOR2_X1 U811 ( .A(n744), .B(KEYINPUT82), .ZN(n748) );
  BUF_X1 U812 ( .A(n745), .Z(n798) );
  NAND2_X1 U813 ( .A1(n798), .A2(n746), .ZN(n747) );
  NAND2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U815 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U816 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n753) );
  XOR2_X1 U817 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n754) );
  XNOR2_X1 U818 ( .A(n459), .B(n754), .ZN(n756) );
  XNOR2_X1 U819 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U820 ( .A1(n758), .A2(n464), .ZN(n760) );
  INV_X1 U821 ( .A(KEYINPUT56), .ZN(n759) );
  XNOR2_X1 U822 ( .A(n760), .B(n759), .ZN(G51) );
  XOR2_X1 U823 ( .A(G101), .B(n764), .Z(G3) );
  NOR2_X1 U824 ( .A1(n777), .A2(n766), .ZN(n765) );
  XOR2_X1 U825 ( .A(G104), .B(n765), .Z(G6) );
  NOR2_X1 U826 ( .A1(n780), .A2(n766), .ZN(n768) );
  XNOR2_X1 U827 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n767) );
  XNOR2_X1 U828 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U829 ( .A(G107), .B(n769), .ZN(G9) );
  XOR2_X1 U830 ( .A(G128), .B(KEYINPUT29), .Z(n773) );
  NAND2_X1 U831 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U832 ( .A(n773), .B(n772), .ZN(G30) );
  NOR2_X1 U833 ( .A1(n777), .A2(n774), .ZN(n776) );
  XNOR2_X1 U834 ( .A(G146), .B(KEYINPUT113), .ZN(n775) );
  XNOR2_X1 U835 ( .A(n776), .B(n775), .ZN(G48) );
  NOR2_X1 U836 ( .A1(n777), .A2(n779), .ZN(n778) );
  XOR2_X1 U837 ( .A(G113), .B(n778), .Z(G15) );
  NOR2_X1 U838 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U839 ( .A(G116), .B(n781), .Z(G18) );
  XNOR2_X1 U840 ( .A(n782), .B(KEYINPUT114), .ZN(n783) );
  XNOR2_X1 U841 ( .A(n783), .B(KEYINPUT37), .ZN(n784) );
  XNOR2_X1 U842 ( .A(G125), .B(n784), .ZN(G27) );
  XNOR2_X1 U843 ( .A(G134), .B(n785), .ZN(G36) );
  XNOR2_X1 U844 ( .A(G140), .B(n786), .ZN(G42) );
  XNOR2_X1 U845 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n789) );
  XNOR2_X1 U846 ( .A(n787), .B(KEYINPUT57), .ZN(n788) );
  XNOR2_X1 U847 ( .A(n789), .B(n788), .ZN(n791) );
  NAND2_X1 U848 ( .A1(n794), .A2(G469), .ZN(n790) );
  NAND2_X1 U849 ( .A1(G478), .A2(n794), .ZN(n792) );
  NAND2_X1 U850 ( .A1(G217), .A2(n794), .ZN(n795) );
  OR2_X1 U851 ( .A1(G953), .A2(n798), .ZN(n803) );
  NAND2_X1 U852 ( .A1(G224), .A2(G953), .ZN(n799) );
  XNOR2_X1 U853 ( .A(n799), .B(KEYINPUT124), .ZN(n800) );
  XNOR2_X1 U854 ( .A(KEYINPUT61), .B(n800), .ZN(n801) );
  NAND2_X1 U855 ( .A1(n801), .A2(G898), .ZN(n802) );
  NAND2_X1 U856 ( .A1(n803), .A2(n802), .ZN(n811) );
  XNOR2_X1 U857 ( .A(n458), .B(n805), .ZN(n806) );
  XNOR2_X1 U858 ( .A(n806), .B(KEYINPUT125), .ZN(n807) );
  XNOR2_X1 U859 ( .A(n807), .B(G101), .ZN(n808) );
  NOR2_X1 U860 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U861 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U862 ( .A(KEYINPUT126), .B(n812), .ZN(G69) );
  XNOR2_X1 U863 ( .A(n813), .B(KEYINPUT127), .ZN(n815) );
  XOR2_X1 U864 ( .A(n814), .B(n815), .Z(n819) );
  XNOR2_X1 U865 ( .A(n819), .B(n816), .ZN(n818) );
  NAND2_X1 U866 ( .A1(n818), .A2(n817), .ZN(n823) );
  XNOR2_X1 U867 ( .A(G227), .B(n819), .ZN(n820) );
  NAND2_X1 U868 ( .A1(n820), .A2(G900), .ZN(n821) );
  NAND2_X1 U869 ( .A1(n821), .A2(G953), .ZN(n822) );
  NAND2_X1 U870 ( .A1(n823), .A2(n822), .ZN(G72) );
  XOR2_X1 U871 ( .A(n824), .B(G119), .Z(G21) );
  XOR2_X1 U872 ( .A(n825), .B(G122), .Z(G24) );
  XNOR2_X1 U873 ( .A(G143), .B(n826), .ZN(G45) );
  XNOR2_X1 U874 ( .A(n827), .B(G137), .ZN(G39) );
  XNOR2_X1 U875 ( .A(G131), .B(n828), .ZN(G33) );
  XOR2_X1 U876 ( .A(n829), .B(G110), .Z(G12) );
endmodule

