//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT93), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(KEYINPUT93), .A3(new_n204), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n203), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n202), .B2(KEYINPUT94), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G57gat), .A2(G64gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G57gat), .A2(G64gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT94), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(new_n203), .B2(new_n210), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n203), .A2(KEYINPUT93), .A3(new_n204), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT93), .B1(new_n203), .B2(new_n204), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(KEYINPUT21), .ZN(new_n224));
  XOR2_X1   g023(.A(G127gat), .B(G155gat), .Z(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  AOI21_X1  g027(.A(G1gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G22gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G15gat), .ZN(new_n231));
  INV_X1    g030(.A(G15gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G8gat), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n227), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(G1gat), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n236), .A2(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(KEYINPUT21), .B2(new_n223), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n226), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT96), .ZN(new_n247));
  NAND2_X1  g046(.A1(G231gat), .A2(G233gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT95), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n247), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G183gat), .B(G211gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n245), .B(new_n252), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(G232gat), .A2(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT41), .ZN(new_n256));
  XNOR2_X1  g055(.A(G134gat), .B(G162gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G50gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G43gat), .ZN(new_n261));
  INV_X1    g060(.A(G43gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G50gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT15), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT15), .ZN(new_n266));
  OR2_X1    g065(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n268));
  AOI21_X1  g067(.A(G50gat), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT85), .B1(new_n260), .B2(G43gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n262), .A3(G50gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n266), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT14), .B(G29gat), .ZN(new_n275));
  INV_X1    g074(.A(G36gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G29gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n265), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n264), .B1(new_n277), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT17), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT17), .ZN(new_n284));
  INV_X1    g083(.A(new_n282), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n260), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n270), .A3(new_n272), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n289), .A2(new_n266), .B1(new_n277), .B2(new_n279), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n284), .B(new_n285), .C1(new_n290), .C2(new_n265), .ZN(new_n291));
  AND2_X1   g090(.A1(G99gat), .A2(G106gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT97), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G99gat), .ZN(new_n295));
  INV_X1    g094(.A(G106gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT97), .ZN(new_n298));
  NAND2_X1  g097(.A1(G99gat), .A2(G106gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G85gat), .A2(G92gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT7), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G85gat), .A3(G92gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G85gat), .ZN(new_n307));
  INV_X1    g106(.A(G92gat), .ZN(new_n308));
  AOI22_X1  g107(.A1(KEYINPUT8), .A2(new_n299), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n294), .A2(new_n300), .A3(new_n306), .A4(new_n309), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n283), .A2(new_n291), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n274), .A2(new_n280), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n282), .B1(new_n316), .B2(new_n264), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n317), .A2(new_n313), .B1(KEYINPUT41), .B2(new_n255), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G190gat), .B(G218gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT98), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n319), .A2(new_n321), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n259), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n319), .A2(new_n321), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n258), .A3(new_n322), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n254), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n218), .A2(new_n221), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n209), .A2(new_n212), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n313), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT10), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT99), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n213), .A2(new_n222), .A3(new_n312), .A4(new_n311), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n314), .A2(KEYINPUT99), .A3(new_n213), .A4(new_n222), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n340), .B2(new_n334), .ZN(new_n341));
  NAND2_X1  g140(.A1(G230gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT100), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT100), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT10), .B1(new_n338), .B2(new_n339), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n345), .B(new_n342), .C1(new_n346), .C2(new_n335), .ZN(new_n347));
  XOR2_X1   g146(.A(G120gat), .B(G148gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT101), .ZN(new_n349));
  XOR2_X1   g148(.A(G176gat), .B(G204gat), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n340), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n343), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n344), .A2(new_n347), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n343), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n341), .B2(new_n343), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n330), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT65), .ZN(new_n363));
  INV_X1    g162(.A(G190gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n362), .B2(new_n364), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G169gat), .ZN(new_n369));
  INV_X1    g168(.A(G176gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(KEYINPUT26), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n372), .A2(KEYINPUT26), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT1), .B1(new_n379), .B2(KEYINPUT66), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(KEYINPUT66), .B2(new_n379), .ZN(new_n381));
  XOR2_X1   g180(.A(G127gat), .B(G134gat), .Z(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n382), .A2(KEYINPUT1), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n384), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n372), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n371), .B1(new_n392), .B2(new_n375), .ZN(new_n393));
  INV_X1    g192(.A(G183gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n364), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT24), .A3(new_n374), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT25), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n389), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n383), .A2(new_n388), .ZN(new_n401));
  INV_X1    g200(.A(new_n377), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n365), .B2(new_n367), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n397), .B(KEYINPUT25), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n406), .B(KEYINPUT64), .Z(new_n407));
  NAND3_X1  g206(.A1(new_n400), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G15gat), .B(G43gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT68), .ZN(new_n410));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT33), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(KEYINPUT32), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT69), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n408), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n412), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n408), .B2(KEYINPUT32), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n408), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n407), .A2(KEYINPUT34), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n400), .B2(new_n405), .ZN(new_n426));
  INV_X1    g225(.A(new_n400), .ZN(new_n427));
  INV_X1    g226(.A(new_n405), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n406), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n429), .B2(KEYINPUT34), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n416), .A2(new_n417), .B1(new_n422), .B2(new_n420), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n424), .A2(new_n438), .A3(new_n431), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT70), .B1(new_n433), .B2(new_n430), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT36), .A4(new_n434), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n403), .A2(new_n404), .ZN(new_n445));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT73), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n378), .A2(new_n399), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT74), .A3(new_n447), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n445), .B2(KEYINPUT29), .ZN(new_n452));
  XNOR2_X1  g251(.A(G197gat), .B(G204gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT22), .ZN(new_n454));
  INV_X1    g253(.A(G211gat), .ZN(new_n455));
  INV_X1    g254(.A(G218gat), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(G211gat), .B(G218gat), .Z(new_n459));
  OR2_X1    g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(KEYINPUT71), .A3(new_n459), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT72), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT72), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n467), .A3(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n447), .B1(new_n450), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n445), .A2(new_n446), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT81), .B(KEYINPUT37), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT75), .ZN(new_n479));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n479), .B(new_n480), .Z(new_n481));
  AND2_X1   g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n448), .B1(new_n445), .B2(KEYINPUT29), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n446), .B2(new_n445), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n485), .B2(new_n469), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n471), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT38), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n475), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n481), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n482), .A2(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493));
  OR2_X1    g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(KEYINPUT2), .ZN(new_n495));
  INV_X1    g294(.A(G141gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G148gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(G148gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(KEYINPUT76), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n500), .A2(new_n496), .A3(G148gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G141gat), .B(G148gat), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n493), .B(new_n494), .C1(new_n503), .C2(KEYINPUT2), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n401), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT77), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n389), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n383), .A2(KEYINPUT77), .A3(new_n388), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(KEYINPUT3), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n517));
  NOR3_X1   g316(.A1(new_n389), .A2(new_n505), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g319(.A1(G225gat), .A2(G233gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n509), .A2(new_n516), .A3(new_n519), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n518), .B1(new_n508), .B2(new_n507), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(KEYINPUT80), .A3(new_n516), .A4(new_n523), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n522), .B1(new_n507), .B2(new_n517), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n389), .A2(new_n505), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT4), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n516), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n511), .A2(new_n512), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n531), .B1(new_n534), .B2(new_n505), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n533), .B(new_n520), .C1(new_n535), .C2(new_n521), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G1gat), .B(G29gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT0), .ZN(new_n539));
  XNOR2_X1  g338(.A(G57gat), .B(G85gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n536), .A3(new_n541), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n492), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT82), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n492), .A2(new_n546), .A3(new_n550), .A4(new_n547), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n482), .B1(new_n483), .B2(new_n490), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT38), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G22gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n515), .A2(new_n472), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n466), .A2(new_n557), .A3(new_n468), .ZN(new_n558));
  NAND2_X1  g357(.A1(G228gat), .A2(G233gat), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT29), .B1(new_n460), .B2(new_n462), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n505), .B1(new_n560), .B2(KEYINPUT3), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n463), .A2(new_n472), .A3(new_n464), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n514), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n505), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n559), .B1(new_n558), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G50gat), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n562), .B2(new_n566), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n556), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  INV_X1    g371(.A(new_n556), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n572), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n521), .B1(new_n527), .B2(new_n516), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n542), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n535), .A2(new_n521), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n543), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n583), .B2(new_n582), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n489), .B2(new_n481), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n489), .B2(new_n481), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n490), .A2(new_n586), .A3(new_n491), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n576), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n443), .B1(new_n554), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n546), .A2(new_n547), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n576), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n573), .B1(new_n572), .B2(new_n568), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n569), .A2(new_n570), .A3(new_n556), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n434), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT83), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n440), .A4(new_n439), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n439), .A2(new_n440), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n434), .A2(new_n597), .A3(new_n598), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT83), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n546), .A2(new_n547), .B1(new_n588), .B2(new_n589), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n607));
  INV_X1    g406(.A(new_n435), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n571), .A2(new_n574), .A3(KEYINPUT35), .ZN(new_n609));
  AND4_X1   g408(.A1(new_n594), .A2(new_n608), .A3(new_n590), .A4(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n593), .A2(new_n596), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n236), .A2(new_n238), .ZN(new_n615));
  INV_X1    g414(.A(new_n229), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n283), .A2(new_n291), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n285), .B1(new_n290), .B2(new_n265), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n621), .A2(new_n619), .A3(KEYINPUT87), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n317), .B2(new_n243), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n614), .B(new_n620), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT18), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT87), .B1(new_n621), .B2(new_n619), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n317), .A2(new_n243), .A3(new_n623), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n627), .A2(new_n628), .B1(new_n621), .B2(new_n619), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT13), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n625), .A2(new_n626), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(KEYINPUT88), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n628), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT88), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n614), .A4(new_n620), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G197gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT11), .B(G169gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n638), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n625), .B2(KEYINPUT88), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n632), .B1(new_n637), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT90), .B1(new_n650), .B2(new_n645), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n633), .A2(new_n639), .A3(KEYINPUT90), .A4(new_n645), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n633), .A2(new_n639), .A3(new_n645), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT90), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n658), .A2(new_n652), .B1(new_n646), .B2(new_n640), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n613), .A2(KEYINPUT92), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT92), .ZN(new_n664));
  INV_X1    g463(.A(new_n662), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n612), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n361), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n594), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AND3_X1   g470(.A1(new_n667), .A2(new_n591), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n237), .B1(new_n667), .B2(new_n591), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  INV_X1    g474(.A(new_n667), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n676), .B2(new_n442), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n232), .A3(new_n608), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n667), .A2(new_n576), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  AOI21_X1  g481(.A(KEYINPUT102), .B1(new_n595), .B2(new_n576), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n605), .A2(new_n684), .A3(new_n575), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n554), .A2(new_n592), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT103), .A4(new_n442), .ZN(new_n688));
  AOI211_X1 g487(.A(KEYINPUT104), .B(new_n610), .C1(new_n606), .C2(KEYINPUT35), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n607), .B2(new_n611), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT103), .B1(new_n593), .B2(new_n686), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n328), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n613), .A2(KEYINPUT44), .A3(new_n328), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n659), .A2(new_n254), .A3(new_n359), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n594), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n663), .A2(new_n666), .ZN(new_n702));
  INV_X1    g501(.A(new_n359), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n253), .A2(new_n328), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G29gat), .A3(new_n594), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n701), .A2(new_n708), .A3(new_n709), .ZN(G1328gat));
  OAI21_X1  g509(.A(G36gat), .B1(new_n700), .B2(new_n590), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n706), .A2(G36gat), .A3(new_n590), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n696), .A2(new_n443), .A3(new_n697), .A4(new_n699), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n286), .A2(new_n287), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n702), .A2(new_n608), .A3(new_n718), .A4(new_n705), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n720), .B(new_n723), .C1(new_n721), .C2(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n702), .A2(new_n576), .A3(new_n705), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(new_n260), .B1(new_n730), .B2(KEYINPUT48), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n730), .A2(KEYINPUT48), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n575), .A2(new_n260), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n696), .A2(new_n697), .A3(new_n699), .A4(new_n733), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n732), .B1(new_n731), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  NAND2_X1  g536(.A1(new_n593), .A2(new_n686), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n740), .B(new_n688), .C1(new_n689), .C2(new_n691), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n659), .A2(new_n254), .A3(new_n329), .A4(new_n359), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n668), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n591), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n443), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G71gat), .ZN(new_n752));
  INV_X1    g551(.A(G71gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n744), .A2(new_n753), .A3(new_n608), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n744), .A2(new_n576), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n654), .A2(new_n254), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT107), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n359), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n698), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n594), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n328), .B(new_n761), .C1(new_n692), .C2(new_n693), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n741), .A2(KEYINPUT51), .A3(new_n328), .A4(new_n761), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n703), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n307), .A3(new_n668), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n770), .ZN(G1336gat));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n768), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n590), .A2(G92gat), .A3(new_n703), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n696), .A2(new_n591), .A3(new_n697), .A4(new_n762), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n776), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n780), .B(new_n776), .C1(new_n777), .C2(new_n772), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1337gat));
  XNOR2_X1  g583(.A(KEYINPUT110), .B(G99gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n608), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n763), .A2(new_n442), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n785), .ZN(G1338gat));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n296), .A3(new_n576), .A4(new_n359), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n696), .A2(new_n576), .A3(new_n697), .A4(new_n762), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G106gat), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n789), .B2(new_n791), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n341), .B2(new_n343), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n344), .A2(new_n798), .A3(new_n347), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n797), .B(new_n342), .C1(new_n346), .C2(new_n335), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n352), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n799), .A2(new_n804), .A3(KEYINPUT55), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n644), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n635), .A2(new_n620), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(G229gat), .A3(G233gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n629), .A2(new_n631), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n658), .B2(new_n652), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(new_n799), .B2(new_n801), .ZN(new_n813));
  INV_X1    g612(.A(new_n355), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n806), .A2(new_n328), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT113), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n811), .B(new_n329), .C1(new_n658), .C2(new_n652), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n806), .A4(new_n815), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n654), .A3(new_n815), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n812), .A2(new_n359), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n328), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n796), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n329), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(KEYINPUT114), .A3(new_n817), .A4(new_n820), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n828), .A3(new_n253), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n361), .A2(new_n654), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n576), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n591), .A2(new_n594), .A3(new_n435), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n665), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n594), .B1(new_n829), .B2(new_n831), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n601), .A2(new_n604), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n591), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n659), .A2(G113gat), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT115), .Z(new_n841));
  OAI21_X1  g640(.A(new_n835), .B1(new_n839), .B2(new_n841), .ZN(G1340gat));
  INV_X1    g641(.A(new_n834), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(G120gat), .A3(new_n359), .ZN(new_n844));
  INV_X1    g643(.A(G120gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n839), .B2(new_n703), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(G1341gat));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n254), .A2(G127gat), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n834), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n834), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n839), .A2(new_n253), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n850), .B(new_n851), .C1(G127gat), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT117), .ZN(G1342gat));
  OR2_X1    g653(.A1(new_n329), .A2(G134gat), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n839), .A2(KEYINPUT56), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n834), .B2(new_n329), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT56), .B1(new_n839), .B2(new_n855), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT118), .Z(G1343gat));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n443), .A2(new_n594), .A3(new_n591), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n575), .B1(new_n829), .B2(new_n831), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(KEYINPUT57), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n576), .A2(KEYINPUT57), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n806), .A2(new_n815), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n655), .B2(new_n661), .ZN(new_n868));
  INV_X1    g667(.A(new_n823), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n329), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n817), .A2(new_n820), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n254), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n830), .B1(new_n872), .B2(KEYINPUT119), .ZN(new_n873));
  INV_X1    g672(.A(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n662), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n328), .B1(new_n875), .B2(new_n823), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n253), .B1(new_n876), .B2(new_n821), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n866), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n654), .B(new_n863), .C1(new_n865), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G141gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n443), .A2(new_n575), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n590), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n665), .A2(G141gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n836), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n862), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n862), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n662), .B(new_n863), .C1(new_n865), .C2(new_n880), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(G141gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n861), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(G141gat), .ZN(new_n894));
  INV_X1    g693(.A(new_n890), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n836), .A2(new_n886), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n881), .A2(G141gat), .B1(new_n898), .B2(new_n887), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n896), .B(KEYINPUT121), .C1(new_n862), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n665), .A2(new_n360), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT122), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n254), .B1(new_n870), .B2(new_n816), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n903), .B(new_n576), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n863), .A2(new_n359), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n907), .B(new_n908), .C1(new_n864), .C2(new_n903), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n902), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n359), .B(new_n863), .C1(new_n865), .C2(new_n880), .ZN(new_n911));
  INV_X1    g710(.A(G148gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(KEYINPUT59), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n897), .A2(G148gat), .A3(new_n703), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT123), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  INV_X1    g716(.A(new_n915), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n911), .A2(new_n913), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n910), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(new_n863), .B1(new_n865), .B2(new_n880), .ZN(new_n922));
  OAI21_X1  g721(.A(G155gat), .B1(new_n922), .B2(new_n253), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n253), .A2(G155gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n897), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n922), .B2(new_n329), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n329), .A2(G162gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n897), .B2(new_n927), .ZN(G1347gat));
  AOI21_X1  g727(.A(new_n668), .B1(new_n829), .B2(new_n831), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n837), .A2(new_n590), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n654), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n668), .A2(new_n590), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n832), .A2(new_n608), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n665), .A2(new_n369), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  NOR3_X1   g736(.A1(new_n931), .A2(G176gat), .A3(new_n703), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n359), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(G176gat), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT124), .ZN(G1349gat));
  AND4_X1   g740(.A1(new_n363), .A2(new_n929), .A3(new_n254), .A4(new_n930), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n935), .A2(new_n254), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(G183gat), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n364), .A3(new_n328), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n935), .A2(new_n328), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G190gat), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  AND3_X1   g750(.A1(new_n929), .A2(new_n591), .A3(new_n883), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n654), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n442), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT125), .Z(new_n955));
  OAI211_X1 g754(.A(new_n907), .B(new_n955), .C1(new_n864), .C2(new_n903), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n662), .A2(G197gat), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n953), .A2(G197gat), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n952), .A2(new_n960), .A3(new_n359), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n956), .A2(new_n963), .A3(new_n703), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n956), .B2(new_n703), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n964), .B2(new_n966), .ZN(G1353gat));
  OAI21_X1  g766(.A(G211gat), .B1(new_n956), .B2(new_n253), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n455), .A3(new_n254), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n956), .B2(new_n329), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n952), .A2(new_n456), .A3(new_n328), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT127), .Z(G1355gat));
endmodule


