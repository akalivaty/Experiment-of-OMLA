//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT7), .ZN(new_n205));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206));
  INV_X1    g005(.A(G85gat), .ZN(new_n207));
  INV_X1    g006(.A(G92gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(KEYINPUT8), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G99gat), .B(G106gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT94), .A2(G57gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(G64gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G71gat), .A2(G78gat), .ZN(new_n215));
  OR2_X1    g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n220));
  AND2_X1   g019(.A1(G57gat), .A2(G64gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n215), .B(new_n216), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n212), .B(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT10), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n212), .A2(KEYINPUT10), .A3(new_n219), .A4(new_n222), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n203), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n224), .A2(new_n202), .ZN(new_n230));
  XOR2_X1   g029(.A(G120gat), .B(G148gat), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT97), .ZN(new_n232));
  XNOR2_X1  g031(.A(G176gat), .B(G204gat), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n232), .B(new_n233), .Z(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(KEYINPUT98), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n228), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n230), .ZN(new_n241));
  INV_X1    g040(.A(new_n234), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n236), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT15), .ZN(new_n244));
  XNOR2_X1  g043(.A(G43gat), .B(G50gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT90), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(KEYINPUT90), .B2(new_n245), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n245), .A2(KEYINPUT15), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT91), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G29gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT14), .B(G29gat), .Z(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(G36gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(KEYINPUT91), .B2(new_n248), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n250), .A2(new_n254), .B1(new_n255), .B2(new_n247), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(new_n212), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT95), .ZN(new_n262));
  AND2_X1   g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n256), .A2(new_n212), .B1(KEYINPUT41), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n264), .A2(new_n262), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT96), .ZN(new_n267));
  XNOR2_X1  g066(.A(G190gat), .B(G218gat), .ZN(new_n268));
  OAI22_X1  g067(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n267), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n263), .A2(KEYINPUT41), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G134gat), .B(G162gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n269), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n223), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G231gat), .A2(G233gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G127gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G22gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT92), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G1gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n286), .A2(KEYINPUT16), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(G8gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n277), .B2(new_n223), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n282), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G155gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n243), .A2(new_n276), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT93), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G127gat), .A2(G134gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  INV_X1    g108(.A(G120gat), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT1), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(KEYINPUT72), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G120gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n309), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n304), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G113gat), .B2(G120gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n307), .B2(new_n306), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n314), .A2(G120gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n310), .A2(KEYINPUT72), .ZN(new_n322));
  OAI21_X1  g121(.A(G113gat), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n323), .A3(KEYINPUT73), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT71), .B(G127gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n311), .A2(new_n327), .B1(new_n281), .B2(new_n305), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n317), .A2(new_n324), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G141gat), .B(G148gat), .ZN(new_n335));
  AND2_X1   g134(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n338));
  INV_X1    g137(.A(G148gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(G141gat), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT80), .B1(new_n341), .B2(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(G148gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n330), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n332), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT81), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G162gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n348), .B1(new_n353), .B2(G155gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n337), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n329), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n328), .A2(new_n326), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n312), .A2(new_n316), .A3(new_n304), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT73), .B1(new_n320), .B2(new_n323), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n355), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n303), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n337), .B(new_n370), .C1(new_n347), .C2(new_n354), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n329), .A2(new_n356), .A3(KEYINPUT4), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n368), .A2(new_n372), .A3(new_n364), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n361), .B2(new_n355), .ZN(new_n377));
  INV_X1    g176(.A(new_n367), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n329), .A2(new_n356), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n377), .A2(new_n372), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n375), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G1gat), .B(G29gat), .Z(new_n386));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n385), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n390), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(KEYINPUT84), .A3(new_n372), .A4(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n382), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n396), .A2(new_n397), .B1(new_n366), .B2(new_n374), .ZN(new_n398));
  INV_X1    g197(.A(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT6), .B1(new_n385), .B2(new_n390), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n393), .A2(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G226gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G169gat), .ZN(new_n406));
  INV_X1    g205(.A(G176gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT26), .ZN(new_n409));
  NAND2_X1  g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT65), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT65), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(G169gat), .A3(G176gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n415), .A2(new_n406), .A3(new_n407), .A4(KEYINPUT70), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n420));
  AND2_X1   g219(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT27), .B(G183gat), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n426));
  INV_X1    g225(.A(G183gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT27), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G183gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n431));
  AND4_X1   g230(.A1(new_n426), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n425), .A2(KEYINPUT69), .B1(new_n432), .B2(KEYINPUT28), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n426), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n434));
  XOR2_X1   g233(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n419), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT24), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT64), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT23), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n406), .A3(new_n407), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n446), .A2(new_n448), .B1(new_n411), .B2(new_n413), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n441), .A2(new_n442), .A3(new_n450), .A4(new_n443), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT66), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT24), .B1(new_n418), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n454), .B2(new_n418), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n423), .A2(new_n427), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n443), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n446), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n459), .A2(new_n414), .A3(KEYINPUT25), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n452), .A2(new_n453), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n405), .B1(new_n439), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n460), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n417), .A2(new_n418), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT28), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n436), .B2(new_n437), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n425), .A2(KEYINPUT69), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n462), .B1(new_n471), .B2(new_n405), .ZN(new_n472));
  XNOR2_X1  g271(.A(G197gat), .B(G204gat), .ZN(new_n473));
  INV_X1    g272(.A(G211gat), .ZN(new_n474));
  INV_X1    g273(.A(G218gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n473), .B1(KEYINPUT22), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G211gat), .B(G218gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n479), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n462), .B(new_n481), .C1(new_n471), .C2(new_n405), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G8gat), .B(G36gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G64gat), .B(G92gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n480), .A2(new_n486), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT30), .A3(new_n489), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n483), .A2(KEYINPUT30), .A3(new_n487), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT87), .B1(new_n402), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  XOR2_X1   g293(.A(G15gat), .B(G43gat), .Z(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT74), .B1(new_n439), .B2(new_n461), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT74), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n465), .A2(new_n470), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n361), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT74), .B(new_n329), .C1(new_n439), .C2(new_n461), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT33), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(KEYINPUT32), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(KEYINPUT32), .C1(new_n508), .C2(new_n499), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n506), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n504), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n514), .A2(new_n518), .A3(new_n515), .A4(new_n504), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n504), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n515), .B1(new_n514), .B2(new_n504), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(KEYINPUT77), .B2(new_n516), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n525), .A2(new_n511), .A3(new_n512), .A4(new_n519), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n481), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n356), .B1(new_n528), .B2(new_n370), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n481), .B1(new_n527), .B2(new_n371), .ZN(new_n530));
  XNOR2_X1  g329(.A(G78gat), .B(G106gat), .ZN(new_n531));
  OR3_X1    g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n529), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g332(.A1(G228gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G22gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G50gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  AND3_X1   g336(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n532), .B2(new_n533), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND4_X1   g339(.A1(new_n494), .A2(new_n523), .A3(new_n526), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n401), .A2(new_n400), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n396), .A2(new_n397), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n399), .B1(new_n543), .B2(new_n375), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT85), .B1(new_n544), .B2(KEYINPUT6), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT6), .ZN(new_n546));
  NOR4_X1   g345(.A1(new_n398), .A2(new_n392), .A3(new_n546), .A4(new_n399), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n490), .A2(new_n491), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n493), .A2(new_n541), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n542), .A2(new_n391), .B1(new_n491), .B2(new_n490), .ZN(new_n554));
  INV_X1    g353(.A(new_n522), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(KEYINPUT78), .B2(new_n513), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n513), .A2(KEYINPUT78), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(new_n522), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n540), .B(new_n554), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n552), .A2(new_n553), .B1(new_n559), .B2(KEYINPUT35), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n493), .A2(new_n541), .A3(new_n551), .A4(KEYINPUT88), .ZN(new_n561));
  INV_X1    g360(.A(new_n540), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n377), .A2(new_n372), .A3(new_n379), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT39), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n365), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n565), .A2(new_n399), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n365), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n567), .B(KEYINPUT39), .C1(new_n365), .C2(new_n363), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT40), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT40), .B1(new_n566), .B2(new_n568), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n569), .A2(new_n570), .A3(new_n544), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n562), .B1(new_n492), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n489), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n480), .A2(new_n482), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT38), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n486), .B1(new_n483), .B2(KEYINPUT37), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n578), .B(new_n542), .C1(new_n545), .C2(new_n547), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT38), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n483), .A2(KEYINPUT37), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n487), .B1(new_n574), .B2(new_n575), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(KEYINPUT86), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT86), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n572), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n542), .A2(new_n391), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n562), .B1(new_n589), .B2(new_n492), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n523), .A2(new_n526), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(KEYINPUT36), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n522), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n555), .A2(KEYINPUT78), .A3(new_n513), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT36), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n560), .A2(new_n561), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n291), .A2(new_n258), .A3(new_n259), .ZN(new_n600));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n289), .B(G8gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n256), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT18), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n602), .B(new_n256), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n601), .B(KEYINPUT13), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n605), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n606), .A2(new_n609), .A3(new_n610), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n302), .B1(new_n599), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n552), .A2(new_n553), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n559), .A2(KEYINPUT35), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n561), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n587), .A2(new_n596), .A3(new_n593), .A4(new_n590), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(KEYINPUT93), .A3(new_n621), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n301), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n589), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT16), .B(G8gat), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n633), .A2(new_n549), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n290), .B1(new_n630), .B2(new_n492), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT42), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(KEYINPUT42), .B2(new_n636), .ZN(G1325gat));
  OR3_X1    g438(.A1(new_n633), .A2(G15gat), .A3(new_n592), .ZN(new_n640));
  OAI21_X1  g439(.A(G15gat), .B1(new_n633), .B2(new_n598), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(G1326gat));
  NAND2_X1  g441(.A1(new_n630), .A2(new_n562), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT43), .B(G22gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n243), .B(KEYINPUT99), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n648), .A2(new_n622), .A3(new_n300), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n628), .B2(new_n275), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n276), .B(new_n653), .C1(new_n626), .C2(new_n627), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n589), .B(new_n649), .C1(new_n651), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT44), .B1(new_n599), .B2(new_n276), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n628), .A2(new_n275), .A3(new_n652), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n589), .A4(new_n649), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n656), .A2(G29gat), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663));
  INV_X1    g462(.A(new_n243), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n664), .A2(new_n276), .A3(new_n300), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT93), .B1(new_n628), .B2(new_n621), .ZN(new_n666));
  AOI211_X1 g465(.A(new_n302), .B(new_n622), .C1(new_n626), .C2(new_n627), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n589), .A2(new_n251), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n665), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n623), .B2(new_n629), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n672), .A2(KEYINPUT45), .A3(new_n251), .A4(new_n589), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n646), .B1(new_n662), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n661), .A3(G29gat), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n670), .A4(new_n673), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(G1328gat));
  NOR3_X1   g477(.A1(new_n668), .A2(G36gat), .A3(new_n549), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  INV_X1    g479(.A(G36gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n659), .A2(new_n492), .A3(new_n649), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n683), .B2(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(G1329gat));
  OAI211_X1 g485(.A(new_n597), .B(new_n649), .C1(new_n651), .C2(new_n654), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G43gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n592), .A2(G43gat), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n665), .B(new_n689), .C1(new_n666), .C2(new_n667), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n672), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(KEYINPUT104), .A2(new_n690), .B1(new_n687), .B2(G43gat), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n699), .A2(KEYINPUT105), .A3(new_n695), .A4(new_n693), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(G1330gat));
  OAI211_X1 g500(.A(new_n562), .B(new_n649), .C1(new_n651), .C2(new_n654), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n702), .A2(new_n703), .A3(G50gat), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n702), .B2(G50gat), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n668), .A2(G50gat), .A3(new_n540), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n702), .A2(G50gat), .ZN(new_n711));
  OAI22_X1  g510(.A1(new_n707), .A2(new_n708), .B1(new_n710), .B2(new_n711), .ZN(G1331gat));
  NAND3_X1  g511(.A1(new_n622), .A2(new_n300), .A3(new_n276), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n599), .A2(new_n647), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n589), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n492), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT49), .B(G64gat), .Z(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(G1333gat));
  NAND2_X1  g519(.A1(new_n714), .A2(new_n597), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n592), .A2(G71gat), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n721), .A2(G71gat), .B1(new_n714), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n562), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n621), .A2(new_n300), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n628), .A2(new_n275), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n732), .A2(new_n207), .A3(new_n589), .A4(new_n664), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n664), .B(new_n727), .C1(new_n651), .C2(new_n654), .ZN(new_n734));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734), .B2(new_n588), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n734), .B2(new_n549), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n628), .A2(new_n275), .A3(new_n727), .A4(new_n731), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n647), .A2(G92gat), .A3(new_n549), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT109), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n740), .C1(new_n728), .C2(new_n729), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT52), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n737), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1337gat));
  NOR3_X1   g547(.A1(new_n243), .A2(new_n592), .A3(G99gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G99gat), .B1(new_n734), .B2(new_n598), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1338gat));
  OAI21_X1  g551(.A(G106gat), .B1(new_n734), .B2(new_n540), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n647), .A2(G106gat), .A3(new_n540), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n738), .B(new_n754), .C1(new_n728), .C2(new_n729), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1339gat));
  INV_X1    g557(.A(new_n300), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n237), .A2(new_n760), .A3(new_n239), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n228), .A2(new_n760), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n226), .A2(new_n203), .A3(new_n227), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(KEYINPUT113), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT113), .B1(new_n762), .B2(new_n763), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n242), .B(new_n761), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n762), .A2(new_n763), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n764), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(KEYINPUT55), .A3(new_n242), .A4(new_n761), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n769), .A2(new_n774), .A3(new_n621), .A4(new_n235), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n607), .A2(new_n608), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n601), .B1(new_n600), .B2(new_n603), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n616), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n616), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n620), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(new_n243), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n275), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n235), .A3(new_n774), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(new_n276), .A3(new_n782), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n759), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n301), .A2(new_n621), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n592), .A2(new_n562), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n588), .A2(new_n492), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G113gat), .B1(new_n792), .B2(new_n622), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n562), .B1(new_n594), .B2(new_n595), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n789), .A2(new_n589), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n588), .B1(new_n787), .B2(new_n788), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n797), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n549), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n621), .A2(new_n309), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n795), .A2(new_n796), .B1(new_n804), .B2(new_n805), .ZN(G1340gat));
  OAI21_X1  g605(.A(G120gat), .B1(new_n792), .B2(new_n647), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(KEYINPUT117), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(KEYINPUT117), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n664), .A2(new_n313), .A3(new_n315), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n808), .A2(new_n809), .B1(new_n804), .B2(new_n810), .ZN(G1341gat));
  OAI21_X1  g610(.A(new_n325), .B1(new_n792), .B2(new_n759), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n759), .A2(new_n325), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n804), .B2(new_n813), .ZN(G1342gat));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n276), .A2(new_n492), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(G134gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G134gat), .B1(new_n792), .B2(new_n276), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n818), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(KEYINPUT56), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT118), .B(new_n815), .C1(new_n803), .C2(new_n818), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n819), .B(new_n820), .C1(new_n823), .C2(new_n824), .ZN(G1343gat));
  NOR3_X1   g624(.A1(new_n597), .A2(new_n588), .A3(new_n492), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n540), .B1(new_n787), .B2(new_n788), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  XOR2_X1   g630(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n832));
  NAND2_X1  g631(.A1(new_n767), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n774), .A3(new_n621), .A4(new_n235), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n275), .B1(new_n834), .B2(new_n783), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n759), .B1(new_n835), .B2(new_n786), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n831), .B(new_n540), .C1(new_n836), .C2(new_n788), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n826), .B(new_n621), .C1(new_n830), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n789), .A2(new_n791), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n598), .A2(new_n562), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n622), .A2(G141gat), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n838), .A2(G141gat), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g642(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(G1344gat));
  OAI211_X1 g644(.A(new_n826), .B(new_n664), .C1(new_n830), .C2(new_n837), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n339), .A2(KEYINPUT59), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(KEYINPUT123), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n826), .A2(new_n664), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n540), .B1(new_n836), .B2(new_n788), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n789), .A2(new_n562), .A3(new_n829), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n856), .B2(new_n339), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n339), .A3(new_n664), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT122), .Z(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1345gat));
  OAI21_X1  g660(.A(new_n826), .B1(new_n830), .B2(new_n837), .ZN(new_n862));
  OAI21_X1  g661(.A(G155gat), .B1(new_n862), .B2(new_n759), .ZN(new_n863));
  INV_X1    g662(.A(G155gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n864), .A3(new_n300), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1346gat));
  OAI21_X1  g665(.A(new_n353), .B1(new_n862), .B2(new_n276), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n840), .A2(new_n353), .A3(new_n817), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n800), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n589), .A2(new_n549), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n787), .B2(new_n788), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n797), .ZN(new_n874));
  AOI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n621), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n790), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n406), .A3(new_n622), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n874), .B2(new_n664), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n873), .A2(G176gat), .A3(new_n790), .A4(new_n648), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(KEYINPUT124), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(KEYINPUT124), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(G1349gat));
  NAND3_X1  g682(.A1(new_n874), .A2(new_n424), .A3(new_n300), .ZN(new_n884));
  OAI21_X1  g683(.A(G183gat), .B1(new_n876), .B2(new_n759), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n874), .A2(new_n423), .A3(new_n275), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT125), .Z(new_n889));
  OAI21_X1  g688(.A(G190gat), .B1(new_n876), .B2(new_n276), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(G1351gat));
  NOR2_X1   g693(.A1(new_n597), .A2(new_n872), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n855), .B1(KEYINPUT57), .B2(new_n853), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(KEYINPUT126), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n855), .B(new_n899), .C1(KEYINPUT57), .C2(new_n853), .ZN(new_n900));
  AND4_X1   g699(.A1(G197gat), .A2(new_n898), .A3(new_n621), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n827), .A2(new_n895), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G197gat), .B1(new_n903), .B2(new_n621), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n904), .ZN(G1352gat));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n648), .A3(new_n900), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G204gat), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n902), .A2(G204gat), .A3(new_n243), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT62), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1353gat));
  NAND3_X1  g709(.A1(new_n903), .A2(new_n474), .A3(new_n300), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n897), .A2(new_n300), .A3(new_n895), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n912), .B2(G211gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1354gat));
  NOR2_X1   g714(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n916));
  AOI211_X1 g715(.A(new_n540), .B(new_n828), .C1(new_n787), .C2(new_n788), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT126), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n276), .A2(new_n475), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n895), .A3(new_n900), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n475), .B1(new_n902), .B2(new_n276), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(KEYINPUT127), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1355gat));
endmodule


