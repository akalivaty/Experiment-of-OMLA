

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U321 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U322 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U323 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U324 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U325 ( .A(n415), .B(KEYINPUT41), .Z(n557) );
  XOR2_X1 U326 ( .A(n305), .B(n304), .Z(n514) );
  XNOR2_X1 U327 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U328 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(G176GAT), .B(KEYINPUT17), .Z(n290) );
  XNOR2_X1 U330 ( .A(KEYINPUT84), .B(KEYINPUT18), .ZN(n289) );
  XNOR2_X1 U331 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U332 ( .A(n291), .B(KEYINPUT19), .Z(n293) );
  XNOR2_X1 U333 ( .A(G183GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n335) );
  XOR2_X1 U335 ( .A(KEYINPUT82), .B(G134GAT), .Z(n295) );
  XNOR2_X1 U336 ( .A(G127GAT), .B(G120GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(KEYINPUT0), .B(n296), .Z(n323) );
  XNOR2_X1 U339 ( .A(n335), .B(n323), .ZN(n305) );
  XOR2_X1 U340 ( .A(G15GAT), .B(G113GAT), .Z(n298) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G43GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n347) );
  XOR2_X1 U343 ( .A(n347), .B(KEYINPUT83), .Z(n300) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(n301), .B(KEYINPUT20), .Z(n303) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G71GAT), .ZN(n369) );
  XOR2_X1 U348 ( .A(n369), .B(KEYINPUT85), .Z(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  INV_X1 U350 ( .A(n514), .ZN(n524) );
  XOR2_X1 U351 ( .A(KEYINPUT1), .B(G1GAT), .Z(n307) );
  XNOR2_X1 U352 ( .A(G29GAT), .B(G113GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U354 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT89), .B(KEYINPUT4), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U357 ( .A(n311), .B(n310), .Z(n321) );
  XNOR2_X1 U358 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n312), .B(KEYINPUT87), .ZN(n313) );
  XOR2_X1 U360 ( .A(n313), .B(KEYINPUT3), .Z(n315) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(G162GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n441) );
  XNOR2_X1 U363 ( .A(G148GAT), .B(G85GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n316), .B(G57GAT), .ZN(n359) );
  XOR2_X1 U365 ( .A(n359), .B(KEYINPUT6), .Z(n318) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n441), .B(n319), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n459) );
  XNOR2_X1 U371 ( .A(KEYINPUT91), .B(n459), .ZN(n509) );
  XOR2_X1 U372 ( .A(G92GAT), .B(G64GAT), .Z(n362) );
  XOR2_X1 U373 ( .A(G204GAT), .B(G8GAT), .Z(n325) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G36GAT), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U376 ( .A(n362), .B(n326), .Z(n328) );
  NAND2_X1 U377 ( .A1(G226GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U379 ( .A(n329), .B(KEYINPUT92), .Z(n333) );
  XOR2_X1 U380 ( .A(G211GAT), .B(KEYINPUT21), .Z(n331) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(G218GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n428) );
  XNOR2_X1 U383 ( .A(n428), .B(KEYINPUT93), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n511) );
  INV_X1 U386 ( .A(n511), .ZN(n424) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(KEYINPUT69), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n336), .B(G29GAT), .ZN(n337) );
  XOR2_X1 U389 ( .A(n337), .B(KEYINPUT7), .Z(n339) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n378) );
  XOR2_X1 U392 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n341) );
  XNOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U395 ( .A(G141GAT), .B(G197GAT), .Z(n343) );
  NAND2_X1 U396 ( .A1(G229GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U398 ( .A(n345), .B(n344), .Z(n349) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(G1GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n346), .B(G8GAT), .ZN(n397) );
  XNOR2_X1 U401 ( .A(n347), .B(n397), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U403 ( .A(n378), .B(n350), .Z(n567) );
  XOR2_X1 U404 ( .A(KEYINPUT71), .B(n567), .Z(n552) );
  XOR2_X1 U405 ( .A(G106GAT), .B(KEYINPUT73), .Z(n374) );
  XOR2_X1 U406 ( .A(G204GAT), .B(G78GAT), .Z(n427) );
  XOR2_X1 U407 ( .A(n374), .B(n427), .Z(n352) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n368) );
  INV_X1 U410 ( .A(KEYINPUT74), .ZN(n353) );
  NAND2_X1 U411 ( .A1(KEYINPUT33), .A2(n353), .ZN(n356) );
  INV_X1 U412 ( .A(KEYINPUT33), .ZN(n354) );
  NAND2_X1 U413 ( .A1(n354), .A2(KEYINPUT74), .ZN(n355) );
  NAND2_X1 U414 ( .A1(n356), .A2(n355), .ZN(n358) );
  XNOR2_X1 U415 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U418 ( .A(KEYINPUT13), .B(KEYINPUT31), .Z(n361) );
  XOR2_X1 U419 ( .A(G176GAT), .B(G120GAT), .Z(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U422 ( .A(n370), .B(n369), .Z(n451) );
  INV_X1 U423 ( .A(n451), .ZN(n415) );
  XOR2_X1 U424 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n411) );
  XOR2_X1 U425 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n372) );
  XNOR2_X1 U426 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U428 ( .A(n373), .B(KEYINPUT11), .Z(n376) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n391) );
  XOR2_X1 U432 ( .A(KEYINPUT64), .B(KEYINPUT78), .Z(n380) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(G85GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U435 ( .A(KEYINPUT76), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U436 ( .A(G99GAT), .B(KEYINPUT75), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U438 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U439 ( .A(G162GAT), .B(G134GAT), .Z(n386) );
  NAND2_X1 U440 ( .A1(G232GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U442 ( .A(G190GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U444 ( .A(n391), .B(n390), .Z(n452) );
  XOR2_X1 U445 ( .A(KEYINPUT36), .B(n452), .Z(n577) );
  XOR2_X1 U446 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n393) );
  XNOR2_X1 U447 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n401) );
  XOR2_X1 U449 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT13), .B(G64GAT), .Z(n395) );
  XNOR2_X1 U451 ( .A(G211GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n409) );
  NAND2_X1 U456 ( .A1(G231GAT), .A2(G233GAT), .ZN(n407) );
  XOR2_X1 U457 ( .A(G78GAT), .B(G155GAT), .Z(n403) );
  XNOR2_X1 U458 ( .A(G15GAT), .B(G127GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U460 ( .A(G183GAT), .B(G71GAT), .Z(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n574) );
  NAND2_X1 U464 ( .A1(n577), .A2(n574), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U466 ( .A1(n415), .A2(n412), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n413), .B(KEYINPUT107), .ZN(n414) );
  NOR2_X1 U468 ( .A1(n552), .A2(n414), .ZN(n422) );
  NAND2_X1 U469 ( .A1(n567), .A2(n557), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n416), .B(KEYINPUT46), .ZN(n417) );
  NAND2_X1 U471 ( .A1(n417), .A2(n452), .ZN(n418) );
  NOR2_X1 U472 ( .A1(n418), .A2(n574), .ZN(n420) );
  INV_X1 U473 ( .A(KEYINPUT47), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  NOR2_X1 U475 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT48), .ZN(n522) );
  NOR2_X1 U477 ( .A1(n424), .A2(n522), .ZN(n425) );
  XOR2_X1 U478 ( .A(n425), .B(KEYINPUT54), .Z(n426) );
  NOR2_X1 U479 ( .A1(n509), .A2(n426), .ZN(n564) );
  XOR2_X1 U480 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U481 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U483 ( .A(KEYINPUT23), .B(G148GAT), .Z(n432) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U486 ( .A(n434), .B(n433), .Z(n439) );
  XOR2_X1 U487 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n436) );
  XNOR2_X1 U488 ( .A(G50GAT), .B(G22GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n437), .B(KEYINPUT88), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n461) );
  NAND2_X1 U493 ( .A1(n564), .A2(n461), .ZN(n445) );
  XOR2_X1 U494 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n443) );
  INV_X1 U495 ( .A(KEYINPUT55), .ZN(n442) );
  NOR2_X1 U496 ( .A1(n524), .A2(n446), .ZN(n560) );
  INV_X1 U497 ( .A(n452), .ZN(n548) );
  NAND2_X1 U498 ( .A1(n560), .A2(n548), .ZN(n450) );
  XOR2_X1 U499 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n448) );
  XNOR2_X1 U500 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n470) );
  NAND2_X1 U502 ( .A1(n552), .A2(n451), .ZN(n483) );
  NAND2_X1 U503 ( .A1(n452), .A2(n574), .ZN(n453) );
  XOR2_X1 U504 ( .A(KEYINPUT16), .B(n453), .Z(n468) );
  XNOR2_X1 U505 ( .A(n511), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U506 ( .A1(n514), .A2(n461), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT26), .B(n454), .Z(n540) );
  INV_X1 U508 ( .A(n540), .ZN(n565) );
  NAND2_X1 U509 ( .A1(n463), .A2(n565), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n514), .A2(n511), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n461), .A2(n455), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT25), .B(n456), .Z(n457) );
  NAND2_X1 U513 ( .A1(n458), .A2(n457), .ZN(n460) );
  NAND2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n467) );
  XOR2_X1 U515 ( .A(n514), .B(KEYINPUT86), .Z(n465) );
  XNOR2_X1 U516 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(n461), .ZN(n527) );
  NAND2_X1 U518 ( .A1(n509), .A2(n463), .ZN(n521) );
  NOR2_X1 U519 ( .A1(n527), .A2(n521), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n480) );
  NAND2_X1 U522 ( .A1(n468), .A2(n480), .ZN(n497) );
  NOR2_X1 U523 ( .A1(n483), .A2(n497), .ZN(n477) );
  NAND2_X1 U524 ( .A1(n477), .A2(n509), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U526 ( .A(G1GAT), .B(n471), .Z(G1324GAT) );
  XOR2_X1 U527 ( .A(G8GAT), .B(KEYINPUT95), .Z(n473) );
  NAND2_X1 U528 ( .A1(n477), .A2(n511), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(G1325GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U531 ( .A1(n477), .A2(n514), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(n476), .ZN(G1326GAT) );
  XOR2_X1 U534 ( .A(G22GAT), .B(KEYINPUT97), .Z(n479) );
  NAND2_X1 U535 ( .A1(n477), .A2(n527), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1327GAT) );
  XOR2_X1 U537 ( .A(G29GAT), .B(KEYINPUT39), .Z(n486) );
  NAND2_X1 U538 ( .A1(n577), .A2(n480), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n574), .A2(n481), .ZN(n482) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(n482), .ZN(n507) );
  NOR2_X1 U541 ( .A1(n507), .A2(n483), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT38), .B(n484), .ZN(n494) );
  NAND2_X1 U543 ( .A1(n509), .A2(n494), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT98), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(G36GAT), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U547 ( .A1(n494), .A2(n511), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1329GAT) );
  XNOR2_X1 U549 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n491) );
  NAND2_X1 U551 ( .A1(n494), .A2(n514), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n494), .A2(n527), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n499) );
  INV_X1 U557 ( .A(n567), .ZN(n496) );
  NAND2_X1 U558 ( .A1(n496), .A2(n557), .ZN(n506) );
  NOR2_X1 U559 ( .A1(n506), .A2(n497), .ZN(n502) );
  NAND2_X1 U560 ( .A1(n509), .A2(n502), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n511), .A2(n502), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U564 ( .A1(n514), .A2(n502), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U567 ( .A1(n502), .A2(n527), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G78GAT), .B(n505), .ZN(G1335GAT) );
  NOR2_X1 U570 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT103), .B(n508), .Z(n517) );
  NAND2_X1 U572 ( .A1(n509), .A2(n517), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n517), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(KEYINPUT104), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  XOR2_X1 U577 ( .A(G99GAT), .B(KEYINPUT105), .Z(n516) );
  NAND2_X1 U578 ( .A1(n517), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n519) );
  NAND2_X1 U581 ( .A1(n517), .A2(n527), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U583 ( .A(G106GAT), .B(n520), .Z(G1339GAT) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT110), .ZN(n529) );
  NOR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT108), .B(n523), .Z(n541) );
  NOR2_X1 U587 ( .A1(n524), .A2(n541), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT109), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n552), .A2(n536), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n531) );
  NAND2_X1 U593 ( .A1(n536), .A2(n557), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n534) );
  NAND2_X1 U597 ( .A1(n536), .A2(n574), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n535), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U601 ( .A1(n536), .A2(n548), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  NOR2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n567), .A2(n549), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  NAND2_X1 U608 ( .A1(n549), .A2(n557), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U611 ( .A1(n574), .A2(n549), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT114), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  XOR2_X1 U614 ( .A(G162GAT), .B(KEYINPUT115), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n560), .A2(n552), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n555) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT118), .B(n556), .Z(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n574), .A2(n560), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n563) );
  XNOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n571) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .Z(n569) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(n566), .Z(n578) );
  NAND2_X1 U633 ( .A1(n578), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n578), .A2(n415), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n578), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

