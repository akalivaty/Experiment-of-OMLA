//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT82), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT67), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT67), .A2(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G128), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT67), .A2(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT67), .A2(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT79), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n201), .B(new_n196), .C1(new_n197), .C2(new_n198), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G110), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n194), .B1(new_n207), .B2(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT24), .B(G110), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT64), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G125), .B(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT80), .A2(G125), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT80), .A2(G125), .ZN(new_n219));
  OAI21_X1  g033(.A(G140), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(G125), .A2(G140), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT16), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT80), .B(G125), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT16), .ZN(new_n226));
  INV_X1    g040(.A(G140), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(G146), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT81), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n224), .A2(KEYINPUT81), .A3(G146), .A4(new_n228), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n211), .A2(new_n217), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n226), .B1(new_n220), .B2(new_n222), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n218), .A2(new_n219), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n236), .A2(KEYINPUT16), .A3(G140), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n229), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n208), .A2(new_n209), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n203), .A2(new_n205), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n239), .B(new_n240), .C1(new_n241), .C2(new_n204), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n233), .A2(KEYINPUT83), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT83), .B1(new_n233), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n191), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT76), .B(G902), .Z(new_n246));
  NAND2_X1  g060(.A1(new_n233), .A2(new_n242), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT83), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n191), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT25), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT77), .B(G217), .Z(new_n254));
  INV_X1    g068(.A(new_n246), .ZN(new_n255));
  INV_X1    g069(.A(G234), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT78), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n245), .A2(new_n259), .A3(new_n251), .A4(new_n246), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n245), .A2(new_n251), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n258), .A2(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n212), .A2(G143), .A3(new_n213), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n267), .A2(KEYINPUT0), .A3(G128), .A4(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT0), .B(G128), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT64), .A2(G146), .ZN(new_n272));
  NOR2_X1   g086(.A1(KEYINPUT64), .A2(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n268), .A2(G146), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI211_X1 g093(.A(KEYINPUT65), .B(new_n271), .C1(new_n274), .C2(new_n276), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n266), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G137), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT11), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n282), .B2(G137), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n284), .A2(new_n290), .A3(new_n286), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n275), .B1(new_n214), .B2(new_n268), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT65), .B1(new_n293), .B2(new_n271), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n277), .A2(new_n278), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT68), .A4(new_n270), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n281), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n192), .A2(G116), .A3(new_n193), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(G116), .B2(new_n207), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT2), .B(G113), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n302), .B(new_n298), .C1(G116), .C2(new_n207), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n267), .A2(G128), .A3(new_n306), .A4(new_n269), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT1), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n196), .B1(new_n267), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n313), .B2(new_n293), .ZN(new_n314));
  INV_X1    g128(.A(new_n287), .ZN(new_n315));
  OAI21_X1  g129(.A(G131), .B1(new_n315), .B2(new_n283), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n291), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n297), .A2(new_n305), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n294), .A2(new_n295), .A3(new_n270), .ZN(new_n323));
  INV_X1    g137(.A(new_n292), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n304), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n329), .A3(new_n320), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(G237), .A2(G953), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G210), .ZN(new_n333));
  XOR2_X1   g147(.A(new_n333), .B(KEYINPUT71), .Z(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G101), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n334), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n305), .B1(new_n325), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT69), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n314), .B2(new_n317), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n297), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n297), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n338), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n319), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT31), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT31), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n346), .A2(new_n350), .A3(new_n319), .A4(new_n347), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n339), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT32), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n338), .B1(new_n327), .B2(KEYINPUT28), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n330), .A3(new_n322), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT73), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n346), .A2(new_n319), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n362), .B2(new_n338), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n319), .A2(new_n329), .A3(new_n320), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n329), .B1(new_n319), .B2(new_n320), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n359), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n319), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n297), .A2(KEYINPUT74), .A3(new_n305), .A4(new_n318), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n297), .A2(new_n318), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n304), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT28), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n338), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n366), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT75), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n376), .A2(new_n366), .A3(new_n381), .A4(new_n378), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n369), .A2(new_n380), .A3(new_n246), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G472), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n265), .B1(new_n358), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G214), .B1(G237), .B2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n298), .B(KEYINPUT5), .C1(G116), .C2(new_n207), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(G113), .C1(KEYINPUT5), .C2(new_n298), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G107), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G101), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT85), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(KEYINPUT3), .C1(new_n390), .C2(G107), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT3), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n392), .A3(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT86), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(new_n401), .A3(new_n392), .A4(G104), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n406), .A3(new_n407), .A4(new_n391), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n389), .A2(new_n395), .A3(new_n408), .A4(new_n303), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n397), .A2(new_n399), .B1(new_n390), .B2(G107), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n407), .B1(new_n411), .B2(new_n406), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  INV_X1    g228(.A(new_n399), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n398), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n391), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n403), .A2(new_n405), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n414), .B(G101), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n304), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n409), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G110), .B(G122), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n422), .B(new_n409), .C1(new_n413), .C2(new_n420), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n427), .A3(new_n423), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n272), .A2(new_n273), .A3(new_n268), .ZN(new_n429));
  OAI21_X1  g243(.A(G128), .B1(new_n429), .B2(new_n306), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n274), .A2(new_n276), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT88), .A3(new_n236), .A4(new_n307), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n236), .B(new_n307), .C1(new_n313), .C2(new_n293), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n323), .A2(new_n225), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G953), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n441), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n426), .A2(new_n428), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n426), .A2(new_n445), .A3(KEYINPUT89), .A4(new_n428), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G210), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n425), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n422), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n409), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n389), .A2(new_n303), .B1(new_n395), .B2(new_n408), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n437), .A2(new_n438), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n437), .B2(new_n438), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n452), .B1(new_n461), .B2(KEYINPUT91), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n457), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n450), .A2(new_n451), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n450), .A2(new_n465), .ZN(new_n467));
  INV_X1    g281(.A(new_n451), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n451), .B1(new_n450), .B2(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT92), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n387), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G113), .B(G122), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(new_n390), .ZN(new_n476));
  INV_X1    g290(.A(G214), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n477), .A2(G237), .A3(G953), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT93), .B1(new_n478), .B2(G143), .ZN(new_n479));
  INV_X1    g293(.A(G237), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n187), .A3(G214), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n268), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n480), .A2(new_n187), .A3(G143), .A4(G214), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT94), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT94), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n332), .A2(new_n486), .A3(G143), .A4(G214), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n479), .A2(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT18), .A2(G131), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n221), .B1(new_n225), .B2(G140), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G146), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n488), .A2(new_n489), .B1(new_n491), .B2(new_n217), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT93), .B(G143), .C1(new_n332), .C2(G214), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n482), .B1(new_n481), .B2(new_n268), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n485), .A2(new_n487), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT18), .B(G131), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n488), .A2(new_n290), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT17), .B(G131), .C1(new_n495), .C2(new_n496), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n238), .A3(new_n229), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n476), .B(new_n498), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(new_n501), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT19), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n216), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(KEYINPUT19), .B2(new_n490), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n215), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n231), .A3(new_n232), .A4(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n476), .B1(new_n512), .B2(new_n498), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT95), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n231), .A2(new_n232), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n499), .A2(new_n501), .B1(new_n510), .B2(new_n215), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n516), .A2(new_n517), .B1(new_n497), .B2(new_n492), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n505), .B(new_n515), .C1(new_n518), .C2(new_n476), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT20), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n505), .B1(new_n518), .B2(new_n476), .ZN(new_n523));
  NOR3_X1   g337(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G952), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n527), .A2(KEYINPUT101), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(KEYINPUT101), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n187), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(G234), .B2(G237), .ZN(new_n531));
  AOI211_X1 g345(.A(new_n187), .B(new_n246), .C1(G234), .C2(G237), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT21), .B(G898), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT9), .B(G234), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n187), .A3(new_n254), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G116), .ZN(new_n540));
  OR2_X1    g354(.A1(KEYINPUT96), .A2(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT96), .A2(G122), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G122), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT97), .B1(new_n544), .B2(G116), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n540), .A3(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n543), .B1(KEYINPUT14), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n392), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n542), .ZN(new_n553));
  NOR2_X1   g367(.A1(KEYINPUT96), .A2(G122), .ZN(new_n554));
  OAI21_X1  g368(.A(G116), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n548), .A3(new_n392), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n196), .A2(G143), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n268), .A2(G128), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G134), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n282), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT100), .B1(new_n552), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n548), .A2(KEYINPUT14), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n551), .A3(new_n555), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G107), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n555), .A2(new_n548), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G107), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n556), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT98), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n575), .A3(new_n556), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  AOI22_X1  g391(.A1(KEYINPUT99), .A2(new_n577), .B1(new_n196), .B2(G143), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(KEYINPUT99), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G134), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n559), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n580), .A2(new_n559), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n574), .A2(new_n576), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n539), .B1(new_n570), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n570), .A2(new_n583), .A3(new_n539), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n255), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G478), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT15), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n587), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(new_n591));
  INV_X1    g405(.A(new_n476), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n593), .B2(new_n505), .ZN(new_n594));
  INV_X1    g408(.A(G475), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n526), .A2(new_n535), .A3(new_n590), .A4(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n594), .A2(new_n595), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n522), .B2(new_n525), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(KEYINPUT102), .A3(new_n535), .A4(new_n590), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G221), .B1(new_n536), .B2(G902), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n408), .A2(new_n395), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n432), .B2(new_n307), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n267), .A2(new_n269), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n196), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n307), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n395), .A3(new_n408), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n607), .A2(new_n609), .B1(new_n613), .B2(new_n608), .ZN(new_n614));
  OAI21_X1  g428(.A(G101), .B1(new_n417), .B2(new_n418), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT4), .A3(new_n408), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n616), .A2(new_n281), .A3(new_n419), .A4(new_n296), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n614), .A2(new_n324), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(G110), .B(G140), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT84), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n187), .A2(G227), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n324), .B1(new_n614), .B2(new_n617), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n614), .A2(new_n617), .A3(new_n324), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n312), .A2(new_n196), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n431), .A2(new_n430), .B1(new_n610), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n606), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n324), .B1(new_n630), .B2(new_n613), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(KEYINPUT87), .A2(KEYINPUT12), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n324), .B(new_n634), .C1(new_n630), .C2(new_n613), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n627), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n624), .A2(new_n626), .B1(new_n636), .B2(new_n623), .ZN(new_n637));
  OAI21_X1  g451(.A(G469), .B1(new_n637), .B2(G902), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n623), .B1(new_n618), .B2(new_n625), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n627), .B(new_n622), .C1(new_n633), .C2(new_n635), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G469), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n246), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n605), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n385), .A2(new_n474), .A3(new_n603), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  OAI211_X1 g460(.A(new_n386), .B(new_n535), .C1(new_n466), .C2(new_n472), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n587), .A2(G478), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n570), .A2(new_n583), .A3(new_n539), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n584), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n649), .B(KEYINPUT33), .C1(new_n650), .C2(new_n584), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n255), .A2(new_n588), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n648), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n647), .A2(new_n601), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(G469), .A2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n636), .A2(new_n623), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n626), .A2(new_n627), .A3(new_n622), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(G469), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n643), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(new_n261), .A3(new_n264), .A4(new_n604), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n352), .A2(new_n353), .ZN(new_n665));
  INV_X1    g479(.A(G472), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n352), .B2(new_n246), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n658), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  NAND2_X1  g485(.A1(new_n585), .A2(new_n586), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n246), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n589), .ZN(new_n674));
  INV_X1    g488(.A(new_n589), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n246), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n596), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n600), .A2(KEYINPUT104), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n521), .B(KEYINPUT20), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n647), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n668), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NOR2_X1   g501(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n247), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n263), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n261), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n644), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n665), .A3(new_n667), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n474), .A2(new_n693), .A3(new_n603), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n532), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n531), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n681), .A2(new_n682), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n358), .B2(new_n384), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n386), .B1(new_n466), .B2(new_n472), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n692), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  NAND3_X1  g520(.A1(new_n450), .A2(new_n451), .A3(new_n465), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n472), .B2(KEYINPUT92), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n470), .B(new_n451), .C1(new_n450), .C2(new_n465), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT38), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n319), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n297), .A2(new_n343), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT69), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n297), .A2(new_n342), .A3(new_n343), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n713), .B1(new_n717), .B2(new_n341), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n338), .ZN(new_n719));
  INV_X1    g533(.A(G902), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n375), .B2(new_n347), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n691), .B1(new_n358), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n601), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n677), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n699), .B(KEYINPUT39), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n644), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n726), .B(new_n386), .C1(KEYINPUT40), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(KEYINPUT40), .B2(new_n728), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n712), .A2(new_n723), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  NAND2_X1  g546(.A1(new_n358), .A2(new_n384), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n601), .A2(new_n657), .A3(new_n699), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n704), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  AOI21_X1  g550(.A(new_n642), .B1(new_n641), .B2(new_n246), .ZN(new_n737));
  AOI211_X1 g551(.A(G469), .B(new_n255), .C1(new_n639), .C2(new_n640), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n605), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n385), .A2(new_n658), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND3_X1  g556(.A1(new_n385), .A2(new_n684), .A3(new_n739), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT105), .B(G116), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G18));
  NAND2_X1  g559(.A1(new_n260), .A2(new_n258), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n747), .A2(new_n253), .B1(new_n263), .B2(new_n689), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n599), .B2(new_n602), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n739), .B(new_n386), .C1(new_n472), .C2(new_n466), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n733), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  NOR2_X1   g567(.A1(new_n703), .A2(new_n725), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n349), .A2(new_n351), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n347), .B1(new_n376), .B2(new_n366), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n353), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n667), .A3(new_n265), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n754), .A2(new_n759), .A3(new_n535), .A4(new_n739), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NOR3_X1   g575(.A1(new_n758), .A2(new_n748), .A3(new_n667), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n751), .A2(new_n762), .A3(new_n734), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  INV_X1    g578(.A(new_n265), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n710), .A2(new_n386), .A3(new_n644), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n377), .B1(new_n718), .B2(new_n347), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n367), .B1(new_n366), .B2(new_n359), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n255), .B1(new_n769), .B2(new_n368), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n380), .A2(new_n382), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n666), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n352), .A2(new_n356), .A3(new_n353), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n356), .B1(new_n352), .B2(new_n353), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n734), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT106), .B1(new_n766), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  INV_X1    g592(.A(new_n734), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n358), .B2(new_n384), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n662), .A2(new_n659), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n604), .B1(new_n781), .B2(new_n738), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n708), .A2(new_n709), .A3(new_n387), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n783), .A3(new_n784), .A4(new_n765), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n777), .A2(new_n778), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n783), .A3(KEYINPUT42), .A4(new_n765), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(KEYINPUT107), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n777), .A2(new_n790), .A3(new_n778), .A4(new_n785), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  NAND3_X1  g607(.A1(new_n702), .A2(new_n783), .A3(new_n765), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  OR2_X1    g609(.A1(new_n637), .A2(KEYINPUT45), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n637), .A2(KEYINPUT45), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(G469), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT46), .B1(new_n798), .B2(new_n659), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n738), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n659), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n605), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n727), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT108), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n708), .A2(new_n387), .A3(new_n709), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n657), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n601), .ZN(new_n808));
  NAND2_X1  g622(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n691), .C1(new_n665), .C2(new_n667), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n806), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n802), .B1(KEYINPUT110), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n802), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n355), .A2(new_n357), .B1(new_n383), .B2(G472), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n805), .A2(new_n823), .A3(new_n265), .A4(new_n734), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G140), .ZN(G42));
  NOR2_X1   g640(.A1(new_n737), .A2(new_n738), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT49), .Z(new_n828));
  NAND2_X1  g642(.A1(new_n604), .A2(new_n386), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n828), .A2(new_n265), .A3(new_n808), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n722), .B1(new_n773), .B2(new_n774), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n711), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n812), .A2(new_n531), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n759), .ZN(new_n836));
  INV_X1    g650(.A(new_n739), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n836), .A2(new_n712), .A3(new_n386), .A4(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT50), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n832), .A2(new_n531), .A3(new_n765), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n806), .A2(new_n837), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n601), .A2(new_n841), .A3(new_n657), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n834), .A2(new_n837), .A3(new_n806), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n762), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n836), .A2(new_n806), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n827), .A2(new_n605), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n822), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(KEYINPUT51), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT114), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n645), .A2(new_n740), .A3(new_n743), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n469), .A2(new_n470), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n473), .A3(new_n707), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n521), .A2(KEYINPUT20), .B1(new_n523), .B2(new_n524), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n657), .B1(new_n600), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n601), .A2(new_n590), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n857), .A2(new_n858), .A3(new_n535), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n668), .A2(new_n855), .A3(new_n859), .A4(new_n386), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n694), .A2(new_n752), .A3(new_n760), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n677), .A2(new_n699), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n682), .A3(new_n679), .A4(new_n680), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n692), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n733), .A2(new_n805), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n701), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n772), .B2(new_n775), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n766), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n667), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n870), .A2(new_n734), .A3(new_n691), .A4(new_n757), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n783), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n783), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT111), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n869), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n789), .A2(new_n791), .A3(new_n862), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n663), .A2(new_n604), .A3(new_n700), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n754), .A2(new_n748), .A3(new_n831), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n705), .A2(new_n735), .A3(new_n880), .A4(new_n763), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT113), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n703), .A2(new_n725), .A3(new_n878), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n704), .A2(new_n780), .B1(new_n723), .B2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n704), .A2(new_n702), .B1(new_n871), .B2(new_n751), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n882), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n469), .A2(new_n707), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n386), .A3(new_n644), .A4(new_n691), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n823), .A2(new_n892), .A3(new_n701), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n870), .A2(new_n734), .A3(new_n691), .A4(new_n757), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n750), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n890), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n705), .A2(KEYINPUT112), .A3(new_n763), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n735), .A3(new_n880), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT52), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n889), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n881), .A2(KEYINPUT113), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n886), .B1(new_n884), .B2(new_n885), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT52), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n889), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n789), .A2(new_n791), .A3(new_n862), .A4(new_n876), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n899), .A2(new_n889), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n901), .B1(new_n910), .B2(new_n906), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n882), .A2(new_n888), .A3(new_n887), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n888), .B1(new_n882), .B2(new_n887), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n877), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(new_n901), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n909), .B1(new_n916), .B2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n844), .A2(new_n385), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT48), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(KEYINPUT116), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n836), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n530), .B1(new_n921), .B2(new_n751), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n841), .A2(new_n842), .A3(new_n724), .A4(new_n807), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n845), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n847), .A3(new_n929), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n920), .B(new_n926), .C1(new_n927), .C2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n852), .A2(new_n917), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(G952), .A2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n833), .B1(new_n932), .B2(new_n933), .ZN(G75));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n914), .B2(new_n877), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n910), .A2(new_n906), .A3(new_n901), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n937), .A2(new_n451), .A3(new_n246), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n426), .A2(new_n428), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT117), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n445), .B(KEYINPUT55), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n187), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n939), .A2(new_n943), .ZN(new_n948));
  OR3_X1    g762(.A1(new_n947), .A2(KEYINPUT118), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT118), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G51));
  XOR2_X1   g765(.A(new_n659), .B(KEYINPUT57), .Z(new_n952));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT54), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n937), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT54), .B1(new_n935), .B2(new_n936), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n900), .A2(new_n907), .A3(new_n953), .A4(new_n954), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n952), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n960), .A3(new_n641), .ZN(new_n961));
  OR3_X1    g775(.A1(new_n937), .A2(new_n246), .A3(new_n798), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n959), .B2(new_n641), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n946), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT121), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n967), .B(new_n946), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G54));
  NAND4_X1  g783(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .A4(new_n255), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n514), .A2(new_n519), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n972), .A2(new_n973), .A3(new_n945), .ZN(G60));
  INV_X1    g788(.A(new_n655), .ZN(new_n975));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT59), .Z(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n917), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n955), .A2(new_n958), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n982), .A2(new_n975), .A3(new_n977), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n980), .A2(new_n981), .A3(new_n945), .A4(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT123), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n908), .A2(new_n689), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT124), .Z(new_n989));
  AOI21_X1  g803(.A(new_n262), .B1(new_n908), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n945), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g807(.A(G953), .B1(new_n533), .B2(new_n440), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n862), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n941), .B1(G898), .B2(new_n187), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G69));
  NAND2_X1  g811(.A1(new_n325), .A2(new_n340), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n717), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n510), .Z(new_n1000));
  AND3_X1   g814(.A1(new_n896), .A2(new_n735), .A3(new_n897), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n731), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  INV_X1    g817(.A(new_n385), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n857), .A2(new_n858), .ZN(new_n1005));
  OR4_X1    g819(.A1(new_n1004), .A2(new_n806), .A3(new_n728), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n825), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1003), .A2(new_n1007), .A3(new_n817), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1000), .B1(new_n1009), .B2(new_n187), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT125), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G900), .A2(G953), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n825), .A2(new_n794), .ZN(new_n1015));
  INV_X1    g829(.A(new_n804), .ZN(new_n1016));
  INV_X1    g830(.A(new_n754), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n816), .B1(new_n1004), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n792), .A3(new_n1001), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1000), .B(new_n1014), .C1(new_n1020), .C2(G953), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1012), .A2(new_n1013), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(G72));
  XNOR2_X1  g838(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n666), .A2(new_n720), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n862), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n362), .A2(new_n347), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n945), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n719), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1030), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n916), .A2(new_n1032), .A3(new_n1033), .A4(new_n1027), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1027), .B1(new_n1009), .B2(new_n1028), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n719), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1031), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(KEYINPUT127), .ZN(G57));
endmodule


