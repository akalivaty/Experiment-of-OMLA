//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n207), .A2(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT85), .B2(new_n207), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT86), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n211), .B2(new_n210), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n205), .A2(KEYINPUT87), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(new_n204), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT86), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n210), .B2(new_n211), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n214), .A2(new_n218), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n213), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT17), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT97), .B(G92gat), .Z(new_n229));
  INV_X1    g028(.A(G85gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT7), .ZN(new_n233));
  INV_X1    g032(.A(G99gat), .ZN(new_n234));
  INV_X1    g033(.A(G106gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT8), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G99gat), .B(G106gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT98), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n228), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G190gat), .B(G218gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT99), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n239), .A2(KEYINPUT98), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n239), .A2(KEYINPUT98), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n227), .ZN(new_n246));
  AND2_X1   g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT41), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n241), .A2(new_n243), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT100), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n246), .A2(new_n248), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(KEYINPUT100), .A3(new_n243), .A4(new_n241), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT101), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n251), .B2(new_n253), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n243), .B1(new_n252), .B2(new_n241), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n247), .A2(KEYINPUT41), .ZN(new_n260));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT102), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT102), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n257), .A2(new_n258), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n265), .B(new_n262), .C1(new_n266), .C2(new_n256), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n258), .A2(new_n262), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n253), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT103), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G155gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT20), .Z(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G64gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT91), .ZN(new_n277));
  NAND2_X1  g076(.A1(G71gat), .A2(G78gat), .ZN(new_n278));
  INV_X1    g077(.A(G71gat), .ZN(new_n279));
  INV_X1    g078(.A(G78gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT9), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT92), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n278), .B(new_n281), .C1(new_n276), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288));
  INV_X1    g087(.A(G231gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n287), .B2(new_n288), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n275), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OR3_X1    g095(.A1(new_n294), .A2(new_n275), .A3(new_n295), .ZN(new_n297));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT16), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(G1gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G1gat), .B2(new_n298), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(G8gat), .Z(new_n302));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT94), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT94), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n304), .A3(new_n286), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(new_n288), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n307), .A2(new_n309), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n296), .B(new_n297), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n296), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n320), .A3(new_n316), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT104), .ZN(new_n326));
  XNOR2_X1  g125(.A(G120gat), .B(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G230gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(new_n290), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT10), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n240), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n303), .A3(new_n305), .ZN(new_n335));
  INV_X1    g134(.A(new_n239), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n287), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n285), .A2(new_n286), .A3(new_n239), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n332), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n332), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n337), .B2(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n330), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n340), .A2(new_n342), .A3(new_n330), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n326), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT104), .A3(new_n343), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G113gat), .B(G141gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(G197gat), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT11), .B(G169gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n353), .B(KEYINPUT12), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n228), .A2(new_n302), .ZN(new_n356));
  NAND2_X1  g155(.A1(G229gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n227), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(new_n302), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT18), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n358), .B(new_n302), .ZN(new_n363));
  XOR2_X1   g162(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(new_n357), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n356), .A2(new_n359), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT18), .A3(new_n357), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n355), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(new_n355), .A3(new_n366), .A4(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT90), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n372), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR4_X1   g174(.A1(new_n273), .A2(new_n325), .A3(new_n349), .A4(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(KEYINPUT24), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382));
  INV_X1    g181(.A(G169gat), .ZN(new_n383));
  INV_X1    g182(.A(G176gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G183gat), .ZN(new_n387));
  INV_X1    g186(.A(G190gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(KEYINPUT24), .A3(new_n379), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n380), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(new_n381), .ZN(new_n393));
  AND4_X1   g192(.A1(KEYINPUT25), .A2(new_n392), .A3(new_n393), .A4(new_n390), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n383), .A2(new_n384), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(KEYINPUT65), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT65), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n396), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n379), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT27), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G183gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n388), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n387), .A2(KEYINPUT27), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n408), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  AND4_X1   g215(.A1(KEYINPUT28), .A2(new_n410), .A3(new_n414), .A4(new_n388), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n406), .A2(new_n407), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n405), .A2(KEYINPUT66), .A3(new_n379), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n395), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT70), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT71), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n377), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n421), .B2(KEYINPUT29), .ZN(new_n427));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G211gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT69), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G211gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT22), .B1(new_n434), .B2(G218gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(G197gat), .B(G204gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n429), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G218gat), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n431), .B2(new_n433), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n436), .B(new_n428), .C1(new_n440), .C2(KEYINPUT22), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n406), .A2(new_n407), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n416), .A2(new_n418), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n420), .A3(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n391), .A2(new_n394), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT72), .A3(new_n424), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n426), .A2(new_n427), .A3(new_n442), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n405), .A2(KEYINPUT66), .A3(new_n379), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT66), .B1(new_n405), .B2(new_n379), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT27), .B(G183gat), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n388), .B(new_n412), .C1(new_n455), .C2(new_n411), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n417), .B1(new_n456), .B2(new_n408), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n452), .B1(new_n458), .B2(new_n395), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n425), .B1(new_n445), .B2(new_n446), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n459), .A2(new_n423), .B1(new_n460), .B2(KEYINPUT72), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(KEYINPUT73), .A3(new_n442), .A4(new_n426), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n424), .B1(new_n447), .B2(new_n452), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n421), .A2(new_n423), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n442), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT37), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n451), .A2(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n426), .A2(new_n427), .A3(new_n467), .A4(new_n448), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n442), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT37), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT83), .A4(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n474), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n467), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n489), .A3(new_n472), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT0), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT75), .ZN(new_n496));
  AND2_X1   g295(.A1(G141gat), .A2(G148gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(G141gat), .A2(G148gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G141gat), .ZN(new_n500));
  INV_X1    g299(.A(G148gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G141gat), .A2(G148gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT75), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT2), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G155gat), .ZN(new_n507));
  INV_X1    g306(.A(G162gat), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT74), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT74), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G155gat), .B(G162gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n498), .ZN(new_n515));
  OR2_X1    g314(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n507), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n514), .B(new_n515), .C1(new_n518), .C2(new_n505), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G127gat), .B(G134gat), .Z(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G120gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(KEYINPUT1), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G113gat), .B(G120gat), .Z(new_n524));
  INV_X1    g323(.A(KEYINPUT1), .ZN(new_n525));
  XNOR2_X1  g324(.A(G127gat), .B(G134gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n519), .A3(new_n527), .A4(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT5), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n523), .A2(new_n527), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n520), .B2(KEYINPUT3), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT3), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n513), .A2(new_n538), .A3(new_n519), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n520), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n541), .A2(KEYINPUT77), .A3(new_n542), .A4(new_n536), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n536), .A2(new_n542), .A3(new_n519), .A4(new_n513), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n530), .A2(KEYINPUT4), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n535), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT78), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n550), .A3(new_n544), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT5), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n541), .A2(KEYINPUT78), .A3(new_n542), .A4(new_n536), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n540), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(KEYINPUT6), .B(new_n495), .C1(new_n549), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n495), .B1(new_n549), .B2(new_n555), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n548), .A2(new_n540), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n494), .B(new_n554), .C1(new_n558), .C2(new_n535), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n490), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n472), .B1(new_n463), .B2(new_n468), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n486), .A2(new_n485), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n563), .A2(KEYINPUT84), .A3(new_n484), .A4(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n478), .A2(new_n488), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n490), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n473), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n475), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n463), .A2(new_n489), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n473), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n537), .A2(new_n539), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n574), .A3(new_n553), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT39), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(new_n533), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n575), .A2(new_n533), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n529), .A2(new_n532), .A3(new_n530), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT39), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT81), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT81), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n582), .A3(KEYINPUT39), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n494), .B(new_n577), .C1(new_n578), .C2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n557), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT82), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G228gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n290), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n441), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT22), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT69), .B(G211gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n439), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n428), .B1(new_n599), .B2(new_n436), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n452), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n541), .B1(new_n601), .B2(new_n538), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n442), .B1(new_n452), .B2(new_n539), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n595), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G22gat), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT29), .B1(new_n438), .B2(new_n441), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n520), .B1(new_n606), .B2(KEYINPUT3), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n539), .A2(new_n452), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n467), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n609), .A3(new_n594), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT79), .ZN(new_n612));
  XNOR2_X1  g411(.A(G78gat), .B(G106gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT31), .B(G50gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT80), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n605), .B1(new_n604), .B2(new_n610), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT80), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n621), .A3(new_n615), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n612), .B2(new_n615), .ZN(new_n624));
  INV_X1    g423(.A(new_n615), .ZN(new_n625));
  AOI211_X1 g424(.A(KEYINPUT80), .B(new_n625), .C1(new_n611), .C2(KEYINPUT79), .ZN(new_n626));
  OAI22_X1  g425(.A1(new_n624), .A2(new_n626), .B1(new_n618), .B2(new_n619), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n573), .A2(new_n592), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n447), .A2(new_n528), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n421), .A2(new_n536), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G227gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n633), .ZN(new_n636));
  INV_X1    g435(.A(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G15gat), .B(G43gat), .Z(new_n639));
  XNOR2_X1  g438(.A(G71gat), .B(G99gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n633), .B1(new_n629), .B2(new_n630), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(KEYINPUT33), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT32), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n645), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n635), .B(new_n638), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n638), .A2(new_n635), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n645), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(KEYINPUT68), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n649), .B2(new_n651), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT68), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n649), .A2(new_n651), .A3(new_n650), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n655), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT36), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n566), .A2(new_n628), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n561), .A2(new_n556), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n568), .A2(new_n663), .A3(new_n572), .A4(new_n570), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n623), .A2(new_n627), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n623), .A2(new_n627), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT35), .B1(new_n668), .B2(new_n664), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n665), .A2(KEYINPUT35), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n657), .ZN(new_n671));
  INV_X1    g470(.A(new_n573), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n663), .A4(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n662), .A2(new_n666), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n376), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n376), .A2(KEYINPUT105), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n663), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g482(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G8gat), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n684), .B2(new_n687), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT108), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n689), .A2(new_n693), .A3(new_n697), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1325gat));
  INV_X1    g498(.A(G15gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n680), .A2(new_n700), .A3(new_n671), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n658), .A2(new_n661), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n678), .B2(new_n679), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n703), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g503(.A1(new_n680), .A2(new_n665), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NOR3_X1   g507(.A1(new_n349), .A2(new_n375), .A3(new_n324), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n566), .A2(new_n628), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n666), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT110), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n710), .A2(new_n702), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n673), .A2(new_n669), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n273), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n268), .A2(new_n272), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n674), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n709), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n663), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n675), .A2(new_n273), .A3(new_n709), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n203), .A3(new_n681), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1328gat));
  OAI21_X1  g532(.A(G36gat), .B1(new_n728), .B2(new_n672), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n730), .A2(new_n204), .A3(new_n573), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT46), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1329gat));
  OAI21_X1  g536(.A(G43gat), .B1(new_n725), .B2(new_n702), .ZN(new_n738));
  INV_X1    g537(.A(G43gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n730), .A2(new_n739), .A3(new_n671), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(KEYINPUT47), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  INV_X1    g541(.A(new_n702), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n743), .A3(new_n727), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n744), .B2(G43gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n745), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g545(.A(G50gat), .B1(new_n725), .B2(new_n667), .ZN(new_n747));
  INV_X1    g546(.A(G50gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n748), .A3(new_n665), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(KEYINPUT48), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n749), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n665), .A3(new_n727), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(G50gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n753), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n717), .A2(new_n718), .ZN(new_n755));
  INV_X1    g554(.A(new_n349), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n370), .A2(new_n372), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n370), .A2(new_n372), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n273), .A2(new_n756), .A3(new_n325), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n681), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n672), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n761), .B2(new_n702), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n671), .A2(new_n279), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g572(.A1(new_n761), .A2(new_n667), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n280), .ZN(G1335gat));
  OAI211_X1 g574(.A(new_n322), .B(new_n323), .C1(new_n757), .C2(new_n758), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n349), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n721), .B2(new_n724), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n714), .A2(new_n716), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT111), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT110), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n664), .B2(new_n665), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n662), .A2(new_n786), .B1(new_n669), .B2(new_n673), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n715), .ZN(new_n788));
  INV_X1    g587(.A(new_n720), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n783), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n778), .B1(new_n790), .B2(new_n723), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n781), .A2(new_n681), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n230), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n776), .B1(new_n268), .B2(new_n272), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n798), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n800), .B(new_n803), .Z(new_n804));
  NAND3_X1  g603(.A1(new_n349), .A2(new_n230), .A3(new_n681), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n797), .B1(new_n804), .B2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(new_n229), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n780), .B2(new_n672), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n756), .A2(G92gat), .A3(new_n672), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n808), .B(new_n809), .C1(new_n804), .C2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n273), .A2(new_n777), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT116), .B1(new_n787), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n782), .A2(new_n816), .A3(new_n798), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT117), .A4(new_n802), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n799), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n817), .A3(new_n802), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n811), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n791), .A2(new_n792), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT113), .B(new_n778), .C1(new_n790), .C2(new_n723), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n825), .A2(new_n826), .A3(new_n672), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n229), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n813), .B1(new_n828), .B2(KEYINPUT52), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n781), .A2(new_n573), .A3(new_n793), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n823), .B1(new_n830), .B2(new_n807), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n809), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n812), .B1(new_n829), .B2(new_n832), .ZN(G1337gat));
  NOR3_X1   g632(.A1(new_n825), .A2(new_n826), .A3(new_n702), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n349), .A2(new_n234), .A3(new_n671), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n834), .A2(new_n234), .B1(new_n804), .B2(new_n835), .ZN(G1338gat));
  OAI21_X1  g635(.A(G106gat), .B1(new_n780), .B2(new_n667), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n756), .A2(G106gat), .A3(new_n667), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n837), .B(new_n838), .C1(new_n804), .C2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n819), .B2(new_n822), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n781), .A2(new_n665), .A3(new_n793), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(G106gat), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n844), .B2(new_n838), .ZN(G1339gat));
  INV_X1    g644(.A(new_n340), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n335), .A2(new_n332), .A3(new_n339), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n329), .B1(new_n340), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n347), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n850), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(new_n374), .A3(new_n373), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n368), .A2(new_n357), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n363), .A2(new_n365), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n353), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n371), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n346), .A2(new_n348), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n346), .A2(new_n348), .A3(KEYINPUT119), .A4(new_n860), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n722), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n273), .A2(new_n855), .A3(new_n852), .A4(new_n860), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n325), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n273), .A2(new_n325), .A3(new_n349), .A4(new_n759), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n681), .A3(new_n667), .A4(new_n660), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n573), .ZN(new_n874));
  AOI21_X1  g673(.A(G113gat), .B1(new_n874), .B2(new_n759), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n324), .B1(new_n866), .B2(new_n867), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n667), .B(new_n671), .C1(new_n876), .C2(new_n870), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n573), .A2(new_n663), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n759), .A2(G113gat), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n880), .B2(new_n349), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT120), .Z(new_n885));
  NAND3_X1  g684(.A1(new_n874), .A2(new_n883), .A3(new_n349), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1341gat));
  INV_X1    g686(.A(G127gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n874), .A2(new_n888), .A3(new_n324), .ZN(new_n889));
  INV_X1    g688(.A(new_n880), .ZN(new_n890));
  OAI21_X1  g689(.A(G127gat), .B1(new_n890), .B2(new_n325), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1342gat));
  OR3_X1    g691(.A1(new_n722), .A2(G134gat), .A3(new_n573), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT56), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT121), .Z(new_n895));
  NOR3_X1   g694(.A1(new_n873), .A2(KEYINPUT56), .A3(new_n893), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n273), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(G134gat), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1343gat));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n665), .B1(new_n876), .B2(new_n870), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n373), .A2(new_n347), .A3(new_n374), .A4(new_n851), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n848), .A2(new_n903), .A3(new_n850), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n848), .B2(new_n850), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT55), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n861), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n722), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n867), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n325), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n871), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n667), .A2(new_n900), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n900), .A2(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n743), .A2(new_n879), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT123), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n872), .B2(new_n665), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n900), .B(new_n667), .C1(new_n910), .C2(new_n871), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n917), .B(new_n914), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n920), .A3(new_n759), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n876), .A2(new_n870), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n663), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n743), .A2(new_n573), .A3(new_n667), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n375), .A2(G141gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n927), .A2(new_n928), .B1(KEYINPUT124), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(KEYINPUT124), .A3(new_n928), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n913), .A2(new_n375), .A3(new_n915), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n500), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n922), .A2(new_n930), .B1(new_n929), .B2(new_n933), .ZN(G1344gat));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n920), .A3(new_n349), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n501), .A2(KEYINPUT59), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n914), .A2(new_n349), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n665), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n900), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n872), .A2(new_n912), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT59), .B1(new_n942), .B2(new_n501), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n926), .A2(G148gat), .A3(new_n756), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1345gat));
  NAND3_X1  g746(.A1(new_n927), .A2(new_n507), .A3(new_n324), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n916), .A2(new_n920), .A3(new_n324), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n507), .ZN(G1346gat));
  AND3_X1   g749(.A1(new_n916), .A2(new_n920), .A3(new_n273), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n516), .A2(new_n517), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n273), .A2(new_n952), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n951), .A2(new_n952), .B1(new_n926), .B2(new_n953), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n672), .A2(new_n681), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n877), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n958), .A2(new_n383), .A3(new_n375), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n668), .A2(new_n672), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n923), .A2(new_n681), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n872), .A2(KEYINPUT126), .A3(new_n663), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n759), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n959), .B1(new_n966), .B2(new_n383), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n965), .B2(new_n349), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n923), .A2(new_n665), .ZN(new_n969));
  AND4_X1   g768(.A1(G176gat), .A2(new_n349), .A3(new_n671), .A4(new_n955), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(G1349gat));
  NAND2_X1  g770(.A1(new_n324), .A2(new_n455), .ZN(new_n972));
  AOI211_X1 g771(.A(new_n961), .B(new_n972), .C1(new_n963), .C2(new_n964), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n387), .B1(new_n957), .B2(new_n324), .ZN(new_n974));
  OAI21_X1  g773(.A(KEYINPUT60), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  INV_X1    g775(.A(new_n974), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT126), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n960), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n976), .B(new_n977), .C1(new_n979), .C2(new_n972), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n975), .A2(new_n980), .ZN(G1350gat));
  NOR2_X1   g780(.A1(new_n722), .A2(G190gat), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n983));
  INV_X1    g782(.A(new_n964), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n960), .B(new_n982), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n957), .A2(new_n273), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(G190gat), .ZN(new_n988));
  AOI211_X1 g787(.A(KEYINPUT61), .B(new_n388), .C1(new_n957), .C2(new_n273), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n992), .B(new_n985), .C1(new_n988), .C2(new_n989), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1351gat));
  NOR2_X1   g793(.A1(new_n743), .A2(new_n956), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n996), .B1(new_n940), .B2(new_n941), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(G197gat), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n998), .A2(new_n999), .A3(new_n375), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n743), .A2(new_n672), .A3(new_n667), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n978), .A2(new_n759), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1000), .B1(new_n1002), .B2(new_n999), .ZN(G1352gat));
  NAND2_X1  g802(.A1(new_n978), .A2(new_n1001), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n756), .A2(G204gat), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n978), .A2(new_n1008), .A3(new_n1001), .A4(new_n1005), .ZN(new_n1009));
  OAI21_X1  g808(.A(G204gat), .B1(new_n998), .B2(new_n756), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(G1353gat));
  NAND2_X1  g810(.A1(new_n997), .A2(new_n324), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1012), .B2(G211gat), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT63), .ZN(new_n1014));
  AOI211_X1 g813(.A(new_n1014), .B(new_n430), .C1(new_n997), .C2(new_n324), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n324), .A2(new_n598), .ZN(new_n1016));
  OAI22_X1  g815(.A1(new_n1013), .A2(new_n1015), .B1(new_n1004), .B2(new_n1016), .ZN(G1354gat));
  OAI21_X1  g816(.A(G218gat), .B1(new_n998), .B2(new_n722), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n273), .A2(new_n439), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1018), .B1(new_n1004), .B2(new_n1019), .ZN(G1355gat));
endmodule


