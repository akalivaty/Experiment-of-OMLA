//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(KEYINPUT82), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  OAI211_X1 g0045(.A(G1), .B(G13), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G41), .A2(G45), .ZN(new_n251));
  OAI211_X1 g0051(.A(G238), .B(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n251), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(new_n206), .A3(G274), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G232), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n246), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT13), .B1(new_n255), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT13), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(new_n254), .A4(new_n252), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT78), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(KEYINPUT78), .B(KEYINPUT13), .C1(new_n255), .C2(new_n265), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G179), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT81), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(new_n271), .A3(KEYINPUT77), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(new_n255), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT77), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(new_n269), .A4(new_n270), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT80), .A2(G169), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n278), .A2(new_n279), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT81), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n275), .A2(new_n287), .A3(G179), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n277), .A2(new_n284), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n213), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n293), .A3(new_n213), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n207), .A2(new_n244), .A3(KEYINPUT71), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G20), .B2(G33), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n202), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n207), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G77), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n300), .A2(new_n301), .B1(new_n207), .B2(G68), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT66), .B(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n291), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(G68), .A3(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n308), .B(KEYINPUT79), .Z(new_n309));
  NAND4_X1  g0109(.A1(new_n247), .A2(new_n249), .A3(G13), .A4(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n304), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n289), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n275), .A2(G190), .ZN(new_n318));
  INV_X1    g0118(.A(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n278), .A2(G200), .A3(new_n282), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n243), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n296), .A2(new_n298), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT70), .ZN(new_n328));
  INV_X1    g0128(.A(G58), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n329), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n326), .B1(new_n331), .B2(new_n300), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n295), .B1(new_n202), .B2(new_n311), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n295), .B1(G20), .B2(new_n305), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G50), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT9), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n333), .A2(KEYINPUT9), .A3(new_n335), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n244), .ZN(new_n339));
  NAND2_X1  g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(G222), .A3(new_n257), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT67), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n261), .A2(new_n262), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n257), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT68), .B(G223), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n346), .A2(new_n347), .B1(G77), .B2(new_n345), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n246), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n268), .B1(new_n305), .B2(new_n253), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G226), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n254), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n336), .B(new_n337), .C1(G190), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n353), .A2(KEYINPUT76), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT76), .B1(new_n353), .B2(new_n355), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n324), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n358), .A3(new_n324), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n333), .A2(new_n335), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n353), .B2(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT72), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT72), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n366), .B(new_n363), .C1(new_n353), .C2(G169), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n353), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n306), .A2(G77), .A3(new_n307), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G77), .B2(new_n310), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n327), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n325), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n377), .B1(new_n207), .B2(new_n301), .C1(new_n300), .C2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n374), .B1(new_n379), .B2(new_n291), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n346), .A2(G238), .ZN(new_n382));
  AOI21_X1  g0182(.A(G1698), .B1(new_n339), .B2(new_n340), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(G232), .B1(new_n345), .B2(G107), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n246), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n350), .A2(G244), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n254), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n368), .ZN(new_n389));
  INV_X1    g0189(.A(G169), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n385), .B2(new_n387), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n381), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(KEYINPUT74), .A3(G190), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n380), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n388), .A2(G190), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT74), .B1(new_n388), .B2(new_n355), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n323), .A2(new_n362), .A3(new_n372), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n339), .A2(new_n207), .A3(new_n340), .ZN(new_n403));
  AND2_X1   g0203(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n404));
  NOR2_X1   g0204(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n340), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n312), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n325), .A2(G159), .ZN(new_n410));
  XNOR2_X1  g0210(.A(G58), .B(G68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G20), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n402), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n325), .A2(G159), .B1(new_n411), .B2(G20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G68), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n403), .A2(new_n405), .A3(new_n404), .ZN(new_n418));
  OAI211_X1 g0218(.A(KEYINPUT16), .B(new_n415), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n291), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT84), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n414), .A2(new_n419), .A3(KEYINPUT84), .A4(new_n291), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n331), .A2(new_n310), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n334), .B2(new_n331), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n350), .A2(G232), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n256), .A2(G1698), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n430), .B1(G223), .B2(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n246), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n433), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(G179), .A3(new_n428), .A4(new_n254), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n401), .B1(new_n427), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n426), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n422), .B2(new_n423), .ZN(new_n440));
  INV_X1    g0240(.A(new_n437), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT85), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n427), .A2(new_n401), .A3(new_n437), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT85), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n440), .B2(new_n441), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n435), .A2(new_n254), .A3(new_n428), .ZN(new_n448));
  INV_X1    g0248(.A(G190), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(G200), .B2(new_n448), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(KEYINPUT17), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT17), .B1(new_n440), .B2(new_n451), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n443), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n317), .A2(new_n243), .A3(new_n322), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n400), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n341), .A2(G244), .A3(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G116), .ZN(new_n460));
  OAI211_X1 g0260(.A(G238), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n268), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  AOI21_X1  g0264(.A(G274), .B1(KEYINPUT90), .B2(G250), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n250), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT90), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G250), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n305), .B2(G45), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n246), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n390), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(G179), .B2(new_n471), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n247), .A2(new_n249), .A3(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n292), .A2(new_n310), .A3(new_n294), .A4(new_n474), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n475), .A2(KEYINPUT93), .A3(new_n378), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT93), .B1(new_n475), .B2(new_n378), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT92), .ZN(new_n479));
  INV_X1    g0279(.A(new_n378), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(new_n310), .ZN(new_n481));
  NAND3_X1  g0281(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n207), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  INV_X1    g0284(.A(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n207), .A2(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT91), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n207), .B(G68), .C1(new_n261), .C2(new_n262), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT19), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n300), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n489), .A2(new_n491), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  AOI211_X1 g0296(.A(new_n479), .B(new_n481), .C1(new_n496), .C2(new_n291), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n492), .B(new_n495), .C1(new_n490), .C2(KEYINPUT91), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n487), .A2(new_n488), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n291), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n481), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT92), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n478), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT94), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(KEYINPUT94), .B(new_n478), .C1(new_n497), .C2(new_n502), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n473), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n407), .A2(new_n408), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G107), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n325), .A2(G77), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n511));
  XNOR2_X1  g0311(.A(G97), .B(G107), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT87), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  MUX2_X1   g0314(.A(new_n513), .B(G97), .S(KEYINPUT6), .Z(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(G20), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n509), .A2(new_n511), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n291), .ZN(new_n519));
  OR3_X1    g0319(.A1(new_n310), .A2(KEYINPUT88), .A3(G97), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT88), .B1(new_n310), .B2(G97), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n494), .C2(new_n475), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT4), .B1(new_n383), .B2(G244), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n268), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G41), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n247), .A2(new_n249), .A3(new_n533), .A4(G45), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n532), .A2(G41), .ZN(new_n535));
  OAI211_X1 g0335(.A(G257), .B(new_n246), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n305), .A2(KEYINPUT89), .A3(G45), .A4(new_n533), .ZN(new_n539));
  OAI21_X1  g0339(.A(G274), .B1(new_n532), .B2(G41), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n268), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n531), .A2(new_n368), .A3(new_n536), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n531), .A2(new_n536), .A3(new_n542), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n390), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n524), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n522), .B1(new_n518), .B2(new_n291), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(G200), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n449), .C2(new_n544), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n497), .A2(new_n502), .B1(new_n485), .B2(new_n475), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n471), .A2(G200), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n449), .B2(new_n471), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n507), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT23), .ZN(new_n557));
  INV_X1    g0357(.A(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT96), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(KEYINPUT96), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n207), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n341), .A2(new_n568), .A3(new_n207), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n565), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n291), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(new_n576), .C1(new_n244), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n268), .ZN(new_n579));
  OAI211_X1 g0379(.A(G264), .B(new_n246), .C1(new_n534), .C2(new_n535), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n579), .A2(G190), .A3(new_n542), .A4(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n475), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n311), .A2(KEYINPUT25), .A3(new_n558), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT25), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n310), .B2(G107), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n582), .A2(G107), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n542), .A3(new_n580), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n574), .A2(new_n581), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G270), .B(new_n246), .C1(new_n534), .C2(new_n535), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n542), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n592));
  OAI211_X1 g0392(.A(G257), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n339), .A2(G303), .A3(new_n340), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT95), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT95), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n592), .A2(new_n593), .A3(new_n597), .A4(new_n594), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n268), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n591), .A2(G190), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n311), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n310), .A2(new_n307), .A3(new_n474), .A4(G116), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n526), .B(new_n207), .C1(G33), .C2(new_n494), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(G20), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n291), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n542), .A2(new_n590), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n246), .B1(new_n595), .B2(KEYINPUT95), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n598), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n600), .B(new_n611), .C1(new_n614), .C2(new_n355), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n589), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n607), .B(KEYINPUT20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n602), .A2(new_n603), .ZN(new_n619));
  OAI21_X1  g0419(.A(G169), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n591), .A2(new_n599), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(KEYINPUT21), .A3(G169), .A4(new_n610), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(G179), .A3(new_n610), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n587), .A2(new_n390), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n579), .A2(new_n368), .A3(new_n542), .A4(new_n580), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n574), .B2(new_n586), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n616), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n458), .A2(new_n555), .A3(new_n630), .ZN(G372));
  NAND2_X1  g0431(.A1(new_n444), .A2(new_n446), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n440), .A2(new_n451), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT17), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n452), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n322), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n316), .A2(new_n392), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n361), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n359), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n372), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT98), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT98), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n644), .B(new_n372), .C1(new_n639), .C2(new_n641), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n458), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT97), .ZN(new_n648));
  INV_X1    g0448(.A(new_n473), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n500), .A2(new_n501), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n479), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n500), .A2(KEYINPUT92), .A3(new_n501), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT94), .B1(new_n653), .B2(new_n478), .ZN(new_n654));
  INV_X1    g0454(.A(new_n506), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n546), .ZN(new_n657));
  INV_X1    g0457(.A(new_n554), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n505), .A2(new_n506), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n554), .B1(new_n661), .B2(new_n649), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n657), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n648), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(KEYINPUT97), .A2(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n589), .ZN(new_n668));
  INV_X1    g0468(.A(new_n625), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n574), .A2(new_n586), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n626), .A3(new_n627), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n546), .A2(new_n549), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n662), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n674), .A3(new_n656), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n646), .B1(new_n647), .B2(new_n676), .ZN(G369));
  INV_X1    g0477(.A(G13), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G20), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n305), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n611), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n615), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n669), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n669), .B2(new_n687), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G330), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n670), .A2(new_n685), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n629), .B1(new_n696), .B2(new_n589), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n671), .A2(new_n685), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n669), .A2(new_n685), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n671), .B2(new_n685), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n701), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n210), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n486), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n216), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n686), .C1(new_n665), .C2(new_n675), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n663), .B1(new_n662), .B2(new_n657), .ZN(new_n715));
  NOR4_X1   g0515(.A1(new_n507), .A2(KEYINPUT26), .A3(new_n546), .A4(new_n554), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n715), .A2(new_n716), .A3(new_n507), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT101), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n656), .A2(new_n673), .A3(new_n658), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n589), .B1(new_n625), .B2(new_n629), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n555), .A2(KEYINPUT101), .A3(new_n672), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n685), .B1(new_n717), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n714), .B1(new_n724), .B2(new_n713), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n591), .A2(G179), .A3(new_n599), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT100), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT100), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n591), .A2(new_n599), .A3(new_n729), .A4(G179), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n463), .A2(new_n579), .A3(new_n470), .A4(new_n580), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n544), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n732), .A4(new_n730), .ZN(new_n736));
  AOI21_X1  g0536(.A(G179), .B1(new_n463), .B2(new_n470), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n622), .A2(new_n544), .A3(new_n587), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n685), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n662), .A2(new_n630), .A3(new_n673), .A4(new_n686), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n726), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n712), .B1(new_n748), .B2(G1), .ZN(G364));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n679), .B2(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n708), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n695), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n692), .A2(new_n693), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n341), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n216), .ZN(new_n764));
  INV_X1    g0564(.A(new_n241), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n764), .B1(G45), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT102), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n706), .A2(new_n345), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G355), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G116), .B2(new_n210), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n767), .B2(new_n770), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n213), .B1(G20), .B2(new_n390), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n760), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT103), .Z(new_n775));
  AOI21_X1  g0575(.A(new_n751), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(new_n368), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n780), .A2(KEYINPUT104), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(KEYINPUT104), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G77), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n778), .A2(new_n449), .A3(G200), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n345), .B1(new_n786), .B2(G58), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n449), .A2(new_n355), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n207), .A2(G179), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G87), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n778), .A2(new_n355), .A3(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n792), .B1(new_n794), .B2(new_n312), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n777), .A2(new_n788), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(G50), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n789), .A2(new_n449), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT106), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G107), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n785), .A2(new_n787), .A3(new_n798), .A4(new_n805), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n368), .A2(new_n355), .A3(KEYINPUT105), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT105), .B1(new_n368), .B2(new_n355), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n207), .B1(new_n810), .B2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n806), .B1(G97), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n809), .A2(new_n207), .A3(G190), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G159), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT32), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n812), .A2(G294), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n341), .B1(new_n779), .B2(G311), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n804), .A2(G283), .B1(G329), .B2(new_n814), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G326), .A2(new_n797), .B1(new_n791), .B2(G303), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT33), .B(G317), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n793), .A2(new_n821), .B1(new_n786), .B2(G322), .ZN(new_n822));
  AND4_X1   g0622(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n813), .A2(new_n816), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n773), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n776), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n754), .A2(new_n757), .B1(new_n762), .B2(new_n826), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n380), .A2(new_n686), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n392), .B1(new_n398), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n393), .A2(new_n686), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n676), .B2(new_n685), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n399), .B(new_n686), .C1(new_n665), .C2(new_n675), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n752), .B1(new_n834), .B2(new_n746), .ZN(new_n835));
  INV_X1    g0635(.A(new_n746), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n773), .A2(new_n758), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G77), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n803), .A2(new_n485), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n784), .B2(G116), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n812), .A2(G97), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n814), .A2(G311), .ZN(new_n845));
  INV_X1    g0645(.A(G283), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n345), .B1(new_n794), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n786), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n848), .A2(new_n577), .B1(new_n796), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n847), .B(new_n850), .C1(G107), .C2(new_n791), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n804), .A2(G68), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n202), .B2(new_n790), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT107), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n786), .A2(G143), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n793), .A2(G150), .B1(new_n797), .B2(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G159), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n858), .C1(new_n783), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n854), .A2(new_n855), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n345), .B1(new_n814), .B2(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n865), .B1(new_n329), .B2(new_n811), .C1(new_n860), .C2(new_n861), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n751), .B(new_n841), .C1(new_n867), .C2(new_n773), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n831), .A2(new_n758), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n838), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(G384));
  OAI21_X1  g0672(.A(G77), .B1(new_n329), .B2(new_n312), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n873), .A2(new_n216), .B1(G50), .B2(new_n312), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n678), .A3(new_n250), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT109), .Z(new_n876));
  OAI21_X1  g0676(.A(new_n514), .B1(new_n512), .B2(new_n515), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT35), .ZN(new_n878));
  OAI211_X1 g0678(.A(G116), .B(new_n214), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n876), .B1(new_n882), .B2(KEYINPUT108), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n315), .A2(new_n685), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n316), .A2(new_n321), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n315), .B(new_n685), .C1(new_n289), .C2(new_n322), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n833), .B2(new_n830), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n402), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n295), .A3(new_n419), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n426), .ZN(new_n894));
  INV_X1    g0694(.A(new_n683), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n636), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n898), .B2(new_n447), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n441), .A2(new_n683), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n894), .A2(new_n900), .B1(new_n440), .B2(new_n451), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT110), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n894), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n633), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT110), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n427), .A2(new_n437), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n427), .A2(new_n895), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n902), .A4(new_n633), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n890), .B1(new_n899), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n896), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n456), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n889), .A2(new_n917), .B1(new_n632), .B2(new_n683), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n633), .B1(new_n440), .B2(new_n441), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n440), .A2(new_n683), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n910), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n636), .B2(new_n632), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n890), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n316), .A2(new_n685), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n918), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n725), .A2(new_n458), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n646), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n829), .A2(new_n830), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n745), .A2(new_n887), .A3(KEYINPUT40), .A4(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n745), .A2(new_n936), .A3(new_n887), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n912), .B2(new_n916), .ZN(new_n941));
  OAI211_X1 g0741(.A(G330), .B(new_n939), .C1(new_n941), .C2(KEYINPUT40), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n458), .A2(new_n836), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT111), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n937), .B1(new_n916), .B2(new_n925), .ZN(new_n946));
  INV_X1    g0746(.A(new_n940), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n899), .A2(new_n890), .A3(new_n911), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n914), .B2(new_n915), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n458), .A3(new_n745), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n935), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n305), .B2(new_n679), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n945), .A2(new_n935), .A3(new_n954), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n883), .B1(KEYINPUT108), .B2(new_n882), .C1(new_n956), .C2(new_n957), .ZN(G367));
  AND2_X1   g0758(.A1(new_n763), .A2(new_n233), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n774), .B1(new_n210), .B2(new_n378), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n784), .A2(G50), .B1(G137), .B2(new_n814), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G143), .A2(new_n797), .B1(new_n791), .B2(G58), .ZN(new_n962));
  INV_X1    g0762(.A(G150), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(new_n848), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n345), .B(new_n964), .C1(G159), .C2(new_n793), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n804), .A2(G77), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n811), .A2(new_n312), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n961), .A2(new_n965), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n786), .A2(G303), .B1(new_n797), .B2(G311), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n577), .B2(new_n794), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n790), .A2(new_n601), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT46), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(new_n784), .C2(G283), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n814), .A2(G317), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n345), .C1(new_n494), .C2(new_n803), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT115), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n974), .B(new_n978), .C1(new_n558), .C2(new_n811), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n969), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT47), .Z(new_n982));
  OAI221_X1 g0782(.A(new_n752), .B1(new_n959), .B2(new_n960), .C1(new_n982), .C2(new_n825), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT116), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n551), .A2(new_n685), .ZN(new_n985));
  MUX2_X1   g0785(.A(new_n662), .B(new_n507), .S(new_n985), .Z(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(new_n761), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n750), .B(KEYINPUT114), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n673), .B1(new_n547), .B2(new_n686), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n657), .A2(new_n685), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n704), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n704), .A2(new_n993), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n700), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n700), .B1(new_n995), .B2(new_n998), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT113), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT112), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n699), .B2(new_n702), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n694), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n694), .B2(new_n1003), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n1007), .A2(new_n703), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n703), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n747), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n707), .B(KEYINPUT41), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n990), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n993), .A2(new_n703), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n546), .B1(new_n991), .B2(new_n671), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1016), .A2(KEYINPUT42), .B1(new_n686), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1017), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n700), .A2(new_n993), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n989), .B1(new_n1015), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT117), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(G387));
  INV_X1    g0827(.A(new_n709), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n768), .A2(new_n1028), .B1(new_n558), .B2(new_n706), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n376), .A2(new_n202), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n464), .B1(new_n312), .B2(new_n301), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1031), .A2(new_n1028), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n763), .B1(new_n230), .B2(new_n464), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n751), .B1(new_n1035), .B2(new_n775), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n699), .B2(new_n761), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n341), .B1(new_n780), .B2(new_n312), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n848), .A2(new_n202), .B1(new_n796), .B2(new_n859), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G77), .C2(new_n791), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n814), .A2(G150), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n331), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n804), .A2(G97), .B1(new_n1042), .B2(new_n793), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n812), .A2(new_n480), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n784), .A2(G303), .B1(G317), .B2(new_n786), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT118), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(KEYINPUT118), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n793), .A2(G311), .B1(new_n797), .B2(G322), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n811), .A2(new_n846), .B1(new_n577), .B2(new_n790), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(KEYINPUT49), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n814), .A2(G326), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n341), .B1(new_n804), .B2(G116), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT49), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1045), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1037), .B1(new_n1060), .B2(new_n773), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n990), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1012), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1012), .A2(new_n748), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n707), .B(KEYINPUT119), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1012), .A2(new_n748), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(G393));
  INV_X1    g0868(.A(new_n1001), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n999), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1002), .A2(new_n1012), .A3(new_n748), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1072), .A3(new_n1065), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n993), .A2(new_n760), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n238), .A2(new_n763), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n774), .B1(new_n494), .B2(new_n210), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n752), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n341), .B1(new_n791), .B2(G283), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G294), .A2(new_n779), .B1(new_n793), .B2(G303), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n805), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G322), .B2(new_n814), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n786), .A2(G311), .B1(new_n797), .B2(G317), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(new_n601), .C2(new_n811), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n784), .A2(new_n376), .B1(G50), .B2(new_n793), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT120), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n341), .B1(new_n790), .B2(new_n312), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1087), .B(new_n842), .C1(G143), .C2(new_n814), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n786), .A2(G159), .B1(new_n797), .B2(G150), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  NAND2_X1  g0890(.A1(new_n812), .A2(G77), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1084), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1077), .B1(new_n1093), .B2(new_n773), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1002), .A2(new_n1062), .B1(new_n1074), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1073), .A2(new_n1095), .ZN(G390));
  NAND4_X1  g0896(.A1(new_n745), .A2(new_n887), .A3(G330), .A4(new_n936), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n399), .A2(new_n686), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n656), .B1(new_n719), .B2(new_n720), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n666), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n662), .B2(new_n657), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT97), .B1(new_n715), .B2(new_n716), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n830), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n887), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n929), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n928), .A2(new_n930), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n721), .A2(new_n722), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n660), .A2(new_n656), .A3(new_n664), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n686), .B(new_n829), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n888), .B1(new_n1112), .B2(new_n830), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n926), .A2(new_n1108), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1098), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1106), .B1(new_n724), .B2(new_n829), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1108), .B(new_n926), .C1(new_n1117), .C2(new_n888), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n928), .A2(new_n930), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n889), .A2(new_n929), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1097), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n745), .A2(G330), .A3(new_n936), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n888), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n1097), .B1(new_n833), .B2(new_n830), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(new_n1097), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n933), .A2(new_n646), .A3(new_n943), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1122), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1065), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1116), .A2(new_n1121), .A3(new_n1062), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n752), .B1(new_n1042), .B2(new_n840), .ZN(new_n1135));
  INV_X1    g0935(.A(G132), .ZN(new_n1136));
  INV_X1    g0936(.A(G137), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1136), .A2(new_n848), .B1(new_n794), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n345), .B(new_n1138), .C1(G128), .C2(new_n797), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n814), .A2(G125), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n859), .C2(new_n811), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n790), .A2(new_n963), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT53), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1143), .B1(new_n202), .B2(new_n803), .C1(new_n783), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n814), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n853), .B1(new_n1146), .B2(new_n577), .C1(new_n783), .C2(new_n494), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n558), .A2(new_n794), .B1(new_n848), .B2(new_n601), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G283), .B2(new_n797), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1149), .A2(new_n345), .A3(new_n792), .A4(new_n1091), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1141), .A2(new_n1145), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1135), .B1(new_n1151), .B2(new_n773), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1119), .B2(new_n759), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1133), .A2(new_n1134), .A3(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n370), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n363), .B(new_n895), .C1(new_n641), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n363), .A2(new_n895), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n362), .A2(new_n370), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n952), .B2(G330), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n942), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n932), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n952), .A2(G330), .A3(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n942), .A2(new_n1166), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1169), .A2(new_n1170), .A3(new_n931), .A4(new_n918), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1166), .A2(new_n758), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n752), .B1(G50), .B2(new_n840), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n793), .A2(G132), .B1(new_n797), .B2(G125), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n790), .A2(new_n1144), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n786), .B2(G128), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n1137), .C2(new_n780), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G150), .B2(new_n812), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT122), .B(G124), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n244), .B(new_n245), .C1(new_n1146), .C2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G159), .B2(new_n804), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n804), .A2(G58), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n345), .A2(new_n245), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G77), .B2(new_n791), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT121), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1187), .B(new_n1191), .C1(new_n846), .C2(new_n1146), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n786), .A2(G107), .B1(new_n797), .B2(G116), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n494), .B2(new_n794), .C1(new_n378), .C2(new_n780), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1190), .A2(KEYINPUT121), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1192), .A2(new_n967), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT58), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT58), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1188), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1186), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1174), .B1(new_n1200), .B2(new_n773), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1172), .A2(new_n1062), .B1(new_n1173), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1128), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1132), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1172), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT57), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1065), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n1204), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT123), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(KEYINPUT123), .B(new_n1208), .C1(new_n1209), .C2(new_n1204), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1202), .B1(new_n1212), .B2(new_n1213), .ZN(G375));
  INV_X1    g1014(.A(new_n1127), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n990), .B(KEYINPUT124), .Z(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n888), .A2(new_n758), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n752), .B1(G68), .B2(new_n840), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n966), .B1(new_n1146), .B2(new_n849), .C1(new_n783), .C2(new_n558), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n848), .A2(new_n846), .B1(new_n494), .B2(new_n790), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G294), .B2(new_n797), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n341), .B1(new_n793), .B2(G116), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1044), .A3(new_n1223), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n1137), .A2(new_n848), .B1(new_n794), .B2(new_n1144), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n780), .A2(new_n963), .B1(new_n1136), .B2(new_n796), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n345), .B1(new_n791), .B2(G159), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n814), .A2(G128), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1227), .A2(new_n1187), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n811), .A2(new_n202), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1220), .A2(new_n1224), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1219), .B1(new_n1232), .B2(new_n773), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1215), .A2(new_n1217), .B1(new_n1218), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1014), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1130), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1215), .A2(new_n1203), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  INV_X1    g1038(.A(G396), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n1063), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1240));
  OR3_X1    g1040(.A1(G390), .A2(G384), .A3(new_n1240), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(G387), .A2(new_n1241), .A3(G378), .A4(G381), .ZN(new_n1242));
  INV_X1    g1042(.A(G375), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT125), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1244), .B(new_n1245), .ZN(G407));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G378), .A2(G343), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G407), .A2(new_n1249), .ZN(G409));
  NOR2_X1   g1050(.A1(new_n1247), .A2(G343), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G378), .B(new_n1202), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1252));
  INV_X1    g1052(.A(G378), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1173), .A2(new_n1201), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1172), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1216), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1205), .A2(new_n1014), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1253), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1252), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1237), .B1(KEYINPUT60), .B2(new_n1130), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT60), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1065), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1234), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(new_n871), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1251), .A2(G2897), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1265), .B(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1260), .B2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n1239), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1025), .B2(G390), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n748), .B1(new_n1070), .B2(new_n1011), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1062), .B1(new_n1271), .B2(new_n1235), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1024), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n988), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1026), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1025), .A2(KEYINPUT117), .ZN(new_n1276));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1270), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1025), .B(G390), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1269), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1264), .B(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1259), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1251), .B(new_n1265), .C1(new_n1252), .C2(new_n1258), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT63), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1268), .A2(new_n1285), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1286), .B(new_n1266), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1259), .ZN(new_n1295));
  AND2_X1   g1095(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1290), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1287), .A2(new_n1297), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1295), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1292), .B1(new_n1301), .B2(new_n1285), .ZN(G405));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1253), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1303), .A2(new_n1252), .A3(new_n1265), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1265), .B1(new_n1303), .B2(new_n1252), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1285), .ZN(G402));
endmodule


