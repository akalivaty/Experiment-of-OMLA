

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n699) );
  XNOR2_X1 U552 ( .A(n700), .B(n699), .ZN(n702) );
  INV_X1 U553 ( .A(n738), .ZN(n724) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT32), .ZN(n745) );
  XNOR2_X1 U555 ( .A(n746), .B(n745), .ZN(n755) );
  NOR2_X2 U556 ( .A1(G2105), .A2(n521), .ZN(n874) );
  NOR2_X1 U557 ( .A1(G651), .A2(n636), .ZN(n652) );
  NOR2_X1 U558 ( .A1(n527), .A2(n526), .ZN(G160) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XOR2_X1 U560 ( .A(KEYINPUT17), .B(n517), .Z(n875) );
  NAND2_X1 U561 ( .A1(n875), .A2(G137), .ZN(n520) );
  INV_X1 U562 ( .A(G2104), .ZN(n521) );
  NAND2_X1 U563 ( .A1(G101), .A2(n874), .ZN(n518) );
  XOR2_X1 U564 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U565 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U566 ( .A1(n521), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U567 ( .A(n522), .B(KEYINPUT65), .ZN(n878) );
  NAND2_X1 U568 ( .A1(n878), .A2(G125), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X1 U570 ( .A(KEYINPUT66), .B(n523), .Z(n879) );
  NAND2_X1 U571 ( .A1(G113), .A2(n879), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U573 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U574 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U575 ( .A1(n875), .A2(G135), .ZN(n528) );
  XNOR2_X1 U576 ( .A(KEYINPUT76), .B(n528), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n878), .A2(G123), .ZN(n529) );
  XNOR2_X1 U578 ( .A(KEYINPUT18), .B(n529), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U580 ( .A(n532), .B(KEYINPUT77), .ZN(n538) );
  NAND2_X1 U581 ( .A1(n874), .A2(G99), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT78), .ZN(n535) );
  NAND2_X1 U583 ( .A1(G111), .A2(n879), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U585 ( .A(KEYINPUT79), .B(n536), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U587 ( .A(n539), .B(KEYINPUT80), .ZN(n993) );
  XNOR2_X1 U588 ( .A(n993), .B(G2096), .ZN(n540) );
  OR2_X1 U589 ( .A1(G2100), .A2(n540), .ZN(G156) );
  INV_X1 U590 ( .A(G132), .ZN(G219) );
  INV_X1 U591 ( .A(G82), .ZN(G220) );
  INV_X1 U592 ( .A(G108), .ZN(G238) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n636) );
  NAND2_X1 U594 ( .A1(G53), .A2(n652), .ZN(n543) );
  INV_X1 U595 ( .A(G651), .ZN(n544) );
  NOR2_X1 U596 ( .A1(G543), .A2(n544), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n541), .Z(n648) );
  NAND2_X1 U598 ( .A1(G65), .A2(n648), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n549) );
  NOR2_X1 U600 ( .A1(n636), .A2(n544), .ZN(n644) );
  NAND2_X1 U601 ( .A1(G78), .A2(n644), .ZN(n547) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n545) );
  XNOR2_X1 U603 ( .A(n545), .B(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U604 ( .A1(G91), .A2(n645), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n705) );
  INV_X1 U607 ( .A(n705), .ZN(G299) );
  NAND2_X1 U608 ( .A1(n875), .A2(G138), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G102), .A2(n874), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT89), .B(n550), .Z(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n878), .A2(G126), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G114), .A2(n879), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U615 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U618 ( .A(G223), .ZN(n817) );
  NAND2_X1 U619 ( .A1(n817), .A2(G567), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  XNOR2_X1 U621 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G81), .A2(n645), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G68), .A2(n644), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n648), .A2(G56), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n652), .A2(G43), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n911) );
  INV_X1 U632 ( .A(n911), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n569), .A2(G860), .ZN(G153) );
  NAND2_X1 U634 ( .A1(G52), .A2(n652), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G64), .A2(n648), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G77), .A2(n644), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G90), .A2(n645), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(KEYINPUT68), .B(n577), .ZN(G171) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(n652), .A2(G54), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G79), .A2(n644), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G92), .A2(n645), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n648), .A2(G66), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT70), .B(n580), .Z(n581) );
  NOR2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U652 ( .A(KEYINPUT15), .B(n585), .Z(n921) );
  INV_X1 U653 ( .A(n921), .ZN(n611) );
  NOR2_X1 U654 ( .A1(n611), .A2(G868), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT71), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(G284) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(KEYINPUT7), .ZN(n601) );
  NAND2_X1 U659 ( .A1(G51), .A2(n652), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G63), .A2(n648), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n591), .B(KEYINPUT6), .ZN(n592) );
  XNOR2_X1 U663 ( .A(n592), .B(KEYINPUT73), .ZN(n599) );
  XNOR2_X1 U664 ( .A(KEYINPUT5), .B(KEYINPUT72), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G89), .A2(n645), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT4), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G76), .A2(n644), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n601), .B(n600), .ZN(G168) );
  XOR2_X1 U672 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U673 ( .A1(G868), .A2(G286), .ZN(n603) );
  INV_X1 U674 ( .A(G868), .ZN(n663) );
  NAND2_X1 U675 ( .A1(G299), .A2(n663), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G297) );
  INV_X1 U677 ( .A(G559), .ZN(n604) );
  NOR2_X1 U678 ( .A1(G860), .A2(n604), .ZN(n605) );
  XNOR2_X1 U679 ( .A(KEYINPUT75), .B(n605), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n606), .A2(n611), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n911), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G868), .A2(n611), .ZN(n608) );
  NOR2_X1 U684 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U686 ( .A1(n611), .A2(G559), .ZN(n661) );
  XNOR2_X1 U687 ( .A(n911), .B(n661), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n612), .A2(G860), .ZN(n619) );
  NAND2_X1 U689 ( .A1(G80), .A2(n644), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G93), .A2(n645), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G55), .A2(n652), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G67), .A2(n648), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n664) );
  XOR2_X1 U696 ( .A(n619), .B(n664), .Z(G145) );
  NAND2_X1 U697 ( .A1(G73), .A2(n644), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT2), .B(n620), .Z(n621) );
  XNOR2_X1 U699 ( .A(n621), .B(KEYINPUT83), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G86), .A2(n645), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G48), .A2(n652), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G61), .A2(n648), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U706 ( .A(KEYINPUT84), .B(n628), .Z(G305) );
  NAND2_X1 U707 ( .A1(G75), .A2(n644), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G88), .A2(n645), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(n631), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n652), .A2(G50), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G62), .A2(n648), .ZN(n632) );
  AND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(G303) );
  INV_X1 U715 ( .A(G303), .ZN(G166) );
  NAND2_X1 U716 ( .A1(n636), .A2(G87), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n637), .B(KEYINPUT82), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n648), .A2(n640), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G49), .A2(n652), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT81), .B(n641), .Z(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G72), .A2(n644), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G85), .A2(n645), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G60), .A2(n648), .ZN(n649) );
  XNOR2_X1 U728 ( .A(KEYINPUT67), .B(n649), .ZN(n650) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n652), .A2(G47), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(G290) );
  XNOR2_X1 U732 ( .A(n664), .B(G166), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(G288), .ZN(n656) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(n656), .ZN(n658) );
  XNOR2_X1 U735 ( .A(G290), .B(n705), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U737 ( .A(G305), .B(n659), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n911), .B(n660), .ZN(n892) );
  XOR2_X1 U739 ( .A(n892), .B(n661), .Z(n662) );
  NOR2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U741 ( .A1(G868), .A2(n664), .ZN(n665) );
  NOR2_X1 U742 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n670), .A2(G2072), .ZN(G158) );
  NAND2_X1 U748 ( .A1(G120), .A2(G69), .ZN(n671) );
  NOR2_X1 U749 ( .A1(G238), .A2(n671), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n672), .A2(G57), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(KEYINPUT86), .ZN(n823) );
  NAND2_X1 U752 ( .A1(n823), .A2(G567), .ZN(n674) );
  XNOR2_X1 U753 ( .A(n674), .B(KEYINPUT87), .ZN(n679) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n675) );
  XNOR2_X1 U755 ( .A(KEYINPUT22), .B(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(n676), .A2(G96), .ZN(n677) );
  OR2_X1 U757 ( .A1(G218), .A2(n677), .ZN(n824) );
  AND2_X1 U758 ( .A1(G2106), .A2(n824), .ZN(n678) );
  NOR2_X1 U759 ( .A1(n679), .A2(n678), .ZN(G319) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n681) );
  INV_X1 U761 ( .A(G319), .ZN(n680) );
  NOR2_X1 U762 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U763 ( .A(n682), .B(KEYINPUT88), .ZN(n822) );
  NAND2_X1 U764 ( .A1(G36), .A2(n822), .ZN(G176) );
  NAND2_X1 U765 ( .A1(G104), .A2(n874), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G140), .A2(n875), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U768 ( .A(KEYINPUT34), .B(n685), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n878), .A2(G128), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G116), .A2(n879), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U772 ( .A(KEYINPUT90), .B(n688), .Z(n689) );
  XNOR2_X1 U773 ( .A(KEYINPUT35), .B(n689), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U775 ( .A(KEYINPUT36), .B(n692), .ZN(n862) );
  XNOR2_X1 U776 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U777 ( .A1(n862), .A2(n810), .ZN(n989) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n696) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n694) );
  NOR2_X1 U780 ( .A1(n696), .A2(n694), .ZN(n812) );
  NAND2_X1 U781 ( .A1(n989), .A2(n812), .ZN(n693) );
  XOR2_X1 U782 ( .A(KEYINPUT91), .B(n693), .Z(n808) );
  INV_X1 U783 ( .A(n808), .ZN(n800) );
  INV_X1 U784 ( .A(n694), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n738) );
  NAND2_X1 U786 ( .A1(G8), .A2(n738), .ZN(n768) );
  XNOR2_X1 U787 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n723) );
  INV_X1 U788 ( .A(KEYINPUT27), .ZN(n698) );
  NAND2_X1 U789 ( .A1(G2072), .A2(n724), .ZN(n697) );
  XNOR2_X1 U790 ( .A(n698), .B(n697), .ZN(n700) );
  XNOR2_X1 U791 ( .A(G1956), .B(KEYINPUT99), .ZN(n972) );
  NOR2_X1 U792 ( .A1(n972), .A2(n724), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n704) );
  XOR2_X1 U795 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n703) );
  XNOR2_X1 U796 ( .A(n704), .B(n703), .ZN(n721) );
  NAND2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n719) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n738), .ZN(n708) );
  NAND2_X1 U799 ( .A1(G2067), .A2(n724), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n921), .A2(n713), .ZN(n717) );
  INV_X1 U802 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U803 ( .A1(n738), .A2(n942), .ZN(n709) );
  XOR2_X1 U804 ( .A(n709), .B(KEYINPUT26), .Z(n711) );
  NAND2_X1 U805 ( .A1(n738), .A2(G1341), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U807 ( .A1(n911), .A2(n712), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n921), .A2(n713), .ZN(n714) );
  OR2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U813 ( .A(n723), .B(n722), .ZN(n728) );
  XOR2_X1 U814 ( .A(G1961), .B(KEYINPUT96), .Z(n967) );
  NAND2_X1 U815 ( .A1(n967), .A2(n738), .ZN(n726) );
  XNOR2_X1 U816 ( .A(KEYINPUT25), .B(G2078), .ZN(n949) );
  NAND2_X1 U817 ( .A1(n724), .A2(n949), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n732), .A2(G171), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n737) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n768), .ZN(n750) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n738), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n750), .A2(n747), .ZN(n729) );
  NAND2_X1 U824 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U826 ( .A1(G168), .A2(n731), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n732), .A2(G171), .ZN(n733) );
  NOR2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U829 ( .A(KEYINPUT31), .B(n735), .Z(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n749) );
  NAND2_X1 U831 ( .A1(n749), .A2(G286), .ZN(n743) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n768), .ZN(n740) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U834 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U835 ( .A1(n741), .A2(G303), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U837 ( .A1(n744), .A2(G8), .ZN(n746) );
  NAND2_X1 U838 ( .A1(G8), .A2(n747), .ZN(n748) );
  XOR2_X1 U839 ( .A(KEYINPUT95), .B(n748), .Z(n753) );
  INV_X1 U840 ( .A(n749), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n769) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U846 ( .A1(n760), .A2(n756), .ZN(n915) );
  NAND2_X1 U847 ( .A1(n769), .A2(n915), .ZN(n757) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n914) );
  NAND2_X1 U849 ( .A1(n757), .A2(n914), .ZN(n758) );
  NOR2_X1 U850 ( .A1(n768), .A2(n758), .ZN(n759) );
  OR2_X1 U851 ( .A1(n759), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n761), .A2(n768), .ZN(n763) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n929) );
  INV_X1 U855 ( .A(n929), .ZN(n762) );
  NOR2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n778) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U859 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n776) );
  INV_X1 U861 ( .A(n768), .ZN(n774) );
  INV_X1 U862 ( .A(n769), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G166), .A2(G8), .ZN(n770) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n770), .ZN(n771) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n798) );
  NAND2_X1 U869 ( .A1(G141), .A2(n875), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G129), .A2(n878), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n874), .A2(G105), .ZN(n781) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G117), .A2(n879), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n858) );
  NAND2_X1 U877 ( .A1(G1996), .A2(n858), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G107), .A2(n879), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G95), .A2(n874), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G119), .A2(n878), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n875), .A2(G131), .ZN(n788) );
  XOR2_X1 U883 ( .A(KEYINPUT92), .B(n788), .Z(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U886 ( .A(KEYINPUT93), .B(n793), .Z(n887) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n887), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n995) );
  NAND2_X1 U889 ( .A1(n995), .A2(n812), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT94), .B(n796), .Z(n805) );
  INV_X1 U891 ( .A(n805), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n802) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n913) );
  NAND2_X1 U895 ( .A1(n913), .A2(n812), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n815) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n858), .ZN(n1001) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n887), .ZN(n988) );
  NOR2_X1 U900 ( .A1(n803), .A2(n988), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n1001), .A2(n806), .ZN(n807) );
  XNOR2_X1 U903 ( .A(KEYINPUT39), .B(n807), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n862), .A2(n810), .ZN(n992) );
  NAND2_X1 U906 ( .A1(n811), .A2(n992), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n817), .ZN(G217) );
  INV_X1 U911 ( .A(G661), .ZN(n819) );
  NAND2_X1 U912 ( .A1(G2), .A2(G15), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U914 ( .A(KEYINPUT104), .B(n820), .Z(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(G188) );
  XNOR2_X1 U917 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U918 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XNOR2_X1 U919 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  XOR2_X1 U923 ( .A(G2096), .B(G2072), .Z(n826) );
  XNOR2_X1 U924 ( .A(G2067), .B(G2090), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n826), .B(n825), .ZN(n836) );
  XOR2_X1 U926 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n828) );
  XNOR2_X1 U927 ( .A(G2678), .B(KEYINPUT111), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U929 ( .A(G2100), .B(KEYINPUT43), .Z(n830) );
  XNOR2_X1 U930 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U932 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2078), .B(G2084), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n836), .B(n835), .Z(G227) );
  XOR2_X1 U936 ( .A(KEYINPUT112), .B(KEYINPUT115), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n839), .B(KEYINPUT113), .Z(n841) );
  XNOR2_X1 U940 ( .A(G1956), .B(G1961), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n849) );
  XOR2_X1 U942 ( .A(G1976), .B(G1981), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1971), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2474), .B(G1966), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U948 ( .A(n847), .B(n846), .Z(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G112), .A2(n879), .ZN(n856) );
  NAND2_X1 U951 ( .A1(G100), .A2(n874), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G136), .A2(n875), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n878), .A2(G124), .ZN(n852) );
  XOR2_X1 U955 ( .A(KEYINPUT44), .B(n852), .Z(n853) );
  NOR2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U958 ( .A(KEYINPUT116), .B(n857), .Z(G162) );
  XNOR2_X1 U959 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT46), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n864) );
  XNOR2_X1 U963 ( .A(G164), .B(G160), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n873) );
  NAND2_X1 U965 ( .A1(n878), .A2(G130), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G118), .A2(n879), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G106), .A2(n874), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G142), .A2(n875), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT45), .B(n869), .Z(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n886) );
  NAND2_X1 U974 ( .A1(G103), .A2(n874), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G139), .A2(n875), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U977 ( .A1(n878), .A2(G127), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n996) );
  XNOR2_X1 U982 ( .A(n996), .B(n993), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U984 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U985 ( .A(G162), .B(n889), .ZN(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G301), .B(G286), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n891), .B(n921), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U990 ( .A1(G37), .A2(n894), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2430), .B(G2451), .Z(n896) );
  XNOR2_X1 U992 ( .A(G2446), .B(G2427), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n903) );
  XOR2_X1 U994 ( .A(G2438), .B(G2435), .Z(n898) );
  XNOR2_X1 U995 ( .A(G2443), .B(KEYINPUT103), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(G2454), .Z(n901) );
  XNOR2_X1 U998 ( .A(G1348), .B(G1341), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(n904), .A2(G14), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n910), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G57), .ZN(G237) );
  INV_X1 U1010 ( .A(n910), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(KEYINPUT56), .B(G16), .ZN(n935) );
  XNOR2_X1 U1012 ( .A(n911), .B(G1341), .ZN(n928) );
  XNOR2_X1 U1013 ( .A(G1956), .B(G299), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n920) );
  AND2_X1 U1015 ( .A1(G303), .A2(G1971), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT122), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(G171), .B(G1961), .ZN(n923) );
  XOR2_X1 U1021 ( .A(G1348), .B(n921), .Z(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT123), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(G168), .B(G1966), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT57), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n1018) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n1010) );
  XOR2_X1 U1032 ( .A(G34), .B(KEYINPUT121), .Z(n937) );
  XNOR2_X1 U1033 ( .A(G2084), .B(KEYINPUT54), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n937), .B(n936), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n956) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G1991), .B(G25), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G32), .B(n942), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n943), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT118), .B(G2072), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G33), .B(n944), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G27), .B(n949), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT119), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(n953), .B(KEYINPUT120), .Z(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n1010), .B(n957), .ZN(n959) );
  INV_X1 U1053 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n960), .ZN(n1016) );
  XOR2_X1 U1056 ( .A(G16), .B(KEYINPUT124), .Z(n987) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n964) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G22), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G23), .B(G1976), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(n966), .B(n965), .ZN(n971) );
  XOR2_X1 U1064 ( .A(n967), .B(G5), .Z(n969) );
  XNOR2_X1 U1065 ( .A(G21), .B(G1966), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n984) );
  XOR2_X1 U1068 ( .A(n972), .B(G20), .Z(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT59), .B(G4), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n973), .B(KEYINPUT125), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n974), .B(G1348), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G1341), .B(G19), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(n981), .B(KEYINPUT60), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n982), .B(KEYINPUT126), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(KEYINPUT61), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n1014) );
  XNOR2_X1 U1082 ( .A(G160), .B(G2084), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n1008) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1006) );
  XOR2_X1 U1087 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1088 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1090 ( .A(KEYINPUT50), .B(n999), .Z(n1004) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT51), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT52), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(G29), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

